module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 325:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 325:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 325:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 262:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 262:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 262:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 262:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 262:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 262:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 264:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 264:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 264:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 264:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 264:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 264:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 288:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 292:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 292:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 292:33:@104.4]
  wire  _T_57; // @[Counter.scala 294:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 300:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 300:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 300:74:@118.4]
  FF bases_0 ( // @[Counter.scala 262:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 264:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 288:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 292:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 292:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 292:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh50); // @[Counter.scala 294:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 300:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 300:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 300:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh50); // @[Counter.scala 334:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 300:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 282:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 285:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 265:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 266:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 267:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@390.2]
  input   clock, // @[:@391.4]
  input   reset, // @[:@392.4]
  input   io_enable, // @[:@393.4]
  output  io_done, // @[:@393.4]
  input   io_rst, // @[:@393.4]
  input   io_ctrDone, // @[:@393.4]
  output  io_ctrInc, // @[:@393.4]
  input   io_doneIn_0, // @[:@393.4]
  input   io_doneIn_1, // @[:@393.4]
  input   io_doneIn_2, // @[:@393.4]
  output  io_enableOut_0, // @[:@393.4]
  output  io_enableOut_1, // @[:@393.4]
  output  io_enableOut_2, // @[:@393.4]
  output  io_childAck_0, // @[:@393.4]
  output  io_childAck_1, // @[:@393.4]
  output  io_childAck_2 // @[:@393.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@396.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@396.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@396.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@396.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@396.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@396.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@399.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@399.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@399.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@399.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@399.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@399.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@402.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@402.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@402.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@402.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@402.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@402.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@405.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@405.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@405.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@405.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@405.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@405.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@408.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@408.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@408.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@408.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@408.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@408.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@411.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@411.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@411.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@411.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@411.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@411.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@452.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@452.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@452.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@452.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@452.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@452.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@455.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@455.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@455.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@455.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@455.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@455.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@458.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@458.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@458.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@458.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@458.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@458.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@497.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@497.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@497.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@497.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@497.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@630.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@630.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@630.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@630.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@630.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@647.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@647.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@647.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@647.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@647.4]
  wire  _T_77; // @[Controllers.scala 80:47:@414.4]
  wire  allDone; // @[Controllers.scala 80:47:@415.4]
  wire  _T_78; // @[Controllers.scala 81:26:@416.4]
  wire  finished; // @[Controllers.scala 81:37:@417.4]
  wire  synchronize; // @[package.scala 96:25:@502.4 package.scala 96:25:@503.4]
  wire  _T_168; // @[Controllers.scala 128:33:@511.4]
  wire  _T_170; // @[Controllers.scala 128:54:@512.4]
  wire  _T_171; // @[Controllers.scala 128:52:@513.4]
  wire  _T_172; // @[Controllers.scala 128:66:@514.4]
  wire  _T_174; // @[Controllers.scala 128:98:@516.4]
  wire  _T_175; // @[Controllers.scala 128:96:@517.4]
  wire  _T_177; // @[Controllers.scala 128:123:@518.4]
  wire  _T_179; // @[Controllers.scala 129:48:@521.4]
  wire  _T_184; // @[Controllers.scala 130:52:@526.4]
  wire  _T_185; // @[Controllers.scala 130:50:@527.4]
  wire  _T_193; // @[Controllers.scala 130:129:@533.4]
  wire  _T_196; // @[Controllers.scala 131:45:@536.4]
  wire  _T_199; // @[Controllers.scala 135:80:@540.4]
  wire  _T_200; // @[Controllers.scala 135:78:@541.4]
  wire  _T_202; // @[Controllers.scala 135:105:@542.4]
  wire  _T_203; // @[Controllers.scala 135:103:@543.4]
  wire  _T_204; // @[Controllers.scala 135:119:@544.4]
  wire  _T_206; // @[Controllers.scala 135:51:@546.4]
  wire  _T_227; // @[Controllers.scala 135:80:@567.4]
  wire  _T_228; // @[Controllers.scala 135:78:@568.4]
  wire  _T_230; // @[Controllers.scala 135:105:@569.4]
  wire  _T_231; // @[Controllers.scala 135:103:@570.4]
  wire  _T_232; // @[Controllers.scala 135:119:@571.4]
  wire  _T_234; // @[Controllers.scala 135:51:@573.4]
  wire  _T_258; // @[Controllers.scala 213:68:@600.4]
  wire  _T_260; // @[Controllers.scala 213:90:@602.4]
  wire  _T_262; // @[Controllers.scala 213:132:@604.4]
  wire  _T_263; // @[Controllers.scala 213:130:@605.4]
  wire  _T_264; // @[Controllers.scala 213:156:@606.4]
  wire  _T_266; // @[Controllers.scala 213:68:@609.4]
  wire  _T_268; // @[Controllers.scala 213:90:@611.4]
  wire  _T_274; // @[Controllers.scala 213:68:@617.4]
  wire  _T_276; // @[Controllers.scala 213:90:@619.4]
  wire  _T_283; // @[package.scala 100:49:@625.4]
  reg  _T_286; // @[package.scala 48:56:@626.4]
  reg [31:0] _RAND_0;
  reg  _T_300; // @[package.scala 48:56:@644.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@396.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@399.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@402.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@405.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@408.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@411.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@452.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@455.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@458.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@497.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@630.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@647.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@414.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@415.4]
  assign _T_78 = allDone | io_done; // @[Controllers.scala 81:26:@416.4]
  assign finished = _T_78 | done_2_io_input_set; // @[Controllers.scala 81:37:@417.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@502.4 package.scala 96:25:@503.4]
  assign _T_168 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@511.4]
  assign _T_170 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@512.4]
  assign _T_171 = _T_168 & _T_170; // @[Controllers.scala 128:52:@513.4]
  assign _T_172 = _T_171 & io_enable; // @[Controllers.scala 128:66:@514.4]
  assign _T_174 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@516.4]
  assign _T_175 = _T_172 & _T_174; // @[Controllers.scala 128:96:@517.4]
  assign _T_177 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@518.4]
  assign _T_179 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@521.4]
  assign _T_184 = synchronize == 1'h0; // @[Controllers.scala 130:52:@526.4]
  assign _T_185 = io_doneIn_0 & _T_184; // @[Controllers.scala 130:50:@527.4]
  assign _T_193 = finished == 1'h0; // @[Controllers.scala 130:129:@533.4]
  assign _T_196 = io_rst == 1'h0; // @[Controllers.scala 131:45:@536.4]
  assign _T_199 = ~ iterDone_1_io_output; // @[Controllers.scala 135:80:@540.4]
  assign _T_200 = iterDone_0_io_output & _T_199; // @[Controllers.scala 135:78:@541.4]
  assign _T_202 = io_doneIn_1 == 1'h0; // @[Controllers.scala 135:105:@542.4]
  assign _T_203 = _T_200 & _T_202; // @[Controllers.scala 135:103:@543.4]
  assign _T_204 = _T_203 & io_enable; // @[Controllers.scala 135:119:@544.4]
  assign _T_206 = io_doneIn_0 | _T_204; // @[Controllers.scala 135:51:@546.4]
  assign _T_227 = ~ iterDone_2_io_output; // @[Controllers.scala 135:80:@567.4]
  assign _T_228 = iterDone_1_io_output & _T_227; // @[Controllers.scala 135:78:@568.4]
  assign _T_230 = io_doneIn_2 == 1'h0; // @[Controllers.scala 135:105:@569.4]
  assign _T_231 = _T_228 & _T_230; // @[Controllers.scala 135:103:@570.4]
  assign _T_232 = _T_231 & io_enable; // @[Controllers.scala 135:119:@571.4]
  assign _T_234 = io_doneIn_1 | _T_232; // @[Controllers.scala 135:51:@573.4]
  assign _T_258 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@600.4]
  assign _T_260 = _T_258 & _T_174; // @[Controllers.scala 213:90:@602.4]
  assign _T_262 = ~ allDone; // @[Controllers.scala 213:132:@604.4]
  assign _T_263 = _T_260 & _T_262; // @[Controllers.scala 213:130:@605.4]
  assign _T_264 = ~ io_ctrDone; // @[Controllers.scala 213:156:@606.4]
  assign _T_266 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@609.4]
  assign _T_268 = _T_266 & _T_199; // @[Controllers.scala 213:90:@611.4]
  assign _T_274 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@617.4]
  assign _T_276 = _T_274 & _T_227; // @[Controllers.scala 213:90:@619.4]
  assign _T_283 = allDone == 1'h0; // @[package.scala 100:49:@625.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@654.4]
  assign io_ctrInc = io_doneIn_2; // @[Controllers.scala 122:17:@496.4]
  assign io_enableOut_0 = _T_263 & _T_264; // @[Controllers.scala 213:55:@608.4]
  assign io_enableOut_1 = _T_268 & _T_262; // @[Controllers.scala 213:55:@616.4]
  assign io_enableOut_2 = _T_276 & _T_262; // @[Controllers.scala 213:55:@624.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@595.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@597.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@599.4]
  assign active_0_clock = clock; // @[:@397.4]
  assign active_0_reset = reset; // @[:@398.4]
  assign active_0_io_input_set = _T_175 & _T_177; // @[Controllers.scala 128:30:@520.4]
  assign active_0_io_input_reset = _T_179 | allDone; // @[Controllers.scala 129:32:@525.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@418.4]
  assign active_1_clock = clock; // @[:@400.4]
  assign active_1_reset = reset; // @[:@401.4]
  assign active_1_io_input_set = _T_206 & _T_184; // @[Controllers.scala 135:32:@549.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_rst; // @[Controllers.scala 136:34:@553.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@419.4]
  assign active_2_clock = clock; // @[:@403.4]
  assign active_2_reset = reset; // @[:@404.4]
  assign active_2_io_input_set = _T_234 & _T_184; // @[Controllers.scala 135:32:@576.4]
  assign active_2_io_input_reset = io_doneIn_2 | io_rst; // @[Controllers.scala 136:34:@580.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@420.4]
  assign done_0_clock = clock; // @[:@406.4]
  assign done_0_reset = reset; // @[:@407.4]
  assign done_0_io_input_set = io_ctrDone & _T_196; // @[Controllers.scala 131:28:@539.4]
  assign done_0_io_input_reset = io_rst | allDone; // @[Controllers.scala 86:33:@432.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@421.4]
  assign done_1_clock = clock; // @[:@409.4]
  assign done_1_reset = reset; // @[:@410.4]
  assign done_1_io_input_set = io_ctrDone & _T_196; // @[Controllers.scala 138:30:@566.4]
  assign done_1_io_input_reset = io_rst | allDone; // @[Controllers.scala 86:33:@441.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@422.4]
  assign done_2_clock = clock; // @[:@412.4]
  assign done_2_reset = reset; // @[:@413.4]
  assign done_2_io_input_set = io_ctrDone & _T_196; // @[Controllers.scala 138:30:@593.4]
  assign done_2_io_input_reset = io_rst | allDone; // @[Controllers.scala 86:33:@450.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@423.4]
  assign iterDone_0_clock = clock; // @[:@453.4]
  assign iterDone_0_reset = reset; // @[:@454.4]
  assign iterDone_0_io_input_set = _T_185 & _T_193; // @[Controllers.scala 130:32:@535.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@472.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@461.4]
  assign iterDone_1_clock = clock; // @[:@456.4]
  assign iterDone_1_reset = reset; // @[:@457.4]
  assign iterDone_1_io_input_set = io_doneIn_1 & _T_184; // @[Controllers.scala 137:34:@562.4]
  assign iterDone_1_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@481.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@462.4]
  assign iterDone_2_clock = clock; // @[:@459.4]
  assign iterDone_2_reset = reset; // @[:@460.4]
  assign iterDone_2_io_input_set = io_doneIn_2 & _T_184; // @[Controllers.scala 137:34:@589.4]
  assign iterDone_2_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@490.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@463.4]
  assign RetimeWrapper_clock = clock; // @[:@498.4]
  assign RetimeWrapper_reset = reset; // @[:@499.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@501.4]
  assign RetimeWrapper_io_in = io_doneIn_2; // @[package.scala 94:16:@500.4]
  assign RetimeWrapper_1_clock = clock; // @[:@631.4]
  assign RetimeWrapper_1_reset = reset; // @[:@632.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@634.4]
  assign RetimeWrapper_1_io_in = allDone & _T_286; // @[package.scala 94:16:@633.4]
  assign RetimeWrapper_2_clock = clock; // @[:@648.4]
  assign RetimeWrapper_2_reset = reset; // @[:@649.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@651.4]
  assign RetimeWrapper_2_io_in = allDone & _T_300; // @[package.scala 94:16:@650.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_286 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_300 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_286 <= 1'h0;
    end else begin
      _T_286 <= _T_283;
    end
    if (reset) begin
      _T_300 <= 1'h0;
    end else begin
      _T_300 <= _T_283;
    end
  end
endmodule
module InstrumentationCounter( // @[:@705.2]
  input         clock, // @[:@706.4]
  input         reset, // @[:@707.4]
  input         io_enable, // @[:@708.4]
  output [63:0] io_count // @[:@708.4]
);
  reg [63:0] ff; // @[Counter.scala 223:19:@710.4]
  reg [63:0] _RAND_0;
  wire [64:0] _T_12; // @[Counter.scala 224:27:@711.4]
  wire [63:0] _T_13; // @[Counter.scala 224:27:@712.4]
  wire [63:0] _T_14; // @[Counter.scala 224:12:@713.4]
  assign _T_12 = ff + 64'h1; // @[Counter.scala 224:27:@711.4]
  assign _T_13 = ff + 64'h1; // @[Counter.scala 224:27:@712.4]
  assign _T_14 = io_enable ? _T_13 : ff; // @[Counter.scala 224:12:@713.4]
  assign io_count = ff; // @[Counter.scala 225:12:@715.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  ff = _RAND_0[63:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 64'h0;
    end else begin
      if (io_enable) begin
        ff <= _T_13;
      end
    end
  end
endmodule
module SRAM( // @[:@745.2]
  input         clock, // @[:@746.4]
  input  [8:0]  io_raddr, // @[:@748.4]
  input         io_wen, // @[:@748.4]
  input  [8:0]  io_waddr, // @[:@748.4]
  input  [31:0] io_wdata, // @[:@748.4]
  output [31:0] io_rdata, // @[:@748.4]
  input         io_backpressure // @[:@748.4]
);
  wire [31:0] SRAMVerilogSim_rdata; // @[SRAM.scala 187:23:@750.4]
  wire [31:0] SRAMVerilogSim_wdata; // @[SRAM.scala 187:23:@750.4]
  wire  SRAMVerilogSim_backpressure; // @[SRAM.scala 187:23:@750.4]
  wire  SRAMVerilogSim_wen; // @[SRAM.scala 187:23:@750.4]
  wire  SRAMVerilogSim_waddrEn; // @[SRAM.scala 187:23:@750.4]
  wire  SRAMVerilogSim_raddrEn; // @[SRAM.scala 187:23:@750.4]
  wire [8:0] SRAMVerilogSim_waddr; // @[SRAM.scala 187:23:@750.4]
  wire [8:0] SRAMVerilogSim_raddr; // @[SRAM.scala 187:23:@750.4]
  wire  SRAMVerilogSim_clk; // @[SRAM.scala 187:23:@750.4]
  SRAMVerilogSim #(.DWIDTH(32), .WORDS(300), .AWIDTH(9)) SRAMVerilogSim ( // @[SRAM.scala 187:23:@750.4]
    .rdata(SRAMVerilogSim_rdata),
    .wdata(SRAMVerilogSim_wdata),
    .backpressure(SRAMVerilogSim_backpressure),
    .wen(SRAMVerilogSim_wen),
    .waddrEn(SRAMVerilogSim_waddrEn),
    .raddrEn(SRAMVerilogSim_raddrEn),
    .waddr(SRAMVerilogSim_waddr),
    .raddr(SRAMVerilogSim_raddr),
    .clk(SRAMVerilogSim_clk)
  );
  assign io_rdata = SRAMVerilogSim_rdata; // @[SRAM.scala 197:16:@770.4]
  assign SRAMVerilogSim_wdata = io_wdata; // @[SRAM.scala 192:20:@764.4]
  assign SRAMVerilogSim_backpressure = io_backpressure; // @[SRAM.scala 193:27:@765.4]
  assign SRAMVerilogSim_wen = io_wen; // @[SRAM.scala 190:18:@762.4]
  assign SRAMVerilogSim_waddrEn = 1'h1; // @[SRAM.scala 195:22:@767.4]
  assign SRAMVerilogSim_raddrEn = 1'h1; // @[SRAM.scala 194:22:@766.4]
  assign SRAMVerilogSim_waddr = io_waddr; // @[SRAM.scala 191:20:@763.4]
  assign SRAMVerilogSim_raddr = io_raddr; // @[SRAM.scala 189:20:@761.4]
  assign SRAMVerilogSim_clk = clock; // @[SRAM.scala 188:18:@760.4]
endmodule
module RetimeWrapper_5( // @[:@784.2]
  input        clock, // @[:@785.4]
  input        reset, // @[:@786.4]
  input        io_flow, // @[:@787.4]
  input  [8:0] io_in, // @[:@787.4]
  output [8:0] io_out // @[:@787.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@789.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@789.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@789.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@789.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@789.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@789.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@789.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@802.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@801.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@800.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@799.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@798.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@796.4]
endmodule
module Mem1D( // @[:@804.2]
  input         clock, // @[:@805.4]
  input         reset, // @[:@806.4]
  input  [8:0]  io_r_ofs_0, // @[:@807.4]
  input         io_r_backpressure, // @[:@807.4]
  input  [8:0]  io_w_ofs_0, // @[:@807.4]
  input  [31:0] io_w_data_0, // @[:@807.4]
  input         io_w_en_0, // @[:@807.4]
  output [31:0] io_output // @[:@807.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 753:21:@811.4]
  wire [8:0] SRAM_io_raddr; // @[MemPrimitives.scala 753:21:@811.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 753:21:@811.4]
  wire [8:0] SRAM_io_waddr; // @[MemPrimitives.scala 753:21:@811.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 753:21:@811.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 753:21:@811.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 753:21:@811.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@814.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@814.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@814.4]
  wire [8:0] RetimeWrapper_io_in; // @[package.scala 93:22:@814.4]
  wire [8:0] RetimeWrapper_io_out; // @[package.scala 93:22:@814.4]
  wire  wInBound; // @[MemPrimitives.scala 740:32:@809.4]
  SRAM SRAM ( // @[MemPrimitives.scala 753:21:@811.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@814.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 9'h12c; // @[MemPrimitives.scala 740:32:@809.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 760:17:@827.4]
  assign SRAM_clock = clock; // @[:@812.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 754:37:@821.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 757:22:@824.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 756:22:@822.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 758:22:@825.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 759:30:@826.4]
  assign RetimeWrapper_clock = clock; // @[:@815.4]
  assign RetimeWrapper_reset = reset; // @[:@816.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@818.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@817.4]
endmodule
module StickySelects( // @[:@829.2]
  input   io_ins_0, // @[:@832.4]
  output  io_outs_0 // @[:@832.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@834.4]
endmodule
module RetimeWrapper_6( // @[:@848.2]
  input   clock, // @[:@849.4]
  input   reset, // @[:@850.4]
  input   io_flow, // @[:@851.4]
  input   io_in, // @[:@851.4]
  output  io_out // @[:@851.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@853.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@853.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@853.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@853.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@853.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@853.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@853.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@866.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@865.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@864.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@863.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@862.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@860.4]
endmodule
module x471_A_sram_0( // @[:@868.2]
  input         clock, // @[:@869.4]
  input         reset, // @[:@870.4]
  input  [8:0]  io_rPort_0_ofs_0, // @[:@871.4]
  input         io_rPort_0_en_0, // @[:@871.4]
  input         io_rPort_0_backpressure, // @[:@871.4]
  output [31:0] io_rPort_0_output_0, // @[:@871.4]
  input  [8:0]  io_wPort_0_ofs_0, // @[:@871.4]
  input  [31:0] io_wPort_0_data_0, // @[:@871.4]
  input         io_wPort_0_en_0 // @[:@871.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@886.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@886.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@886.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@886.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@886.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@886.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@886.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@886.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@912.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@912.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@926.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@926.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@926.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@926.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@926.4]
  wire [41:0] _T_70; // @[Cat.scala 30:58:@904.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@916.4]
  wire [10:0] _T_78; // @[Cat.scala 30:58:@918.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@886.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@912.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@926.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_70 = {io_wPort_0_en_0,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@904.4]
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@916.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@918.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@933.4]
  assign Mem1D_clock = clock; // @[:@887.4]
  assign Mem1D_reset = reset; // @[:@888.4]
  assign Mem1D_io_r_ofs_0 = _T_78[8:0]; // @[MemPrimitives.scala 131:28:@922.4]
  assign Mem1D_io_r_backpressure = _T_78[9]; // @[MemPrimitives.scala 132:32:@923.4]
  assign Mem1D_io_w_ofs_0 = _T_70[8:0]; // @[MemPrimitives.scala 94:28:@908.4]
  assign Mem1D_io_w_data_0 = _T_70[40:9]; // @[MemPrimitives.scala 95:29:@909.4]
  assign Mem1D_io_w_en_0 = _T_70[41]; // @[MemPrimitives.scala 96:27:@910.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@915.4]
  assign RetimeWrapper_clock = clock; // @[:@927.4]
  assign RetimeWrapper_reset = reset; // @[:@928.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@930.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@929.4]
endmodule
module x538_outr_UnitPipe_DenseTransfer_sm( // @[:@1681.2]
  input   clock, // @[:@1682.4]
  input   reset, // @[:@1683.4]
  input   io_enable, // @[:@1684.4]
  output  io_done, // @[:@1684.4]
  input   io_parentAck, // @[:@1684.4]
  input   io_doneIn_0, // @[:@1684.4]
  input   io_doneIn_1, // @[:@1684.4]
  output  io_enableOut_0, // @[:@1684.4]
  output  io_enableOut_1, // @[:@1684.4]
  output  io_childAck_0, // @[:@1684.4]
  output  io_childAck_1, // @[:@1684.4]
  input   io_ctrCopyDone_0, // @[:@1684.4]
  input   io_ctrCopyDone_1 // @[:@1684.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1687.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1687.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1687.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1687.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1687.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1687.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1690.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1690.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1690.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1690.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1690.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1690.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1693.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1693.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1693.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1693.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1693.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1693.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1696.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1696.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1696.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1696.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1696.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1696.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1725.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1725.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1725.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1725.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1725.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1725.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1728.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1728.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1728.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1728.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1728.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1728.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1769.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1769.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1769.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1769.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1769.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1783.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1783.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1783.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1783.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1783.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1801.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1801.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1801.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1801.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1801.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1838.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1838.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1838.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1838.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1838.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1852.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1852.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1852.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1852.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1852.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1870.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1870.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1870.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1870.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1870.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1917.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1917.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1917.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1917.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1917.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1934.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1934.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1934.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1934.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1934.4]
  wire  allDone; // @[Controllers.scala 80:47:@1699.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1753.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1754.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1755.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1756.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1757.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1760.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1762.4]
  wire  _T_148; // @[package.scala 96:25:@1774.4 package.scala 96:25:@1775.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1777.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1778.4]
  wire  _T_160; // @[package.scala 96:25:@1788.4 package.scala 96:25:@1789.4]
  wire  _T_178; // @[package.scala 96:25:@1806.4 package.scala 96:25:@1807.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1809.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1810.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1822.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1823.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1824.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1825.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1826.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1829.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1831.4]
  wire  _T_216; // @[package.scala 96:25:@1843.4 package.scala 96:25:@1844.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1846.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1847.4]
  wire  _T_228; // @[package.scala 96:25:@1857.4 package.scala 96:25:@1858.4]
  wire  _T_246; // @[package.scala 96:25:@1875.4 package.scala 96:25:@1876.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1878.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1879.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1895.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1897.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1899.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1904.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1906.4]
  wire  _T_282; // @[package.scala 100:49:@1912.4]
  reg  _T_285; // @[package.scala 48:56:@1913.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1915.4]
  reg  _T_299; // @[package.scala 48:56:@1931.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1687.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1690.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1693.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1696.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1725.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1728.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1769.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1783.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1801.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1838.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1852.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1870.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1917.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1934.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1699.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1753.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1754.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1755.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1756.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1757.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1760.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1762.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1774.4 package.scala 96:25:@1775.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1777.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1778.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1788.4 package.scala 96:25:@1789.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1806.4 package.scala 96:25:@1807.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1809.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1810.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1822.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1823.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1824.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1825.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1826.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1829.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1831.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1843.4 package.scala 96:25:@1844.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1846.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1847.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1857.4 package.scala 96:25:@1858.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1875.4 package.scala 96:25:@1876.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1878.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1879.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1895.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1897.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1899.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1904.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1906.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1912.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1915.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1941.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1903.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1911.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1892.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1894.4]
  assign active_0_clock = clock; // @[:@1688.4]
  assign active_0_reset = reset; // @[:@1689.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1764.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1768.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1702.4]
  assign active_1_clock = clock; // @[:@1691.4]
  assign active_1_reset = reset; // @[:@1692.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1833.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1837.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1703.4]
  assign done_0_clock = clock; // @[:@1694.4]
  assign done_0_reset = reset; // @[:@1695.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1814.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1714.4 Controllers.scala 170:32:@1821.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1704.4]
  assign done_1_clock = clock; // @[:@1697.4]
  assign done_1_reset = reset; // @[:@1698.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1883.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1723.4 Controllers.scala 170:32:@1890.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1705.4]
  assign iterDone_0_clock = clock; // @[:@1726.4]
  assign iterDone_0_reset = reset; // @[:@1727.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1782.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1741.4 Controllers.scala 168:36:@1798.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1731.4]
  assign iterDone_1_clock = clock; // @[:@1729.4]
  assign iterDone_1_reset = reset; // @[:@1730.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1851.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1750.4 Controllers.scala 168:36:@1867.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1732.4]
  assign RetimeWrapper_clock = clock; // @[:@1770.4]
  assign RetimeWrapper_reset = reset; // @[:@1771.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1773.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1772.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1784.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1785.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1787.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1786.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1802.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1803.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1805.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1804.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1839.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1840.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1842.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1841.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1853.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1854.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1856.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1855.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1871.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1872.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1874.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1873.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1918.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1919.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1921.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1920.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1935.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1936.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1938.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1937.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module FF_1( // @[:@2048.2]
  input        clock, // @[:@2049.4]
  input        reset, // @[:@2050.4]
  output [6:0] io_rPort_0_output_0, // @[:@2051.4]
  input  [6:0] io_wPort_0_data_0, // @[:@2051.4]
  input        io_wPort_0_reset, // @[:@2051.4]
  input  [6:0] io_wPort_0_init, // @[:@2051.4]
  input        io_wPort_0_en_0, // @[:@2051.4]
  input        io_reset // @[:@2051.4]
);
  reg [6:0] ff; // @[MemPrimitives.scala 321:19:@2066.4]
  reg [31:0] _RAND_0;
  wire  anyReset; // @[MemPrimitives.scala 322:65:@2067.4]
  wire [6:0] _T_68; // @[MemPrimitives.scala 325:32:@2068.4]
  wire [6:0] _T_69; // @[MemPrimitives.scala 325:12:@2069.4]
  assign anyReset = io_wPort_0_reset | io_reset; // @[MemPrimitives.scala 322:65:@2067.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@2068.4]
  assign _T_69 = anyReset ? io_wPort_0_init : _T_68; // @[MemPrimitives.scala 325:12:@2069.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@2071.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= io_wPort_0_init;
    end else begin
      if (anyReset) begin
        ff <= io_wPort_0_init;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module CompactingCounter( // @[:@2073.2]
  input        clock, // @[:@2074.4]
  input        reset, // @[:@2075.4]
  input        io_input_reset, // @[:@2076.4]
  input        io_input_enables_0, // @[:@2076.4]
  output [6:0] io_output_count // @[:@2076.4]
);
  wire  base_clock; // @[Counter.scala 200:20:@2078.4]
  wire  base_reset; // @[Counter.scala 200:20:@2078.4]
  wire [6:0] base_io_rPort_0_output_0; // @[Counter.scala 200:20:@2078.4]
  wire [6:0] base_io_wPort_0_data_0; // @[Counter.scala 200:20:@2078.4]
  wire  base_io_wPort_0_reset; // @[Counter.scala 200:20:@2078.4]
  wire [6:0] base_io_wPort_0_init; // @[Counter.scala 200:20:@2078.4]
  wire  base_io_wPort_0_en_0; // @[Counter.scala 200:20:@2078.4]
  wire  base_io_reset; // @[Counter.scala 200:20:@2078.4]
  wire [6:0] count; // @[Counter.scala 206:42:@2097.4]
  wire [6:0] num_enabled; // @[Counter.scala 207:56:@2098.4]
  wire [7:0] _T_27; // @[Counter.scala 208:22:@2103.4]
  wire [6:0] _T_28; // @[Counter.scala 208:22:@2104.4]
  wire [6:0] newval; // @[Counter.scala 208:22:@2105.4]
  wire  isMax; // @[Counter.scala 209:40:@2106.4]
  wire [7:0] _T_34; // @[Counter.scala 210:32:@2109.4]
  wire [6:0] _T_35; // @[Counter.scala 210:32:@2110.4]
  wire [6:0] _T_36; // @[Counter.scala 210:32:@2111.4]
  wire [6:0] next; // @[Counter.scala 210:17:@2112.4]
  wire [6:0] _T_38; // @[Counter.scala 211:68:@2113.4]
  FF_1 base ( // @[Counter.scala 200:20:@2078.4]
    .clock(base_clock),
    .reset(base_reset),
    .io_rPort_0_output_0(base_io_rPort_0_output_0),
    .io_wPort_0_data_0(base_io_wPort_0_data_0),
    .io_wPort_0_reset(base_io_wPort_0_reset),
    .io_wPort_0_init(base_io_wPort_0_init),
    .io_wPort_0_en_0(base_io_wPort_0_en_0),
    .io_reset(base_io_reset)
  );
  assign count = $signed(base_io_rPort_0_output_0); // @[Counter.scala 206:42:@2097.4]
  assign num_enabled = io_input_enables_0 ? $signed(7'sh1) : $signed(7'sh0); // @[Counter.scala 207:56:@2098.4]
  assign _T_27 = $signed(count) + $signed(num_enabled); // @[Counter.scala 208:22:@2103.4]
  assign _T_28 = $signed(count) + $signed(num_enabled); // @[Counter.scala 208:22:@2104.4]
  assign newval = $signed(_T_28); // @[Counter.scala 208:22:@2105.4]
  assign isMax = $signed(newval) >= $signed(7'sh10); // @[Counter.scala 209:40:@2106.4]
  assign _T_34 = $signed(newval) - $signed(7'sh10); // @[Counter.scala 210:32:@2109.4]
  assign _T_35 = $signed(newval) - $signed(7'sh10); // @[Counter.scala 210:32:@2110.4]
  assign _T_36 = $signed(_T_35); // @[Counter.scala 210:32:@2111.4]
  assign next = isMax ? $signed(_T_36) : $signed(newval); // @[Counter.scala 210:17:@2112.4]
  assign _T_38 = $unsigned(next); // @[Counter.scala 211:68:@2113.4]
  assign io_output_count = $signed(base_io_rPort_0_output_0); // @[Counter.scala 213:19:@2117.4]
  assign base_clock = clock; // @[:@2079.4]
  assign base_reset = reset; // @[:@2080.4]
  assign base_io_wPort_0_data_0 = io_input_reset ? 7'h0 : _T_38; // @[Counter.scala 211:30:@2115.4]
  assign base_io_wPort_0_reset = io_input_reset; // @[Counter.scala 203:26:@2095.4]
  assign base_io_wPort_0_init = 7'h0; // @[Counter.scala 202:25:@2094.4]
  assign base_io_wPort_0_en_0 = io_input_enables_0; // @[Counter.scala 204:28:@2096.4]
  assign base_io_reset = 1'h0;
endmodule
module CompactingIncDincCtr( // @[:@2194.2]
  input   clock, // @[:@2195.4]
  input   reset, // @[:@2196.4]
  input   io_input_inc_en_0, // @[:@2197.4]
  input   io_input_dinc_en_0, // @[:@2197.4]
  output  io_output_empty, // @[:@2197.4]
  output  io_output_full // @[:@2197.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@2199.4]
  reg [31:0] _RAND_0;
  wire [6:0] numPushed; // @[Counter.scala 172:47:@2200.4]
  wire [6:0] numPopped; // @[Counter.scala 173:48:@2201.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@2202.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@2202.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@2203.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@2204.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@2205.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@2205.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@2206.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@2207.4]
  assign numPushed = io_input_inc_en_0 ? $signed(7'sh1) : $signed(7'sh0); // @[Counter.scala 172:47:@2200.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(7'sh1) : $signed(7'sh0); // @[Counter.scala 173:48:@2201.4]
  assign _GEN_0 = {{25{numPushed[6]}},numPushed}; // @[Counter.scala 174:14:@2202.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@2202.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@2203.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@2204.4]
  assign _GEN_1 = {{25{numPopped[6]}},numPopped}; // @[Counter.scala 174:26:@2205.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@2205.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@2206.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@2207.4]
  assign io_output_empty = $signed(cnt) < $signed(32'sh1); // @[Counter.scala 179:19:@2214.4]
  assign io_output_full = $signed(cnt) > $signed(32'shf); // @[Counter.scala 181:18:@2221.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module Mem1D_3( // @[:@2229.2]
  input         clock, // @[:@2230.4]
  input  [4:0]  io_r_ofs_0, // @[:@2232.4]
  input  [4:0]  io_w_ofs_0, // @[:@2232.4]
  input  [95:0] io_w_data_0, // @[:@2232.4]
  input         io_w_en_0, // @[:@2232.4]
  output [95:0] io_output // @[:@2232.4]
);
  reg [95:0] _T_127 [0:15]; // @[MemPrimitives.scala 771:18:@2236.4]
  reg [95:0] _RAND_0;
  wire [95:0] _T_127__T_132_data; // @[MemPrimitives.scala 771:18:@2236.4]
  wire [3:0] _T_127__T_132_addr; // @[MemPrimitives.scala 771:18:@2236.4]
  wire [95:0] _T_127__T_130_data; // @[MemPrimitives.scala 771:18:@2236.4]
  wire [3:0] _T_127__T_130_addr; // @[MemPrimitives.scala 771:18:@2236.4]
  wire  _T_127__T_130_mask; // @[MemPrimitives.scala 771:18:@2236.4]
  wire  _T_127__T_130_en; // @[MemPrimitives.scala 771:18:@2236.4]
  wire  wInBound; // @[MemPrimitives.scala 740:32:@2234.4]
  assign _T_127__T_132_addr = io_r_ofs_0[3:0];
  assign _T_127__T_132_data = _T_127[_T_127__T_132_addr]; // @[MemPrimitives.scala 771:18:@2236.4]
  assign _T_127__T_130_data = io_w_data_0;
  assign _T_127__T_130_addr = io_w_ofs_0[3:0];
  assign _T_127__T_130_mask = 1'h1;
  assign _T_127__T_130_en = io_w_en_0 & wInBound;
  assign wInBound = io_w_ofs_0 <= 5'h10; // @[MemPrimitives.scala 740:32:@2234.4]
  assign io_output = _T_127__T_132_data; // @[MemPrimitives.scala 773:17:@2245.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {3{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    _T_127[initvar] = _RAND_0[95:0];
  `endif // RANDOMIZE_MEM_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T_127__T_130_en & _T_127__T_130_mask) begin
      _T_127[_T_127__T_130_addr] <= _T_127__T_130_data; // @[MemPrimitives.scala 771:18:@2236.4]
    end
  end
endmodule
module Compactor( // @[:@2247.2]
  input  [95:0] io_in_0_data, // @[:@2250.4]
  output [95:0] io_out_0_data // @[:@2250.4]
);
  assign io_out_0_data = io_in_0_data; // @[MemPrimitives.scala 848:22:@2254.4]
endmodule
module CompactingEnqNetwork( // @[:@2258.2]
  input  [6:0]  io_headCnt, // @[:@2261.4]
  input  [95:0] io_in_0_data, // @[:@2261.4]
  input         io_in_0_en, // @[:@2261.4]
  output [95:0] io_out_0_data, // @[:@2261.4]
  output        io_out_0_en // @[:@2261.4]
);
  wire [95:0] compactor_io_in_0_data; // @[MemPrimitives.scala 870:25:@2264.4]
  wire [95:0] compactor_io_out_0_data; // @[MemPrimitives.scala 870:25:@2264.4]
  wire [6:0] numEnabled; // @[MemPrimitives.scala 866:38:@2263.4]
  wire [6:0] _GEN_0; // @[Math.scala 53:59:@2270.4]
  wire [6:0] current_base_bank; // @[Math.scala 53:59:@2270.4]
  wire [6:0] _T_22; // @[MemPrimitives.scala 876:46:@2271.4]
  wire [7:0] _T_23; // @[MemPrimitives.scala 876:33:@2272.4]
  wire [6:0] _T_24; // @[MemPrimitives.scala 876:33:@2273.4]
  wire [6:0] _T_25; // @[MemPrimitives.scala 876:33:@2274.4]
  wire [7:0] _T_27; // @[MemPrimitives.scala 876:53:@2275.4]
  wire [6:0] _T_28; // @[MemPrimitives.scala 876:53:@2276.4]
  wire [6:0] upper; // @[MemPrimitives.scala 876:53:@2277.4]
  wire  _T_30; // @[MemPrimitives.scala 877:34:@2278.4]
  wire [6:0] num_straddling; // @[MemPrimitives.scala 877:27:@2279.4]
  wire [7:0] _T_33; // @[MemPrimitives.scala 878:40:@2281.4]
  wire [6:0] _T_34; // @[MemPrimitives.scala 878:40:@2282.4]
  wire [6:0] num_straight; // @[MemPrimitives.scala 878:40:@2283.4]
  wire  _T_36; // @[MemPrimitives.scala 880:40:@2284.4]
  wire  _T_38; // @[MemPrimitives.scala 880:73:@2285.4]
  wire  _T_44; // @[MemPrimitives.scala 880:109:@2290.4]
  wire  _T_45; // @[MemPrimitives.scala 880:94:@2291.4]
  wire [7:0] _T_53; // @[MemPrimitives.scala 881:72:@2295.4]
  wire [6:0] _T_54; // @[MemPrimitives.scala 881:72:@2296.4]
  wire [6:0] _T_55; // @[MemPrimitives.scala 881:72:@2297.4]
  wire [7:0] _T_57; // @[MemPrimitives.scala 881:101:@2298.4]
  wire [6:0] _T_58; // @[MemPrimitives.scala 881:101:@2299.4]
  wire [6:0] _T_59; // @[MemPrimitives.scala 881:101:@2300.4]
  wire [6:0] _T_60; // @[MemPrimitives.scala 881:27:@2301.4]
  wire [6:0] _T_62; // @[MemPrimitives.scala 885:57:@2302.4]
  wire  _T_64; // @[Mux.scala 46:19:@2303.4]
  Compactor compactor ( // @[MemPrimitives.scala 870:25:@2264.4]
    .io_in_0_data(compactor_io_in_0_data),
    .io_out_0_data(compactor_io_out_0_data)
  );
  assign numEnabled = io_in_0_en ? 7'h1 : 7'h0; // @[MemPrimitives.scala 866:38:@2263.4]
  assign _GEN_0 = $signed(io_headCnt) % $signed(7'sh1); // @[Math.scala 53:59:@2270.4]
  assign current_base_bank = _GEN_0[6:0]; // @[Math.scala 53:59:@2270.4]
  assign _T_22 = $signed(numEnabled); // @[MemPrimitives.scala 876:46:@2271.4]
  assign _T_23 = $signed(current_base_bank) + $signed(_T_22); // @[MemPrimitives.scala 876:33:@2272.4]
  assign _T_24 = $signed(current_base_bank) + $signed(_T_22); // @[MemPrimitives.scala 876:33:@2273.4]
  assign _T_25 = $signed(_T_24); // @[MemPrimitives.scala 876:33:@2274.4]
  assign _T_27 = $signed(_T_25) - $signed(7'sh1); // @[MemPrimitives.scala 876:53:@2275.4]
  assign _T_28 = $signed(_T_25) - $signed(7'sh1); // @[MemPrimitives.scala 876:53:@2276.4]
  assign upper = $signed(_T_28); // @[MemPrimitives.scala 876:53:@2277.4]
  assign _T_30 = $signed(upper) < $signed(7'sh0); // @[MemPrimitives.scala 877:34:@2278.4]
  assign num_straddling = _T_30 ? $signed(7'sh0) : $signed(upper); // @[MemPrimitives.scala 877:27:@2279.4]
  assign _T_33 = $signed(_T_22) - $signed(num_straddling); // @[MemPrimitives.scala 878:40:@2281.4]
  assign _T_34 = $signed(_T_22) - $signed(num_straddling); // @[MemPrimitives.scala 878:40:@2282.4]
  assign num_straight = $signed(_T_34); // @[MemPrimitives.scala 878:40:@2283.4]
  assign _T_36 = $signed(7'sh0) < $signed(num_straddling); // @[MemPrimitives.scala 880:40:@2284.4]
  assign _T_38 = $signed(7'sh0) >= $signed(current_base_bank); // @[MemPrimitives.scala 880:73:@2285.4]
  assign _T_44 = $signed(7'sh0) < $signed(_T_25); // @[MemPrimitives.scala 880:109:@2290.4]
  assign _T_45 = _T_38 & _T_44; // @[MemPrimitives.scala 880:94:@2291.4]
  assign _T_53 = {{1{num_straight[6]}},num_straight}; // @[MemPrimitives.scala 881:72:@2295.4]
  assign _T_54 = _T_53[6:0]; // @[MemPrimitives.scala 881:72:@2296.4]
  assign _T_55 = $signed(_T_54); // @[MemPrimitives.scala 881:72:@2297.4]
  assign _T_57 = $signed(7'sh0) - $signed(current_base_bank); // @[MemPrimitives.scala 881:101:@2298.4]
  assign _T_58 = $signed(7'sh0) - $signed(current_base_bank); // @[MemPrimitives.scala 881:101:@2299.4]
  assign _T_59 = $signed(_T_58); // @[MemPrimitives.scala 881:101:@2300.4]
  assign _T_60 = _T_36 ? $signed(_T_55) : $signed(_T_59); // @[MemPrimitives.scala 881:27:@2301.4]
  assign _T_62 = $unsigned(_T_60); // @[MemPrimitives.scala 885:57:@2302.4]
  assign _T_64 = 7'h0 == _T_62; // @[Mux.scala 46:19:@2303.4]
  assign io_out_0_data = _T_64 ? compactor_io_out_0_data : 96'h0; // @[MemPrimitives.scala 890:63:@2305.4]
  assign io_out_0_en = _T_36 | _T_45; // @[MemPrimitives.scala 891:63:@2306.4]
  assign compactor_io_in_0_data = io_in_0_data; // @[MemPrimitives.scala 871:19:@2268.4]
endmodule
module CompactingDeqNetwork( // @[:@2308.2]
  input  [6:0]  io_tailCnt, // @[:@2311.4]
  input  [95:0] io_input_data_0, // @[:@2311.4]
  output [95:0] io_output_0 // @[:@2311.4]
);
  wire [6:0] _GEN_0; // @[Math.scala 53:59:@2315.4]
  wire [6:0] current_base_bank; // @[Math.scala 53:59:@2315.4]
  wire [6:0] _T_55; // @[MemPrimitives.scala 917:64:@2338.4]
  wire [7:0] _T_56; // @[MemPrimitives.scala 917:71:@2339.4]
  wire [6:0] _T_57; // @[MemPrimitives.scala 917:71:@2340.4]
  wire [6:0] _GEN_1; // @[Math.scala 55:59:@2341.4]
  wire [6:0] _T_59; // @[Math.scala 55:59:@2341.4]
  wire  _T_62; // @[Mux.scala 46:19:@2342.4]
  assign _GEN_0 = $signed(io_tailCnt) % $signed(7'sh1); // @[Math.scala 53:59:@2315.4]
  assign current_base_bank = _GEN_0[6:0]; // @[Math.scala 53:59:@2315.4]
  assign _T_55 = $unsigned(current_base_bank); // @[MemPrimitives.scala 917:64:@2338.4]
  assign _T_56 = {{1'd0}, _T_55}; // @[MemPrimitives.scala 917:71:@2339.4]
  assign _T_57 = _T_56[6:0]; // @[MemPrimitives.scala 917:71:@2340.4]
  assign _GEN_1 = _T_57 % 7'h1; // @[Math.scala 55:59:@2341.4]
  assign _T_59 = _GEN_1[6:0]; // @[Math.scala 55:59:@2341.4]
  assign _T_62 = 7'h0 == _T_59; // @[Mux.scala 46:19:@2342.4]
  assign io_output_0 = _T_62 ? io_input_data_0 : 96'h0; // @[MemPrimitives.scala 921:18:@2344.4]
endmodule
module x475_fifo( // @[:@2346.2]
  input         clock, // @[:@2347.4]
  input         reset, // @[:@2348.4]
  input         io_rPort_0_en_0, // @[:@2349.4]
  output [95:0] io_rPort_0_output_0, // @[:@2349.4]
  input  [95:0] io_wPort_0_data_0, // @[:@2349.4]
  input         io_wPort_0_en_0, // @[:@2349.4]
  output        io_full, // @[:@2349.4]
  output        io_empty, // @[:@2349.4]
  input         io_active_0_in, // @[:@2349.4]
  output        io_active_0_out // @[:@2349.4]
);
  wire  headCtr_clock; // @[MemPrimitives.scala 381:23:@2373.4]
  wire  headCtr_reset; // @[MemPrimitives.scala 381:23:@2373.4]
  wire  headCtr_io_input_reset; // @[MemPrimitives.scala 381:23:@2373.4]
  wire  headCtr_io_input_enables_0; // @[MemPrimitives.scala 381:23:@2373.4]
  wire [6:0] headCtr_io_output_count; // @[MemPrimitives.scala 381:23:@2373.4]
  wire  tailCtr_clock; // @[MemPrimitives.scala 382:23:@2381.4]
  wire  tailCtr_reset; // @[MemPrimitives.scala 382:23:@2381.4]
  wire  tailCtr_io_input_reset; // @[MemPrimitives.scala 382:23:@2381.4]
  wire  tailCtr_io_input_enables_0; // @[MemPrimitives.scala 382:23:@2381.4]
  wire [6:0] tailCtr_io_output_count; // @[MemPrimitives.scala 382:23:@2381.4]
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2395.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2395.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2395.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2395.4]
  wire  elements_io_output_empty; // @[MemPrimitives.scala 392:24:@2395.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2395.4]
  wire  m_0_clock; // @[MemPrimitives.scala 398:56:@2409.4]
  wire [4:0] m_0_io_r_ofs_0; // @[MemPrimitives.scala 398:56:@2409.4]
  wire [4:0] m_0_io_w_ofs_0; // @[MemPrimitives.scala 398:56:@2409.4]
  wire [95:0] m_0_io_w_data_0; // @[MemPrimitives.scala 398:56:@2409.4]
  wire  m_0_io_w_en_0; // @[MemPrimitives.scala 398:56:@2409.4]
  wire [95:0] m_0_io_output; // @[MemPrimitives.scala 398:56:@2409.4]
  wire [6:0] enqCompactor_io_headCnt; // @[MemPrimitives.scala 402:28:@2425.4]
  wire [95:0] enqCompactor_io_in_0_data; // @[MemPrimitives.scala 402:28:@2425.4]
  wire  enqCompactor_io_in_0_en; // @[MemPrimitives.scala 402:28:@2425.4]
  wire [95:0] enqCompactor_io_out_0_data; // @[MemPrimitives.scala 402:28:@2425.4]
  wire  enqCompactor_io_out_0_en; // @[MemPrimitives.scala 402:28:@2425.4]
  wire [6:0] deqCompactor_io_tailCnt; // @[MemPrimitives.scala 421:28:@2447.4]
  wire [95:0] deqCompactor_io_input_data_0; // @[MemPrimitives.scala 421:28:@2447.4]
  wire [95:0] deqCompactor_io_output_0; // @[MemPrimitives.scala 421:28:@2447.4]
  wire [6:0] _GEN_0; // @[Math.scala 53:59:@2436.4]
  wire [6:0] active_w_bank; // @[Math.scala 53:59:@2436.4]
  wire [7:0] active_w_addr; // @[Math.scala 52:59:@2437.4]
  wire  _T_102; // @[MemPrimitives.scala 414:38:@2438.4]
  wire [8:0] _T_104; // @[MemPrimitives.scala 414:69:@2439.4]
  wire [7:0] _T_105; // @[MemPrimitives.scala 414:69:@2440.4]
  wire [7:0] _T_106; // @[MemPrimitives.scala 414:69:@2441.4]
  wire [7:0] _T_107; // @[MemPrimitives.scala 414:19:@2442.4]
  wire [7:0] _T_108; // @[MemPrimitives.scala 415:32:@2443.4]
  wire [6:0] _GEN_1; // @[Math.scala 53:59:@2455.4]
  wire [6:0] active_r_bank; // @[Math.scala 53:59:@2455.4]
  wire [7:0] active_r_addr; // @[Math.scala 52:59:@2456.4]
  wire  _T_112; // @[MemPrimitives.scala 427:38:@2457.4]
  wire [8:0] _T_114; // @[MemPrimitives.scala 427:69:@2458.4]
  wire [7:0] _T_115; // @[MemPrimitives.scala 427:69:@2459.4]
  wire [7:0] _T_116; // @[MemPrimitives.scala 427:69:@2460.4]
  wire [7:0] _T_117; // @[MemPrimitives.scala 427:19:@2461.4]
  wire [7:0] _T_118; // @[MemPrimitives.scala 428:32:@2462.4]
  CompactingCounter headCtr ( // @[MemPrimitives.scala 381:23:@2373.4]
    .clock(headCtr_clock),
    .reset(headCtr_reset),
    .io_input_reset(headCtr_io_input_reset),
    .io_input_enables_0(headCtr_io_input_enables_0),
    .io_output_count(headCtr_io_output_count)
  );
  CompactingCounter tailCtr ( // @[MemPrimitives.scala 382:23:@2381.4]
    .clock(tailCtr_clock),
    .reset(tailCtr_reset),
    .io_input_reset(tailCtr_io_input_reset),
    .io_input_enables_0(tailCtr_io_input_enables_0),
    .io_output_count(tailCtr_io_output_count)
  );
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2395.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_empty(elements_io_output_empty),
    .io_output_full(elements_io_output_full)
  );
  Mem1D_3 m_0 ( // @[MemPrimitives.scala 398:56:@2409.4]
    .clock(m_0_clock),
    .io_r_ofs_0(m_0_io_r_ofs_0),
    .io_w_ofs_0(m_0_io_w_ofs_0),
    .io_w_data_0(m_0_io_w_data_0),
    .io_w_en_0(m_0_io_w_en_0),
    .io_output(m_0_io_output)
  );
  CompactingEnqNetwork enqCompactor ( // @[MemPrimitives.scala 402:28:@2425.4]
    .io_headCnt(enqCompactor_io_headCnt),
    .io_in_0_data(enqCompactor_io_in_0_data),
    .io_in_0_en(enqCompactor_io_in_0_en),
    .io_out_0_data(enqCompactor_io_out_0_data),
    .io_out_0_en(enqCompactor_io_out_0_en)
  );
  CompactingDeqNetwork deqCompactor ( // @[MemPrimitives.scala 421:28:@2447.4]
    .io_tailCnt(deqCompactor_io_tailCnt),
    .io_input_data_0(deqCompactor_io_input_data_0),
    .io_output_0(deqCompactor_io_output_0)
  );
  assign _GEN_0 = $signed(headCtr_io_output_count) % $signed(7'sh1); // @[Math.scala 53:59:@2436.4]
  assign active_w_bank = _GEN_0[6:0]; // @[Math.scala 53:59:@2436.4]
  assign active_w_addr = $signed(headCtr_io_output_count) / $signed(7'sh1); // @[Math.scala 52:59:@2437.4]
  assign _T_102 = $signed(7'sh0) < $signed(active_w_bank); // @[MemPrimitives.scala 414:38:@2438.4]
  assign _T_104 = $signed(active_w_addr) + $signed(8'sh1); // @[MemPrimitives.scala 414:69:@2439.4]
  assign _T_105 = $signed(active_w_addr) + $signed(8'sh1); // @[MemPrimitives.scala 414:69:@2440.4]
  assign _T_106 = $signed(_T_105); // @[MemPrimitives.scala 414:69:@2441.4]
  assign _T_107 = _T_102 ? $signed(_T_106) : $signed(active_w_addr); // @[MemPrimitives.scala 414:19:@2442.4]
  assign _T_108 = $unsigned(_T_107); // @[MemPrimitives.scala 415:32:@2443.4]
  assign _GEN_1 = $signed(tailCtr_io_output_count) % $signed(7'sh1); // @[Math.scala 53:59:@2455.4]
  assign active_r_bank = _GEN_1[6:0]; // @[Math.scala 53:59:@2455.4]
  assign active_r_addr = $signed(tailCtr_io_output_count) / $signed(7'sh1); // @[Math.scala 52:59:@2456.4]
  assign _T_112 = $signed(7'sh0) < $signed(active_r_bank); // @[MemPrimitives.scala 427:38:@2457.4]
  assign _T_114 = $signed(active_r_addr) + $signed(8'sh1); // @[MemPrimitives.scala 427:69:@2458.4]
  assign _T_115 = $signed(active_r_addr) + $signed(8'sh1); // @[MemPrimitives.scala 427:69:@2459.4]
  assign _T_116 = $signed(_T_115); // @[MemPrimitives.scala 427:69:@2460.4]
  assign _T_117 = _T_112 ? $signed(_T_116) : $signed(active_r_addr); // @[MemPrimitives.scala 427:19:@2461.4]
  assign _T_118 = $unsigned(_T_117); // @[MemPrimitives.scala 428:32:@2462.4]
  assign io_rPort_0_output_0 = deqCompactor_io_output_0; // @[MemPrimitives.scala 432:82:@2466.4]
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 439:39:@2470.4]
  assign io_empty = elements_io_output_empty; // @[MemPrimitives.scala 438:40:@2469.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 437:129:@2467.4]
  assign headCtr_clock = clock; // @[:@2374.4]
  assign headCtr_reset = reset; // @[:@2375.4]
  assign headCtr_io_input_reset = reset; // @[MemPrimitives.scala 385:26:@2391.4]
  assign headCtr_io_input_enables_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 383:129:@2389.4]
  assign tailCtr_clock = clock; // @[:@2382.4]
  assign tailCtr_reset = reset; // @[:@2383.4]
  assign tailCtr_io_input_reset = reset; // @[MemPrimitives.scala 386:26:@2392.4]
  assign tailCtr_io_input_enables_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 384:129:@2390.4]
  assign elements_clock = clock; // @[:@2396.4]
  assign elements_reset = reset; // @[:@2397.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 394:79:@2407.4]
  assign elements_io_input_dinc_en_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 395:80:@2408.4]
  assign m_0_clock = clock; // @[:@2410.4]
  assign m_0_io_r_ofs_0 = _T_118[4:0]; // @[MemPrimitives.scala 428:24:@2463.4]
  assign m_0_io_w_ofs_0 = _T_108[4:0]; // @[MemPrimitives.scala 415:24:@2444.4]
  assign m_0_io_w_data_0 = enqCompactor_io_out_0_data; // @[MemPrimitives.scala 416:25:@2445.4]
  assign m_0_io_w_en_0 = enqCompactor_io_out_0_en; // @[MemPrimitives.scala 417:25:@2446.4]
  assign enqCompactor_io_headCnt = headCtr_io_output_count; // @[MemPrimitives.scala 404:27:@2433.4]
  assign enqCompactor_io_in_0_data = io_wPort_0_data_0; // @[MemPrimitives.scala 406:90:@2434.4]
  assign enqCompactor_io_in_0_en = io_wPort_0_en_0; // @[MemPrimitives.scala 407:85:@2435.4]
  assign deqCompactor_io_tailCnt = tailCtr_io_output_count; // @[MemPrimitives.scala 423:27:@2454.4]
  assign deqCompactor_io_input_data_0 = m_0_io_output; // @[MemPrimitives.scala 429:35:@2464.4]
endmodule
module FF_3( // @[:@2476.2]
  input        clock, // @[:@2477.4]
  input        reset, // @[:@2478.4]
  output [8:0] io_rPort_0_output_0, // @[:@2479.4]
  input  [8:0] io_wPort_0_data_0, // @[:@2479.4]
  input        io_wPort_0_reset, // @[:@2479.4]
  input        io_wPort_0_en_0 // @[:@2479.4]
);
  reg [8:0] ff; // @[MemPrimitives.scala 321:19:@2494.4]
  reg [31:0] _RAND_0;
  wire [8:0] _T_68; // @[MemPrimitives.scala 325:32:@2496.4]
  wire [8:0] _T_69; // @[MemPrimitives.scala 325:12:@2497.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@2496.4]
  assign _T_69 = io_wPort_0_reset ? 9'h0 : _T_68; // @[MemPrimitives.scala 325:12:@2497.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@2499.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 9'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 9'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@2514.2]
  input        clock, // @[:@2515.4]
  input        reset, // @[:@2516.4]
  input        io_setup_saturate, // @[:@2517.4]
  input        io_input_reset, // @[:@2517.4]
  input        io_input_enable, // @[:@2517.4]
  output [8:0] io_output_count_0, // @[:@2517.4]
  output       io_output_oobs_0, // @[:@2517.4]
  output       io_output_done // @[:@2517.4]
);
  wire  bases_0_clock; // @[Counter.scala 262:53:@2530.4]
  wire  bases_0_reset; // @[Counter.scala 262:53:@2530.4]
  wire [8:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 262:53:@2530.4]
  wire [8:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 262:53:@2530.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 262:53:@2530.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 262:53:@2530.4]
  wire  SRFF_clock; // @[Counter.scala 264:22:@2546.4]
  wire  SRFF_reset; // @[Counter.scala 264:22:@2546.4]
  wire  SRFF_io_input_set; // @[Counter.scala 264:22:@2546.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 264:22:@2546.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 264:22:@2546.4]
  wire  SRFF_io_output; // @[Counter.scala 264:22:@2546.4]
  wire  _T_36; // @[Counter.scala 265:45:@2549.4]
  wire [8:0] _T_48; // @[Counter.scala 288:52:@2574.4]
  wire [9:0] _T_50; // @[Counter.scala 292:33:@2575.4]
  wire [8:0] _T_51; // @[Counter.scala 292:33:@2576.4]
  wire [8:0] _T_52; // @[Counter.scala 292:33:@2577.4]
  wire  _T_57; // @[Counter.scala 294:18:@2579.4]
  wire [8:0] _T_68; // @[Counter.scala 300:115:@2587.4]
  wire [8:0] _T_70; // @[Counter.scala 300:85:@2589.4]
  wire [8:0] _T_71; // @[Counter.scala 300:152:@2590.4]
  wire [8:0] _T_72; // @[Counter.scala 300:74:@2591.4]
  wire  _T_75; // @[Counter.scala 323:102:@2595.4]
  wire  _T_77; // @[Counter.scala 323:130:@2596.4]
  FF_3 bases_0 ( // @[Counter.scala 262:53:@2530.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 264:22:@2546.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 265:45:@2549.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 288:52:@2574.4]
  assign _T_50 = $signed(_T_48) + $signed(9'sh1); // @[Counter.scala 292:33:@2575.4]
  assign _T_51 = $signed(_T_48) + $signed(9'sh1); // @[Counter.scala 292:33:@2576.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 292:33:@2577.4]
  assign _T_57 = $signed(_T_52) >= $signed(9'sh64); // @[Counter.scala 294:18:@2579.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 300:115:@2587.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 9'h0; // @[Counter.scala 300:85:@2589.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 300:152:@2590.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 300:74:@2591.4]
  assign _T_75 = $signed(_T_48) < $signed(9'sh0); // @[Counter.scala 323:102:@2595.4]
  assign _T_77 = $signed(_T_48) >= $signed(9'sh64); // @[Counter.scala 323:130:@2596.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 305:28:@2594.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 323:60:@2598.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 334:20:@2600.4]
  assign bases_0_clock = clock; // @[:@2531.4]
  assign bases_0_reset = reset; // @[:@2532.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 9'h0 : _T_72; // @[Counter.scala 300:31:@2593.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 282:27:@2572.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 285:29:@2573.4]
  assign SRFF_clock = clock; // @[:@2547.4]
  assign SRFF_reset = reset; // @[:@2548.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 265:23:@2551.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 266:25:@2553.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 267:30:@2554.4]
endmodule
module x478_ctrchain( // @[:@2605.2]
  input        clock, // @[:@2606.4]
  input        reset, // @[:@2607.4]
  input        io_input_reset, // @[:@2608.4]
  input        io_input_enable, // @[:@2608.4]
  output [8:0] io_output_counts_0, // @[:@2608.4]
  output       io_output_oobs_0, // @[:@2608.4]
  output       io_output_done // @[:@2608.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 514:46:@2610.4]
  wire  ctrs_0_reset; // @[Counter.scala 514:46:@2610.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 514:46:@2610.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 514:46:@2610.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 514:46:@2610.4]
  wire [8:0] ctrs_0_io_output_count_0; // @[Counter.scala 514:46:@2610.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 514:46:@2610.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 514:46:@2610.4]
  reg  wasDone; // @[Counter.scala 543:24:@2619.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 547:69:@2625.4]
  wire  _T_47; // @[Counter.scala 547:80:@2626.4]
  reg  doneLatch; // @[Counter.scala 551:26:@2631.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 552:48:@2632.4]
  wire  _T_55; // @[Counter.scala 552:19:@2633.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 514:46:@2610.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 547:69:@2625.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 547:80:@2626.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 552:48:@2632.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 552:19:@2633.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 558:32:@2635.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 559:30:@2637.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 547:18:@2628.4]
  assign ctrs_0_clock = clock; // @[:@2611.4]
  assign ctrs_0_reset = reset; // @[:@2612.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 531:29:@2618.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 521:24:@2616.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 525:33:@2617.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@2677.2]
  input   clock, // @[:@2678.4]
  input   reset, // @[:@2679.4]
  input   io_flow, // @[:@2680.4]
  input   io_in, // @[:@2680.4]
  output  io_out // @[:@2680.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2682.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2682.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2682.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2682.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2682.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2682.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@2682.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2695.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2694.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2693.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2692.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2691.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2689.4]
endmodule
module RetimeWrapper_25( // @[:@2805.2]
  input   clock, // @[:@2806.4]
  input   reset, // @[:@2807.4]
  input   io_flow, // @[:@2808.4]
  input   io_in, // @[:@2808.4]
  output  io_out // @[:@2808.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2810.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2810.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2810.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2810.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2810.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2810.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@2810.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2823.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2822.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2821.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2820.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2819.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2817.4]
endmodule
module x499_inr_Foreach_sm( // @[:@2825.2]
  input   clock, // @[:@2826.4]
  input   reset, // @[:@2827.4]
  input   io_enable, // @[:@2828.4]
  output  io_done, // @[:@2828.4]
  output  io_doneLatch, // @[:@2828.4]
  input   io_rst, // @[:@2828.4]
  input   io_ctrDone, // @[:@2828.4]
  output  io_datapathEn, // @[:@2828.4]
  output  io_ctrInc, // @[:@2828.4]
  output  io_ctrRst, // @[:@2828.4]
  input   io_parentAck, // @[:@2828.4]
  input   io_backpressure, // @[:@2828.4]
  input   io_break // @[:@2828.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@2830.4]
  wire  active_reset; // @[Controllers.scala 261:22:@2830.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@2830.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@2830.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@2830.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@2830.4]
  wire  done_clock; // @[Controllers.scala 262:20:@2833.4]
  wire  done_reset; // @[Controllers.scala 262:20:@2833.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@2833.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@2833.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@2833.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@2833.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2867.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2867.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2867.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2867.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2867.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2889.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2889.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2889.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2889.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2889.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2901.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2901.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2901.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2901.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2901.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2909.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2909.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2909.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2909.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2909.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2925.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2925.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2925.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2925.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2925.4]
  wire  _T_80; // @[Controllers.scala 264:48:@2838.4]
  wire  _T_81; // @[Controllers.scala 264:46:@2839.4]
  wire  _T_82; // @[Controllers.scala 264:62:@2840.4]
  wire  _T_83; // @[Controllers.scala 264:60:@2841.4]
  wire  _T_100; // @[package.scala 100:49:@2858.4]
  reg  _T_103; // @[package.scala 48:56:@2859.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@2872.4 package.scala 96:25:@2873.4]
  wire  _T_110; // @[package.scala 100:49:@2874.4]
  reg  _T_113; // @[package.scala 48:56:@2875.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@2877.4]
  wire  _T_118; // @[Controllers.scala 283:41:@2882.4]
  wire  _T_119; // @[Controllers.scala 283:59:@2883.4]
  wire  _T_121; // @[Controllers.scala 284:37:@2886.4]
  wire  _T_124; // @[package.scala 96:25:@2894.4 package.scala 96:25:@2895.4]
  wire  _T_126; // @[package.scala 100:49:@2896.4]
  reg  _T_129; // @[package.scala 48:56:@2897.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@2919.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@2921.4]
  reg  _T_153; // @[package.scala 48:56:@2922.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@2930.4 package.scala 96:25:@2931.4]
  wire  _T_158; // @[Controllers.scala 292:61:@2932.4]
  wire  _T_159; // @[Controllers.scala 292:24:@2933.4]
  SRFF active ( // @[Controllers.scala 261:22:@2830.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@2833.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@2867.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@2889.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2901.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2909.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@2925.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@2838.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@2839.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@2840.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@2841.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@2858.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@2872.4 package.scala 96:25:@2873.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@2874.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@2877.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@2882.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@2883.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@2886.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2894.4 package.scala 96:25:@2895.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@2896.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@2921.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@2930.4 package.scala 96:25:@2931.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@2932.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@2933.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@2900.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@2935.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@2885.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@2888.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@2880.4]
  assign active_clock = clock; // @[:@2831.4]
  assign active_reset = reset; // @[:@2832.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@2843.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@2847.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@2848.4]
  assign done_clock = clock; // @[:@2834.4]
  assign done_reset = reset; // @[:@2835.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@2863.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@2856.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@2857.4]
  assign RetimeWrapper_clock = clock; // @[:@2868.4]
  assign RetimeWrapper_reset = reset; // @[:@2869.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@2871.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@2870.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2890.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2891.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@2893.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@2892.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2902.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2903.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2905.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@2904.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2910.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2911.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2913.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@2912.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2926.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2927.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@2929.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@2928.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x499_inr_Foreach_iiCtr( // @[:@2938.2]
  input   clock, // @[:@2939.4]
  input   reset, // @[:@2940.4]
  input   io_input_enable, // @[:@2941.4]
  input   io_input_reset, // @[:@2941.4]
  output  io_output_issue, // @[:@2941.4]
  output  io_output_done // @[:@2941.4]
);
  reg [4:0] _T_15; // @[Counter.scala 135:22:@2943.4]
  reg [31:0] _RAND_0;
  wire  _T_17; // @[Counter.scala 138:24:@2944.4]
  wire  _T_20; // @[Counter.scala 139:23:@2946.4]
  wire [5:0] _T_26; // @[Counter.scala 141:68:@2949.4]
  wire [4:0] _T_27; // @[Counter.scala 141:68:@2950.4]
  wire [4:0] _T_28; // @[Counter.scala 141:68:@2951.4]
  wire [4:0] _T_29; // @[Counter.scala 141:23:@2952.4]
  wire [4:0] _T_30; // @[Counter.scala 142:19:@2953.4]
  wire [4:0] _T_32; // @[Counter.scala 143:15:@2954.4]
  assign _T_17 = $signed(_T_15) == $signed(5'sh4); // @[Counter.scala 138:24:@2944.4]
  assign _T_20 = $signed(_T_15) == $signed(5'sh0); // @[Counter.scala 139:23:@2946.4]
  assign _T_26 = $signed(_T_15) - $signed(5'sh1); // @[Counter.scala 141:68:@2949.4]
  assign _T_27 = $signed(_T_15) - $signed(5'sh1); // @[Counter.scala 141:68:@2950.4]
  assign _T_28 = $signed(_T_27); // @[Counter.scala 141:68:@2951.4]
  assign _T_29 = _T_20 ? $signed(5'sh4) : $signed(_T_28); // @[Counter.scala 141:23:@2952.4]
  assign _T_30 = io_input_enable ? $signed(_T_29) : $signed(_T_15); // @[Counter.scala 142:19:@2953.4]
  assign _T_32 = io_input_reset ? $signed(5'sh4) : $signed(_T_30); // @[Counter.scala 143:15:@2954.4]
  assign io_output_issue = _T_17 & io_input_enable; // @[Counter.scala 146:21:@2957.4]
  assign io_output_done = _T_20 & io_input_enable; // @[Counter.scala 145:20:@2956.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 5'sh4;
    end else begin
      if (io_input_reset) begin
        _T_15 <= 5'sh4;
      end else begin
        if (io_input_enable) begin
          if (_T_20) begin
            _T_15 <= 5'sh4;
          end else begin
            _T_15 <= _T_28;
          end
        end
      end
    end
  end
endmodule
module SimBlackBoxesfix2fixBox( // @[:@3167.2]
  input  [31:0] io_a, // @[:@3170.4]
  output [31:0] io_b // @[:@3170.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@3183.4]
endmodule
module _( // @[:@3185.2]
  input  [31:0] io_b, // @[:@3188.4]
  output [31:0] io_result // @[:@3188.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3193.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3193.4]
  SimBlackBoxesfix2fixBox SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3193.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 717:17:@3206.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3201.4]
endmodule
module SimBlackBoxesfix2fixBox_1( // @[:@3240.2]
  input  [31:0] io_a, // @[:@3243.4]
  output [32:0] io_b // @[:@3243.4]
);
  wire  _T_20; // @[implicits.scala 70:16:@3253.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 70:16:@3253.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@3258.4]
endmodule
module __1( // @[:@3260.2]
  input  [31:0] io_b, // @[:@3263.4]
  output [32:0] io_result // @[:@3263.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3268.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3268.4]
  SimBlackBoxesfix2fixBox_1 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3268.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 717:17:@3281.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3276.4]
endmodule
module RetimeWrapper_32( // @[:@3338.2]
  input         clock, // @[:@3339.4]
  input         reset, // @[:@3340.4]
  input         io_flow, // @[:@3341.4]
  input  [31:0] io_in, // @[:@3341.4]
  output [31:0] io_out // @[:@3341.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3343.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3343.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3343.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3343.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3343.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3343.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3343.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3356.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3355.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3354.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3353.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3352.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3350.4]
endmodule
module fix2fixBox( // @[:@3358.2]
  input         clock, // @[:@3359.4]
  input         reset, // @[:@3360.4]
  input  [32:0] io_a, // @[:@3361.4]
  input         io_flow, // @[:@3361.4]
  output [31:0] io_b // @[:@3361.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3374.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3374.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3374.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3374.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3374.4]
  RetimeWrapper_32 RetimeWrapper ( // @[package.scala 93:22:@3374.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3381.4]
  assign RetimeWrapper_clock = clock; // @[:@3375.4]
  assign RetimeWrapper_reset = reset; // @[:@3376.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3378.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3377.4]
endmodule
module x739_sum( // @[:@3383.2]
  input         clock, // @[:@3384.4]
  input         reset, // @[:@3385.4]
  input  [31:0] io_a, // @[:@3386.4]
  input  [31:0] io_b, // @[:@3386.4]
  input         io_flow, // @[:@3386.4]
  output [31:0] io_result // @[:@3386.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@3394.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@3394.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@3401.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@3401.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@3419.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@3419.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@3419.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@3419.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@3419.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@3399.4 Math.scala 724:14:@3400.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@3406.4 Math.scala 724:14:@3407.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@3408.4]
  __1 _ ( // @[Math.scala 720:24:@3394.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __1 __1 ( // @[Math.scala 720:24:@3401.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 141:30:@3419.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@3399.4 Math.scala 724:14:@3400.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@3406.4 Math.scala 724:14:@3407.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@3408.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@3427.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@3397.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@3404.4]
  assign fix2fixBox_clock = clock; // @[:@3420.4]
  assign fix2fixBox_reset = reset; // @[:@3421.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@3422.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@3425.4]
endmodule
module x485_sub( // @[:@3572.2]
  input         clock, // @[:@3573.4]
  input         reset, // @[:@3574.4]
  input  [31:0] io_a, // @[:@3575.4]
  input  [31:0] io_b, // @[:@3575.4]
  input         io_flow, // @[:@3575.4]
  output [31:0] io_result // @[:@3575.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@3583.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@3583.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@3590.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@3590.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@3609.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@3609.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@3609.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@3609.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@3609.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@3588.4 Math.scala 724:14:@3589.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@3595.4 Math.scala 724:14:@3596.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@3597.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@3598.4]
  __1 _ ( // @[Math.scala 720:24:@3583.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __1 __1 ( // @[Math.scala 720:24:@3590.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 182:30:@3609.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@3588.4 Math.scala 724:14:@3589.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@3595.4 Math.scala 724:14:@3596.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@3597.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@3598.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@3617.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@3586.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@3593.4]
  assign fix2fixBox_clock = clock; // @[:@3610.4]
  assign fix2fixBox_reset = reset; // @[:@3611.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@3612.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@3615.4]
endmodule
module RetimeWrapper_36( // @[:@4009.2]
  input         clock, // @[:@4010.4]
  input         reset, // @[:@4011.4]
  input         io_flow, // @[:@4012.4]
  input  [35:0] io_in, // @[:@4012.4]
  output [35:0] io_out // @[:@4012.4]
);
  wire [35:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@4014.4]
  wire [35:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@4014.4]
  wire [35:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@4014.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@4014.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@4014.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@4014.4]
  RetimeShiftRegister #(.WIDTH(36), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@4014.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@4027.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@4026.4]
  assign sr_init = 36'h0; // @[RetimeShiftRegister.scala 19:16:@4025.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@4024.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@4023.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@4021.4]
endmodule
module RetimeWrapper_37( // @[:@4041.2]
  input         clock, // @[:@4042.4]
  input         reset, // @[:@4043.4]
  input         io_flow, // @[:@4044.4]
  input  [37:0] io_in, // @[:@4044.4]
  output [37:0] io_out // @[:@4044.4]
);
  wire [37:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@4046.4]
  wire [37:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@4046.4]
  wire [37:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@4046.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@4046.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@4046.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@4046.4]
  RetimeShiftRegister #(.WIDTH(38), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@4046.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@4059.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@4058.4]
  assign sr_init = 38'h0; // @[RetimeShiftRegister.scala 19:16:@4057.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@4056.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@4055.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@4053.4]
endmodule
module SimBlackBoxesfix2fixBox_9( // @[:@4061.2]
  input  [31:0] io_a, // @[:@4064.4]
  output [63:0] io_b // @[:@4064.4]
);
  wire  _T_20; // @[implicits.scala 70:16:@4074.4]
  wire [31:0] _T_24; // @[Bitwise.scala 72:12:@4077.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 70:16:@4074.4]
  assign _T_24 = _T_20 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@4077.4]
  assign io_b = {_T_24,io_a}; // @[SimBlackBoxes.scala 99:40:@4081.4]
endmodule
module x491( // @[:@4083.2]
  input  [31:0] io_b, // @[:@4086.4]
  output [63:0] io_result // @[:@4086.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@4091.4]
  wire [63:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@4091.4]
  SimBlackBoxesfix2fixBox_9 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@4091.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 717:17:@4104.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@4099.4]
endmodule
module RetimeWrapper_38( // @[:@4118.2]
  input         clock, // @[:@4119.4]
  input         reset, // @[:@4120.4]
  input         io_flow, // @[:@4121.4]
  input  [63:0] io_in, // @[:@4121.4]
  output [63:0] io_out // @[:@4121.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@4123.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@4123.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@4123.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@4123.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@4123.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@4123.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@4123.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@4136.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@4135.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@4134.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@4133.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@4132.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@4130.4]
endmodule
module SimBlackBoxesfix2fixBox_10( // @[:@4138.2]
  input  [63:0] io_a, // @[:@4141.4]
  output [64:0] io_b // @[:@4141.4]
);
  wire  _T_20; // @[implicits.scala 70:16:@4151.4]
  assign _T_20 = io_a[63]; // @[implicits.scala 70:16:@4151.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@4156.4]
endmodule
module __9( // @[:@4158.2]
  input  [63:0] io_b, // @[:@4161.4]
  output [64:0] io_result // @[:@4161.4]
);
  wire [63:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@4166.4]
  wire [64:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@4166.4]
  SimBlackBoxesfix2fixBox_10 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@4166.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 717:17:@4179.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@4174.4]
endmodule
module RetimeWrapper_39( // @[:@4236.2]
  input         clock, // @[:@4237.4]
  input         reset, // @[:@4238.4]
  input         io_flow, // @[:@4239.4]
  input  [63:0] io_in, // @[:@4239.4]
  output [63:0] io_out // @[:@4239.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@4241.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@4241.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@4241.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@4241.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@4241.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@4241.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@4241.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@4254.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@4253.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@4252.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@4251.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@4250.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@4248.4]
endmodule
module fix2fixBox_4( // @[:@4256.2]
  input         clock, // @[:@4257.4]
  input         reset, // @[:@4258.4]
  input  [64:0] io_a, // @[:@4259.4]
  input         io_flow, // @[:@4259.4]
  output [63:0] io_b // @[:@4259.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4272.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4272.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4272.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@4272.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@4272.4]
  RetimeWrapper_39 RetimeWrapper ( // @[package.scala 93:22:@4272.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@4279.4]
  assign RetimeWrapper_clock = clock; // @[:@4273.4]
  assign RetimeWrapper_reset = reset; // @[:@4274.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@4276.4]
  assign RetimeWrapper_io_in = io_a[63:0]; // @[package.scala 94:16:@4275.4]
endmodule
module x493_sum( // @[:@4281.2]
  input         clock, // @[:@4282.4]
  input         reset, // @[:@4283.4]
  input  [63:0] io_a, // @[:@4284.4]
  input  [63:0] io_b, // @[:@4284.4]
  input         io_flow, // @[:@4284.4]
  output [63:0] io_result // @[:@4284.4]
);
  wire [63:0] __io_b; // @[Math.scala 720:24:@4292.4]
  wire [64:0] __io_result; // @[Math.scala 720:24:@4292.4]
  wire [63:0] __1_io_b; // @[Math.scala 720:24:@4299.4]
  wire [64:0] __1_io_result; // @[Math.scala 720:24:@4299.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4317.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4317.4]
  wire [64:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4317.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4317.4]
  wire [63:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4317.4]
  wire [64:0] a_upcast_number; // @[Math.scala 723:22:@4297.4 Math.scala 724:14:@4298.4]
  wire [64:0] b_upcast_number; // @[Math.scala 723:22:@4304.4 Math.scala 724:14:@4305.4]
  wire [65:0] _T_21; // @[Math.scala 136:37:@4306.4]
  __9 _ ( // @[Math.scala 720:24:@4292.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __9 __1 ( // @[Math.scala 720:24:@4299.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@4317.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@4297.4 Math.scala 724:14:@4298.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@4304.4 Math.scala 724:14:@4305.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4306.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4325.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@4295.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@4302.4]
  assign fix2fixBox_clock = clock; // @[:@4318.4]
  assign fix2fixBox_reset = reset; // @[:@4319.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4320.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4323.4]
endmodule
module RetimeWrapper_45( // @[:@4499.2]
  input         clock, // @[:@4500.4]
  input         reset, // @[:@4501.4]
  input         io_flow, // @[:@4502.4]
  input  [31:0] io_in, // @[:@4502.4]
  output [31:0] io_out // @[:@4502.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@4504.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@4504.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@4504.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@4504.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@4504.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@4504.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@4504.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@4517.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@4516.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@4515.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@4514.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@4513.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@4511.4]
endmodule
module x499_inr_Foreach_kernelx499_inr_Foreach_concrete1( // @[:@4551.2]
  input         clock, // @[:@4552.4]
  input         reset, // @[:@4553.4]
  input  [63:0] io_in_x468_A_dram_number, // @[:@4554.4]
  output [95:0] io_in_x475_fifo_wPort_0_data_0, // @[:@4554.4]
  output        io_in_x475_fifo_wPort_0_en_0, // @[:@4554.4]
  input         io_in_x475_fifo_full, // @[:@4554.4]
  output        io_in_x475_fifo_active_0_in, // @[:@4554.4]
  input         io_in_x475_fifo_active_0_out, // @[:@4554.4]
  input         io_in_x474_ready, // @[:@4554.4]
  output        io_in_x474_valid, // @[:@4554.4]
  output [63:0] io_in_x474_bits_addr, // @[:@4554.4]
  output [31:0] io_in_x474_bits_size, // @[:@4554.4]
  output [63:0] io_in_instrctrs_2_cycs, // @[:@4554.4]
  output [63:0] io_in_instrctrs_2_iters, // @[:@4554.4]
  output [63:0] io_in_instrctrs_2_stalls, // @[:@4554.4]
  output [63:0] io_in_instrctrs_2_idles, // @[:@4554.4]
  input         io_sigsIn_done, // @[:@4554.4]
  input         io_sigsIn_iiIssue, // @[:@4554.4]
  input         io_sigsIn_backpressure, // @[:@4554.4]
  input         io_sigsIn_datapathEn, // @[:@4554.4]
  input         io_sigsIn_baseEn, // @[:@4554.4]
  input         io_sigsIn_break, // @[:@4554.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@4554.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@4554.4]
  input         io_rr // @[:@4554.4]
);
  wire  cycles_x499_inr_Foreach_clock; // @[sm_x499_inr_Foreach.scala 68:43:@4682.4]
  wire  cycles_x499_inr_Foreach_reset; // @[sm_x499_inr_Foreach.scala 68:43:@4682.4]
  wire  cycles_x499_inr_Foreach_io_enable; // @[sm_x499_inr_Foreach.scala 68:43:@4682.4]
  wire [63:0] cycles_x499_inr_Foreach_io_count; // @[sm_x499_inr_Foreach.scala 68:43:@4682.4]
  wire  iters_x499_inr_Foreach_clock; // @[sm_x499_inr_Foreach.scala 69:42:@4685.4]
  wire  iters_x499_inr_Foreach_reset; // @[sm_x499_inr_Foreach.scala 69:42:@4685.4]
  wire  iters_x499_inr_Foreach_io_enable; // @[sm_x499_inr_Foreach.scala 69:42:@4685.4]
  wire [63:0] iters_x499_inr_Foreach_io_count; // @[sm_x499_inr_Foreach.scala 69:42:@4685.4]
  wire  stalls_x499_inr_Foreach_clock; // @[sm_x499_inr_Foreach.scala 72:43:@4694.4]
  wire  stalls_x499_inr_Foreach_reset; // @[sm_x499_inr_Foreach.scala 72:43:@4694.4]
  wire  stalls_x499_inr_Foreach_io_enable; // @[sm_x499_inr_Foreach.scala 72:43:@4694.4]
  wire [63:0] stalls_x499_inr_Foreach_io_count; // @[sm_x499_inr_Foreach.scala 72:43:@4694.4]
  wire  idles_x499_inr_Foreach_clock; // @[sm_x499_inr_Foreach.scala 73:42:@4697.4]
  wire  idles_x499_inr_Foreach_reset; // @[sm_x499_inr_Foreach.scala 73:42:@4697.4]
  wire  idles_x499_inr_Foreach_io_enable; // @[sm_x499_inr_Foreach.scala 73:42:@4697.4]
  wire [63:0] idles_x499_inr_Foreach_io_count; // @[sm_x499_inr_Foreach.scala 73:42:@4697.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4700.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4700.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4700.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@4700.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@4700.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@4727.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@4727.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4738.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4738.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@4738.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@4738.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@4738.4]
  wire  x739_sum_1_clock; // @[Math.scala 150:24:@4756.4]
  wire  x739_sum_1_reset; // @[Math.scala 150:24:@4756.4]
  wire [31:0] x739_sum_1_io_a; // @[Math.scala 150:24:@4756.4]
  wire [31:0] x739_sum_1_io_b; // @[Math.scala 150:24:@4756.4]
  wire  x739_sum_1_io_flow; // @[Math.scala 150:24:@4756.4]
  wire [31:0] x739_sum_1_io_result; // @[Math.scala 150:24:@4756.4]
  wire  x485_sub_1_clock; // @[Math.scala 191:24:@4793.4]
  wire  x485_sub_1_reset; // @[Math.scala 191:24:@4793.4]
  wire [31:0] x485_sub_1_io_a; // @[Math.scala 191:24:@4793.4]
  wire [31:0] x485_sub_1_io_b; // @[Math.scala 191:24:@4793.4]
  wire  x485_sub_1_io_flow; // @[Math.scala 191:24:@4793.4]
  wire [31:0] x485_sub_1_io_result; // @[Math.scala 191:24:@4793.4]
  wire  x486_sum_1_clock; // @[Math.scala 150:24:@4805.4]
  wire  x486_sum_1_reset; // @[Math.scala 150:24:@4805.4]
  wire [31:0] x486_sum_1_io_a; // @[Math.scala 150:24:@4805.4]
  wire [31:0] x486_sum_1_io_b; // @[Math.scala 150:24:@4805.4]
  wire  x486_sum_1_io_flow; // @[Math.scala 150:24:@4805.4]
  wire [31:0] x486_sum_1_io_result; // @[Math.scala 150:24:@4805.4]
  wire  x487_sum_1_clock; // @[Math.scala 150:24:@4817.4]
  wire  x487_sum_1_reset; // @[Math.scala 150:24:@4817.4]
  wire [31:0] x487_sum_1_io_a; // @[Math.scala 150:24:@4817.4]
  wire [31:0] x487_sum_1_io_b; // @[Math.scala 150:24:@4817.4]
  wire  x487_sum_1_io_flow; // @[Math.scala 150:24:@4817.4]
  wire [31:0] x487_sum_1_io_result; // @[Math.scala 150:24:@4817.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@4846.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@4846.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@4846.4]
  wire [35:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@4846.4]
  wire [35:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@4846.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@4858.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@4858.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@4858.4]
  wire [37:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@4858.4]
  wire [37:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@4858.4]
  wire [31:0] x491_1_io_b; // @[Math.scala 720:24:@4868.4]
  wire [63:0] x491_1_io_result; // @[Math.scala 720:24:@4868.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@4878.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@4878.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@4878.4]
  wire [63:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@4878.4]
  wire [63:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@4878.4]
  wire  x493_sum_1_clock; // @[Math.scala 150:24:@4887.4]
  wire  x493_sum_1_reset; // @[Math.scala 150:24:@4887.4]
  wire [63:0] x493_sum_1_io_a; // @[Math.scala 150:24:@4887.4]
  wire [63:0] x493_sum_1_io_b; // @[Math.scala 150:24:@4887.4]
  wire  x493_sum_1_io_flow; // @[Math.scala 150:24:@4887.4]
  wire [63:0] x493_sum_1_io_result; // @[Math.scala 150:24:@4887.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@4898.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@4898.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@4898.4]
  wire [63:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@4898.4]
  wire [63:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@4898.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@4912.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@4912.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@4912.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@4912.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@4912.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@4922.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@4922.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@4922.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@4922.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@4922.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@4932.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@4932.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@4932.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@4932.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@4932.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@4950.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@4950.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@4950.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@4950.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@4950.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@4960.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@4960.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@4960.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@4960.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@4960.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@4976.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@4976.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@4976.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@4976.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@4976.4]
  wire  _T_318; // @[package.scala 100:49:@4689.4]
  reg  _T_321; // @[package.scala 48:56:@4690.4]
  reg [31:0] _RAND_0;
  wire  _T_326; // @[package.scala 96:25:@4705.4 package.scala 96:25:@4706.4]
  wire  _T_329; // @[sm_x499_inr_Foreach.scala 74:66:@4708.4]
  wire  _T_330; // @[sm_x499_inr_Foreach.scala 74:93:@4709.4]
  wire  _T_331; // @[sm_x499_inr_Foreach.scala 74:91:@4710.4]
  wire  _T_332; // @[sm_x499_inr_Foreach.scala 74:121:@4711.4]
  wire  _T_333; // @[sm_x499_inr_Foreach.scala 74:63:@4712.4]
  wire  _T_352; // @[package.scala 96:25:@4743.4 package.scala 96:25:@4744.4]
  wire  _T_355; // @[sm_x499_inr_Foreach.scala 81:18:@4746.4]
  wire  _T_357; // @[sm_x499_inr_Foreach.scala 81:43:@4748.4]
  wire [31:0] b479_number; // @[Math.scala 723:22:@4732.4 Math.scala 724:14:@4733.4]
  wire [32:0] _GEN_0; // @[Math.scala 461:32:@4752.4]
  wire [32:0] _T_360; // @[Math.scala 461:32:@4752.4]
  wire [31:0] x739_sum_number; // @[Math.scala 154:22:@4762.4 Math.scala 155:14:@4763.4]
  wire  _T_366; // @[FixedPoint.scala 50:25:@4767.4]
  wire [3:0] _T_370; // @[Bitwise.scala 72:12:@4769.4]
  wire [27:0] _T_371; // @[FixedPoint.scala 18:52:@4770.4]
  wire  _T_377; // @[Math.scala 451:55:@4772.4]
  wire [3:0] _T_378; // @[FixedPoint.scala 18:52:@4773.4]
  wire  _T_384; // @[Math.scala 451:110:@4775.4]
  wire  _T_385; // @[Math.scala 451:94:@4776.4]
  wire [31:0] _T_387; // @[Cat.scala 30:58:@4778.4]
  wire [31:0] x482_1_number; // @[Math.scala 454:20:@4779.4]
  wire [35:0] _GEN_1; // @[Math.scala 461:32:@4784.4]
  wire [35:0] _T_392; // @[Math.scala 461:32:@4784.4]
  wire [37:0] _GEN_2; // @[Math.scala 461:32:@4789.4]
  wire [37:0] _T_395; // @[Math.scala 461:32:@4789.4]
  wire [31:0] x487_sum_number; // @[Math.scala 154:22:@4823.4 Math.scala 155:14:@4824.4]
  wire  _T_415; // @[FixedPoint.scala 50:25:@4828.4]
  wire [3:0] _T_419; // @[Bitwise.scala 72:12:@4830.4]
  wire [27:0] _T_420; // @[FixedPoint.scala 18:52:@4831.4]
  wire  _T_426; // @[Math.scala 451:55:@4833.4]
  wire [3:0] _T_427; // @[FixedPoint.scala 18:52:@4834.4]
  wire  _T_433; // @[Math.scala 451:110:@4836.4]
  wire  _T_434; // @[Math.scala 451:94:@4837.4]
  wire [31:0] _T_436; // @[Cat.scala 30:58:@4839.4]
  wire [31:0] x488_1_number; // @[Math.scala 454:20:@4840.4]
  wire [35:0] _GEN_3; // @[Math.scala 461:32:@4845.4]
  wire [37:0] _GEN_4; // @[Math.scala 461:32:@4857.4]
  wire [37:0] _T_448; // @[package.scala 96:25:@4863.4 package.scala 96:25:@4864.4]
  wire [31:0] x741_1_number; // @[Math.scala 459:22:@4856.4 Math.scala 461:14:@4865.4]
  wire [63:0] x759_x493_sum_D1_number; // @[package.scala 96:25:@4903.4 package.scala 96:25:@4904.4]
  wire [96:0] x494_tuple; // @[Cat.scala 30:58:@4908.4]
  wire  _T_483; // @[package.scala 96:25:@4937.4 package.scala 96:25:@4938.4]
  wire  _T_485; // @[implicits.scala 56:10:@4939.4]
  wire  x760_x495_D4; // @[package.scala 96:25:@4917.4 package.scala 96:25:@4918.4]
  wire  _T_486; // @[sm_x499_inr_Foreach.scala 119:121:@4940.4]
  wire  x761_b480_D4; // @[package.scala 96:25:@4927.4 package.scala 96:25:@4928.4]
  wire  _T_487; // @[sm_x499_inr_Foreach.scala 119:127:@4941.4]
  wire [31:0] x762_x486_sum_D1_number; // @[package.scala 96:25:@4955.4 package.scala 96:25:@4956.4]
  wire [31:0] x763_x485_sub_D2_number; // @[package.scala 96:25:@4965.4 package.scala 96:25:@4966.4]
  wire [63:0] _T_502; // @[Cat.scala 30:58:@4969.4]
  wire [35:0] _T_443; // @[package.scala 96:25:@4851.4 package.scala 96:25:@4852.4]
  wire [31:0] x489_1_number; // @[Math.scala 459:22:@4844.4 Math.scala 461:14:@4853.4]
  wire  _T_504; // @[sm_x499_inr_Foreach.scala 132:121:@4972.4]
  wire  _T_510; // @[package.scala 96:25:@4981.4 package.scala 96:25:@4982.4]
  wire  _T_512; // @[implicits.scala 56:10:@4983.4]
  wire  _T_513; // @[sm_x499_inr_Foreach.scala 132:138:@4984.4]
  wire  _T_515; // @[sm_x499_inr_Foreach.scala 132:235:@4986.4]
  wire  _T_516; // @[sm_x499_inr_Foreach.scala 132:254:@4987.4]
  InstrumentationCounter cycles_x499_inr_Foreach ( // @[sm_x499_inr_Foreach.scala 68:43:@4682.4]
    .clock(cycles_x499_inr_Foreach_clock),
    .reset(cycles_x499_inr_Foreach_reset),
    .io_enable(cycles_x499_inr_Foreach_io_enable),
    .io_count(cycles_x499_inr_Foreach_io_count)
  );
  InstrumentationCounter iters_x499_inr_Foreach ( // @[sm_x499_inr_Foreach.scala 69:42:@4685.4]
    .clock(iters_x499_inr_Foreach_clock),
    .reset(iters_x499_inr_Foreach_reset),
    .io_enable(iters_x499_inr_Foreach_io_enable),
    .io_count(iters_x499_inr_Foreach_io_count)
  );
  InstrumentationCounter stalls_x499_inr_Foreach ( // @[sm_x499_inr_Foreach.scala 72:43:@4694.4]
    .clock(stalls_x499_inr_Foreach_clock),
    .reset(stalls_x499_inr_Foreach_reset),
    .io_enable(stalls_x499_inr_Foreach_io_enable),
    .io_count(stalls_x499_inr_Foreach_io_count)
  );
  InstrumentationCounter idles_x499_inr_Foreach ( // @[sm_x499_inr_Foreach.scala 73:42:@4697.4]
    .clock(idles_x499_inr_Foreach_clock),
    .reset(idles_x499_inr_Foreach_reset),
    .io_enable(idles_x499_inr_Foreach_io_enable),
    .io_count(idles_x499_inr_Foreach_io_count)
  );
  RetimeWrapper_25 RetimeWrapper ( // @[package.scala 93:22:@4700.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  _ _ ( // @[Math.scala 720:24:@4727.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@4738.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x739_sum x739_sum_1 ( // @[Math.scala 150:24:@4756.4]
    .clock(x739_sum_1_clock),
    .reset(x739_sum_1_reset),
    .io_a(x739_sum_1_io_a),
    .io_b(x739_sum_1_io_b),
    .io_flow(x739_sum_1_io_flow),
    .io_result(x739_sum_1_io_result)
  );
  x485_sub x485_sub_1 ( // @[Math.scala 191:24:@4793.4]
    .clock(x485_sub_1_clock),
    .reset(x485_sub_1_reset),
    .io_a(x485_sub_1_io_a),
    .io_b(x485_sub_1_io_b),
    .io_flow(x485_sub_1_io_flow),
    .io_result(x485_sub_1_io_result)
  );
  x739_sum x486_sum_1 ( // @[Math.scala 150:24:@4805.4]
    .clock(x486_sum_1_clock),
    .reset(x486_sum_1_reset),
    .io_a(x486_sum_1_io_a),
    .io_b(x486_sum_1_io_b),
    .io_flow(x486_sum_1_io_flow),
    .io_result(x486_sum_1_io_result)
  );
  x739_sum x487_sum_1 ( // @[Math.scala 150:24:@4817.4]
    .clock(x487_sum_1_clock),
    .reset(x487_sum_1_reset),
    .io_a(x487_sum_1_io_a),
    .io_b(x487_sum_1_io_b),
    .io_flow(x487_sum_1_io_flow),
    .io_result(x487_sum_1_io_result)
  );
  RetimeWrapper_36 RetimeWrapper_2 ( // @[package.scala 93:22:@4846.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_3 ( // @[package.scala 93:22:@4858.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x491 x491_1 ( // @[Math.scala 720:24:@4868.4]
    .io_b(x491_1_io_b),
    .io_result(x491_1_io_result)
  );
  RetimeWrapper_38 RetimeWrapper_4 ( // @[package.scala 93:22:@4878.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x493_sum x493_sum_1 ( // @[Math.scala 150:24:@4887.4]
    .clock(x493_sum_1_clock),
    .reset(x493_sum_1_reset),
    .io_a(x493_sum_1_io_a),
    .io_b(x493_sum_1_io_b),
    .io_flow(x493_sum_1_io_flow),
    .io_result(x493_sum_1_io_result)
  );
  RetimeWrapper_38 RetimeWrapper_5 ( // @[package.scala 93:22:@4898.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_6 ( // @[package.scala 93:22:@4912.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_7 ( // @[package.scala 93:22:@4922.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_8 ( // @[package.scala 93:22:@4932.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_9 ( // @[package.scala 93:22:@4950.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_45 RetimeWrapper_10 ( // @[package.scala 93:22:@4960.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_11 ( // @[package.scala 93:22:@4976.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  assign _T_318 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@4689.4]
  assign _T_326 = RetimeWrapper_io_out; // @[package.scala 96:25:@4705.4 package.scala 96:25:@4706.4]
  assign _T_329 = ~ _T_326; // @[sm_x499_inr_Foreach.scala 74:66:@4708.4]
  assign _T_330 = ~ io_in_x475_fifo_active_0_out; // @[sm_x499_inr_Foreach.scala 74:93:@4709.4]
  assign _T_331 = _T_329 | _T_330; // @[sm_x499_inr_Foreach.scala 74:91:@4710.4]
  assign _T_332 = _T_331 & io_in_x474_ready; // @[sm_x499_inr_Foreach.scala 74:121:@4711.4]
  assign _T_333 = ~ _T_332; // @[sm_x499_inr_Foreach.scala 74:63:@4712.4]
  assign _T_352 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@4743.4 package.scala 96:25:@4744.4]
  assign _T_355 = ~ _T_352; // @[sm_x499_inr_Foreach.scala 81:18:@4746.4]
  assign _T_357 = _T_355 | _T_330; // @[sm_x499_inr_Foreach.scala 81:43:@4748.4]
  assign b479_number = __io_result; // @[Math.scala 723:22:@4732.4 Math.scala 724:14:@4733.4]
  assign _GEN_0 = {{1'd0}, b479_number}; // @[Math.scala 461:32:@4752.4]
  assign _T_360 = _GEN_0 << 1; // @[Math.scala 461:32:@4752.4]
  assign x739_sum_number = x739_sum_1_io_result; // @[Math.scala 154:22:@4762.4 Math.scala 155:14:@4763.4]
  assign _T_366 = x739_sum_number[31]; // @[FixedPoint.scala 50:25:@4767.4]
  assign _T_370 = _T_366 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@4769.4]
  assign _T_371 = x739_sum_number[31:4]; // @[FixedPoint.scala 18:52:@4770.4]
  assign _T_377 = _T_371 == 28'hfffffff; // @[Math.scala 451:55:@4772.4]
  assign _T_378 = x739_sum_number[3:0]; // @[FixedPoint.scala 18:52:@4773.4]
  assign _T_384 = _T_378 != 4'h0; // @[Math.scala 451:110:@4775.4]
  assign _T_385 = _T_377 & _T_384; // @[Math.scala 451:94:@4776.4]
  assign _T_387 = {_T_370,_T_371}; // @[Cat.scala 30:58:@4778.4]
  assign x482_1_number = _T_385 ? 32'h0 : _T_387; // @[Math.scala 454:20:@4779.4]
  assign _GEN_1 = {{4'd0}, x482_1_number}; // @[Math.scala 461:32:@4784.4]
  assign _T_392 = _GEN_1 << 4; // @[Math.scala 461:32:@4784.4]
  assign _GEN_2 = {{6'd0}, x482_1_number}; // @[Math.scala 461:32:@4789.4]
  assign _T_395 = _GEN_2 << 6; // @[Math.scala 461:32:@4789.4]
  assign x487_sum_number = x487_sum_1_io_result; // @[Math.scala 154:22:@4823.4 Math.scala 155:14:@4824.4]
  assign _T_415 = x487_sum_number[31]; // @[FixedPoint.scala 50:25:@4828.4]
  assign _T_419 = _T_415 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@4830.4]
  assign _T_420 = x487_sum_number[31:4]; // @[FixedPoint.scala 18:52:@4831.4]
  assign _T_426 = _T_420 == 28'hfffffff; // @[Math.scala 451:55:@4833.4]
  assign _T_427 = x487_sum_number[3:0]; // @[FixedPoint.scala 18:52:@4834.4]
  assign _T_433 = _T_427 != 4'h0; // @[Math.scala 451:110:@4836.4]
  assign _T_434 = _T_426 & _T_433; // @[Math.scala 451:94:@4837.4]
  assign _T_436 = {_T_419,_T_420}; // @[Cat.scala 30:58:@4839.4]
  assign x488_1_number = _T_434 ? 32'h0 : _T_436; // @[Math.scala 454:20:@4840.4]
  assign _GEN_3 = {{4'd0}, x488_1_number}; // @[Math.scala 461:32:@4845.4]
  assign _GEN_4 = {{6'd0}, x488_1_number}; // @[Math.scala 461:32:@4857.4]
  assign _T_448 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@4863.4 package.scala 96:25:@4864.4]
  assign x741_1_number = _T_448[31:0]; // @[Math.scala 459:22:@4856.4 Math.scala 461:14:@4865.4]
  assign x759_x493_sum_D1_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@4903.4 package.scala 96:25:@4904.4]
  assign x494_tuple = {1'h1,x741_1_number,x759_x493_sum_D1_number}; // @[Cat.scala 30:58:@4908.4]
  assign _T_483 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@4937.4 package.scala 96:25:@4938.4]
  assign _T_485 = io_rr ? _T_483 : 1'h0; // @[implicits.scala 56:10:@4939.4]
  assign x760_x495_D4 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@4917.4 package.scala 96:25:@4918.4]
  assign _T_486 = _T_485 & x760_x495_D4; // @[sm_x499_inr_Foreach.scala 119:121:@4940.4]
  assign x761_b480_D4 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@4927.4 package.scala 96:25:@4928.4]
  assign _T_487 = _T_486 & x761_b480_D4; // @[sm_x499_inr_Foreach.scala 119:127:@4941.4]
  assign x762_x486_sum_D1_number = RetimeWrapper_9_io_out; // @[package.scala 96:25:@4955.4 package.scala 96:25:@4956.4]
  assign x763_x485_sub_D2_number = RetimeWrapper_10_io_out; // @[package.scala 96:25:@4965.4 package.scala 96:25:@4966.4]
  assign _T_502 = {x762_x486_sum_D1_number,x763_x485_sub_D2_number}; // @[Cat.scala 30:58:@4969.4]
  assign _T_443 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@4851.4 package.scala 96:25:@4852.4]
  assign x489_1_number = _T_443[31:0]; // @[Math.scala 459:22:@4844.4 Math.scala 461:14:@4853.4]
  assign _T_504 = ~ io_sigsIn_break; // @[sm_x499_inr_Foreach.scala 132:121:@4972.4]
  assign _T_510 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@4981.4 package.scala 96:25:@4982.4]
  assign _T_512 = io_rr ? _T_510 : 1'h0; // @[implicits.scala 56:10:@4983.4]
  assign _T_513 = _T_504 & _T_512; // @[sm_x499_inr_Foreach.scala 132:138:@4984.4]
  assign _T_515 = _T_513 & _T_504; // @[sm_x499_inr_Foreach.scala 132:235:@4986.4]
  assign _T_516 = _T_515 & io_sigsIn_backpressure; // @[sm_x499_inr_Foreach.scala 132:254:@4987.4]
  assign io_in_x475_fifo_wPort_0_data_0 = {_T_502,x489_1_number}; // @[MemInterfaceType.scala 90:56:@4990.4]
  assign io_in_x475_fifo_wPort_0_en_0 = _T_516 & x761_b480_D4; // @[MemInterfaceType.scala 93:57:@4992.4]
  assign io_in_x475_fifo_active_0_in = RetimeWrapper_7_io_out; // @[MemInterfaceType.scala 147:18:@4994.4]
  assign io_in_x474_valid = _T_487 & io_sigsIn_backpressure; // @[sm_x499_inr_Foreach.scala 119:18:@4943.4]
  assign io_in_x474_bits_addr = x494_tuple[63:0]; // @[sm_x499_inr_Foreach.scala 120:22:@4945.4]
  assign io_in_x474_bits_size = x494_tuple[95:64]; // @[sm_x499_inr_Foreach.scala 121:22:@4947.4]
  assign io_in_instrctrs_2_cycs = cycles_x499_inr_Foreach_io_count; // @[Ledger.scala 293:21:@4719.4]
  assign io_in_instrctrs_2_iters = iters_x499_inr_Foreach_io_count; // @[Ledger.scala 294:22:@4720.4]
  assign io_in_instrctrs_2_stalls = stalls_x499_inr_Foreach_io_count; // @[Ledger.scala 295:23:@4721.4]
  assign io_in_instrctrs_2_idles = idles_x499_inr_Foreach_io_count; // @[Ledger.scala 296:22:@4722.4]
  assign cycles_x499_inr_Foreach_clock = clock; // @[:@4683.4]
  assign cycles_x499_inr_Foreach_reset = reset; // @[:@4684.4]
  assign cycles_x499_inr_Foreach_io_enable = io_sigsIn_baseEn; // @[sm_x499_inr_Foreach.scala 70:41:@4688.4]
  assign iters_x499_inr_Foreach_clock = clock; // @[:@4686.4]
  assign iters_x499_inr_Foreach_reset = reset; // @[:@4687.4]
  assign iters_x499_inr_Foreach_io_enable = io_sigsIn_done & _T_321; // @[sm_x499_inr_Foreach.scala 71:40:@4693.4]
  assign stalls_x499_inr_Foreach_clock = clock; // @[:@4695.4]
  assign stalls_x499_inr_Foreach_reset = reset; // @[:@4696.4]
  assign stalls_x499_inr_Foreach_io_enable = io_sigsIn_baseEn & _T_333; // @[sm_x499_inr_Foreach.scala 74:41:@4714.4]
  assign idles_x499_inr_Foreach_clock = clock; // @[:@4698.4]
  assign idles_x499_inr_Foreach_reset = reset; // @[:@4699.4]
  assign idles_x499_inr_Foreach_io_enable = 1'h0; // @[sm_x499_inr_Foreach.scala 75:40:@4718.4]
  assign RetimeWrapper_clock = clock; // @[:@4701.4]
  assign RetimeWrapper_reset = reset; // @[:@4702.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@4704.4]
  assign RetimeWrapper_io_in = io_in_x475_fifo_full; // @[package.scala 94:16:@4703.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@4730.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4739.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4740.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@4742.4]
  assign RetimeWrapper_1_io_in = io_in_x475_fifo_full; // @[package.scala 94:16:@4741.4]
  assign x739_sum_1_clock = clock; // @[:@4757.4]
  assign x739_sum_1_reset = reset; // @[:@4758.4]
  assign x739_sum_1_io_a = _T_360[31:0]; // @[Math.scala 151:17:@4759.4]
  assign x739_sum_1_io_b = __io_result; // @[Math.scala 152:17:@4760.4]
  assign x739_sum_1_io_flow = _T_357 & io_in_x474_ready; // @[Math.scala 153:20:@4761.4]
  assign x485_sub_1_clock = clock; // @[:@4794.4]
  assign x485_sub_1_reset = reset; // @[:@4795.4]
  assign x485_sub_1_io_a = x739_sum_1_io_result; // @[Math.scala 192:17:@4796.4]
  assign x485_sub_1_io_b = _T_392[31:0]; // @[Math.scala 193:17:@4797.4]
  assign x485_sub_1_io_flow = _T_357 & io_in_x474_ready; // @[Math.scala 194:20:@4798.4]
  assign x486_sum_1_clock = clock; // @[:@4806.4]
  assign x486_sum_1_reset = reset; // @[:@4807.4]
  assign x486_sum_1_io_a = x485_sub_1_io_result; // @[Math.scala 151:17:@4808.4]
  assign x486_sum_1_io_b = 32'h3; // @[Math.scala 152:17:@4809.4]
  assign x486_sum_1_io_flow = _T_357 & io_in_x474_ready; // @[Math.scala 153:20:@4810.4]
  assign x487_sum_1_clock = clock; // @[:@4818.4]
  assign x487_sum_1_reset = reset; // @[:@4819.4]
  assign x487_sum_1_io_a = x485_sub_1_io_result; // @[Math.scala 151:17:@4820.4]
  assign x487_sum_1_io_b = 32'h12; // @[Math.scala 152:17:@4821.4]
  assign x487_sum_1_io_flow = _T_357 & io_in_x474_ready; // @[Math.scala 153:20:@4822.4]
  assign RetimeWrapper_2_clock = clock; // @[:@4847.4]
  assign RetimeWrapper_2_reset = reset; // @[:@4848.4]
  assign RetimeWrapper_2_io_flow = _T_357 & io_in_x474_ready; // @[package.scala 95:18:@4850.4]
  assign RetimeWrapper_2_io_in = _GEN_3 << 4; // @[package.scala 94:16:@4849.4]
  assign RetimeWrapper_3_clock = clock; // @[:@4859.4]
  assign RetimeWrapper_3_reset = reset; // @[:@4860.4]
  assign RetimeWrapper_3_io_flow = _T_357 & io_in_x474_ready; // @[package.scala 95:18:@4862.4]
  assign RetimeWrapper_3_io_in = _GEN_4 << 6; // @[package.scala 94:16:@4861.4]
  assign x491_1_io_b = _T_395[31:0]; // @[Math.scala 721:17:@4871.4]
  assign RetimeWrapper_4_clock = clock; // @[:@4879.4]
  assign RetimeWrapper_4_reset = reset; // @[:@4880.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4882.4]
  assign RetimeWrapper_4_io_in = io_in_x468_A_dram_number; // @[package.scala 94:16:@4881.4]
  assign x493_sum_1_clock = clock; // @[:@4888.4]
  assign x493_sum_1_reset = reset; // @[:@4889.4]
  assign x493_sum_1_io_a = x491_1_io_result; // @[Math.scala 151:17:@4890.4]
  assign x493_sum_1_io_b = RetimeWrapper_4_io_out; // @[Math.scala 152:17:@4891.4]
  assign x493_sum_1_io_flow = _T_357 & io_in_x474_ready; // @[Math.scala 153:20:@4892.4]
  assign RetimeWrapper_5_clock = clock; // @[:@4899.4]
  assign RetimeWrapper_5_reset = reset; // @[:@4900.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4902.4]
  assign RetimeWrapper_5_io_in = x493_sum_1_io_result; // @[package.scala 94:16:@4901.4]
  assign RetimeWrapper_6_clock = clock; // @[:@4913.4]
  assign RetimeWrapper_6_reset = reset; // @[:@4914.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4916.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@4915.4]
  assign RetimeWrapper_7_clock = clock; // @[:@4923.4]
  assign RetimeWrapper_7_reset = reset; // @[:@4924.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4926.4]
  assign RetimeWrapper_7_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@4925.4]
  assign RetimeWrapper_8_clock = clock; // @[:@4933.4]
  assign RetimeWrapper_8_reset = reset; // @[:@4934.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4936.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_datapathEn & io_sigsIn_iiIssue; // @[package.scala 94:16:@4935.4]
  assign RetimeWrapper_9_clock = clock; // @[:@4951.4]
  assign RetimeWrapper_9_reset = reset; // @[:@4952.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4954.4]
  assign RetimeWrapper_9_io_in = x486_sum_1_io_result; // @[package.scala 94:16:@4953.4]
  assign RetimeWrapper_10_clock = clock; // @[:@4961.4]
  assign RetimeWrapper_10_reset = reset; // @[:@4962.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4964.4]
  assign RetimeWrapper_10_io_in = x485_sub_1_io_result; // @[package.scala 94:16:@4963.4]
  assign RetimeWrapper_11_clock = clock; // @[:@4977.4]
  assign RetimeWrapper_11_reset = reset; // @[:@4978.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4980.4]
  assign RetimeWrapper_11_io_in = io_sigsIn_datapathEn & io_sigsIn_iiIssue; // @[package.scala 94:16:@4979.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_321 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_321 <= 1'h0;
    end else begin
      _T_321 <= _T_318;
    end
  end
endmodule
module x537_outr_Foreach_sm( // @[:@5333.2]
  input   clock, // @[:@5334.4]
  input   reset, // @[:@5335.4]
  input   io_enable, // @[:@5336.4]
  output  io_done, // @[:@5336.4]
  input   io_ctrDone, // @[:@5336.4]
  output  io_ctrInc, // @[:@5336.4]
  output  io_ctrRst, // @[:@5336.4]
  input   io_parentAck, // @[:@5336.4]
  input   io_doneIn_0, // @[:@5336.4]
  input   io_doneIn_1, // @[:@5336.4]
  input   io_maskIn_0, // @[:@5336.4]
  input   io_maskIn_1, // @[:@5336.4]
  output  io_enableOut_0, // @[:@5336.4]
  output  io_enableOut_1, // @[:@5336.4]
  output  io_childAck_0, // @[:@5336.4]
  output  io_childAck_1 // @[:@5336.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@5339.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@5339.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@5339.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@5339.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@5339.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@5339.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@5342.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@5342.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@5342.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@5342.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@5342.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@5342.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@5345.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@5345.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@5345.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@5345.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@5345.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@5345.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@5348.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@5348.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@5348.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@5348.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@5348.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@5348.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@5377.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@5377.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@5377.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@5377.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@5377.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@5377.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@5380.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@5380.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@5380.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@5380.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@5380.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@5380.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@5409.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@5409.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@5409.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@5409.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@5409.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@5505.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@5505.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@5505.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@5505.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@5505.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@5522.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@5522.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@5522.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@5522.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@5522.4]
  wire  allDone; // @[Controllers.scala 80:47:@5351.4]
  wire  _T_77; // @[Controllers.scala 81:26:@5352.4]
  wire  finished; // @[Controllers.scala 81:37:@5353.4]
  wire  _T_134; // @[package.scala 96:25:@5414.4 package.scala 96:25:@5415.4]
  wire  _T_138; // @[Controllers.scala 125:45:@5417.4]
  wire  _T_139; // @[Controllers.scala 125:61:@5418.4]
  wire  _T_140; // @[Controllers.scala 125:87:@5419.4]
  wire  synchronize; // @[Controllers.scala 125:42:@5421.4]
  wire  _T_144; // @[Controllers.scala 128:33:@5423.4]
  wire  _T_146; // @[Controllers.scala 128:54:@5424.4]
  wire  _T_147; // @[Controllers.scala 128:52:@5425.4]
  wire  _T_148; // @[Controllers.scala 128:66:@5426.4]
  wire  _T_150; // @[Controllers.scala 128:98:@5428.4]
  wire  _T_151; // @[Controllers.scala 128:96:@5429.4]
  wire  _T_153; // @[Controllers.scala 128:123:@5430.4]
  wire  _T_156; // @[Controllers.scala 129:57:@5434.4]
  wire  _T_160; // @[Controllers.scala 130:52:@5438.4]
  wire  _T_161; // @[Controllers.scala 130:50:@5439.4]
  wire  _T_163; // @[Controllers.scala 130:69:@5440.4]
  wire  _T_164; // @[Controllers.scala 130:83:@5441.4]
  wire  _T_166; // @[Controllers.scala 130:66:@5443.4]
  wire  _T_169; // @[Controllers.scala 130:129:@5445.4]
  wire  _T_175; // @[Controllers.scala 135:80:@5452.4]
  wire  _T_176; // @[Controllers.scala 135:78:@5453.4]
  wire  _T_178; // @[Controllers.scala 135:105:@5454.4]
  wire  _T_179; // @[Controllers.scala 135:103:@5455.4]
  wire  _T_180; // @[Controllers.scala 135:119:@5456.4]
  wire  _T_182; // @[Controllers.scala 135:51:@5458.4]
  wire  _T_191; // @[Controllers.scala 137:79:@5467.4]
  wire  _T_192; // @[Controllers.scala 137:95:@5468.4]
  wire  _T_194; // @[Controllers.scala 137:52:@5470.4]
  wire  _T_205; // @[Controllers.scala 213:68:@5483.4]
  wire  _T_207; // @[Controllers.scala 213:90:@5485.4]
  wire  _T_208; // @[Controllers.scala 213:115:@5486.4]
  wire  _T_209; // @[Controllers.scala 213:132:@5487.4]
  wire  _T_210; // @[Controllers.scala 213:130:@5488.4]
  wire  _T_211; // @[Controllers.scala 213:156:@5489.4]
  wire  _T_213; // @[Controllers.scala 213:68:@5492.4]
  wire  _T_215; // @[Controllers.scala 213:90:@5494.4]
  wire  _T_216; // @[Controllers.scala 213:115:@5495.4]
  wire  _T_222; // @[package.scala 100:49:@5500.4]
  reg  _T_225; // @[package.scala 48:56:@5501.4]
  reg [31:0] _RAND_0;
  wire  _T_226; // @[package.scala 100:41:@5503.4]
  reg  _T_239; // @[package.scala 48:56:@5519.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@5339.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@5342.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@5345.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@5348.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@5377.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@5380.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@5409.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@5505.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@5522.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@5351.4]
  assign _T_77 = allDone | io_done; // @[Controllers.scala 81:26:@5352.4]
  assign finished = _T_77 | done_1_io_input_set; // @[Controllers.scala 81:37:@5353.4]
  assign _T_134 = RetimeWrapper_io_out; // @[package.scala 96:25:@5414.4 package.scala 96:25:@5415.4]
  assign _T_138 = io_maskIn_1 == 1'h0; // @[Controllers.scala 125:45:@5417.4]
  assign _T_139 = _T_138 & iterDone_1_io_output; // @[Controllers.scala 125:61:@5418.4]
  assign _T_140 = _T_139 & io_enable; // @[Controllers.scala 125:87:@5419.4]
  assign synchronize = _T_134 | _T_140; // @[Controllers.scala 125:42:@5421.4]
  assign _T_144 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@5423.4]
  assign _T_146 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@5424.4]
  assign _T_147 = _T_144 & _T_146; // @[Controllers.scala 128:52:@5425.4]
  assign _T_148 = _T_147 & io_enable; // @[Controllers.scala 128:66:@5426.4]
  assign _T_150 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@5428.4]
  assign _T_151 = _T_148 & _T_150; // @[Controllers.scala 128:96:@5429.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@5430.4]
  assign _T_156 = io_doneIn_0 | io_parentAck; // @[Controllers.scala 129:57:@5434.4]
  assign _T_160 = synchronize == 1'h0; // @[Controllers.scala 130:52:@5438.4]
  assign _T_161 = io_doneIn_0 & _T_160; // @[Controllers.scala 130:50:@5439.4]
  assign _T_163 = io_maskIn_0 == 1'h0; // @[Controllers.scala 130:69:@5440.4]
  assign _T_164 = _T_163 & io_enable; // @[Controllers.scala 130:83:@5441.4]
  assign _T_166 = _T_161 | _T_164; // @[Controllers.scala 130:66:@5443.4]
  assign _T_169 = finished == 1'h0; // @[Controllers.scala 130:129:@5445.4]
  assign _T_175 = ~ iterDone_1_io_output; // @[Controllers.scala 135:80:@5452.4]
  assign _T_176 = iterDone_0_io_output & _T_175; // @[Controllers.scala 135:78:@5453.4]
  assign _T_178 = io_doneIn_1 == 1'h0; // @[Controllers.scala 135:105:@5454.4]
  assign _T_179 = _T_176 & _T_178; // @[Controllers.scala 135:103:@5455.4]
  assign _T_180 = _T_179 & io_enable; // @[Controllers.scala 135:119:@5456.4]
  assign _T_182 = io_doneIn_0 | _T_180; // @[Controllers.scala 135:51:@5458.4]
  assign _T_191 = iterDone_0_io_output & _T_138; // @[Controllers.scala 137:79:@5467.4]
  assign _T_192 = _T_191 & io_enable; // @[Controllers.scala 137:95:@5468.4]
  assign _T_194 = io_doneIn_1 | _T_192; // @[Controllers.scala 137:52:@5470.4]
  assign _T_205 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@5483.4]
  assign _T_207 = _T_205 & _T_150; // @[Controllers.scala 213:90:@5485.4]
  assign _T_208 = _T_207 & io_maskIn_0; // @[Controllers.scala 213:115:@5486.4]
  assign _T_209 = ~ allDone; // @[Controllers.scala 213:132:@5487.4]
  assign _T_210 = _T_208 & _T_209; // @[Controllers.scala 213:130:@5488.4]
  assign _T_211 = ~ io_ctrDone; // @[Controllers.scala 213:156:@5489.4]
  assign _T_213 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@5492.4]
  assign _T_215 = _T_213 & _T_175; // @[Controllers.scala 213:90:@5494.4]
  assign _T_216 = _T_215 & io_maskIn_1; // @[Controllers.scala 213:115:@5495.4]
  assign _T_222 = allDone == 1'h0; // @[package.scala 100:49:@5500.4]
  assign _T_226 = allDone & _T_225; // @[package.scala 100:41:@5503.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@5529.4]
  assign io_ctrInc = io_doneIn_1 | _T_140; // @[Controllers.scala 122:17:@5408.4]
  assign io_ctrRst = RetimeWrapper_1_io_out; // @[Controllers.scala 215:13:@5512.4]
  assign io_enableOut_0 = _T_210 & _T_211; // @[Controllers.scala 213:55:@5491.4]
  assign io_enableOut_1 = _T_216 & _T_209; // @[Controllers.scala 213:55:@5499.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@5480.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@5482.4]
  assign active_0_clock = clock; // @[:@5340.4]
  assign active_0_reset = reset; // @[:@5341.4]
  assign active_0_io_input_set = _T_151 & _T_153; // @[Controllers.scala 128:30:@5432.4]
  assign active_0_io_input_reset = _T_156 | allDone; // @[Controllers.scala 129:32:@5437.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@5354.4]
  assign active_1_clock = clock; // @[:@5343.4]
  assign active_1_reset = reset; // @[:@5344.4]
  assign active_1_io_input_set = _T_182 & _T_160; // @[Controllers.scala 135:32:@5461.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 136:34:@5465.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@5355.4]
  assign done_0_clock = clock; // @[:@5346.4]
  assign done_0_reset = reset; // @[:@5347.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 131:28:@5451.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@5366.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@5356.4]
  assign done_1_clock = clock; // @[:@5349.4]
  assign done_1_reset = reset; // @[:@5350.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 138:30:@5478.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@5375.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@5357.4]
  assign iterDone_0_clock = clock; // @[:@5378.4]
  assign iterDone_0_reset = reset; // @[:@5379.4]
  assign iterDone_0_io_input_set = _T_166 & _T_169; // @[Controllers.scala 130:32:@5447.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@5393.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@5383.4]
  assign iterDone_1_clock = clock; // @[:@5381.4]
  assign iterDone_1_reset = reset; // @[:@5382.4]
  assign iterDone_1_io_input_set = _T_194 & _T_160; // @[Controllers.scala 137:34:@5474.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@5402.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@5384.4]
  assign RetimeWrapper_clock = clock; // @[:@5410.4]
  assign RetimeWrapper_reset = reset; // @[:@5411.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@5413.4]
  assign RetimeWrapper_io_in = io_doneIn_1; // @[package.scala 94:16:@5412.4]
  assign RetimeWrapper_1_clock = clock; // @[:@5506.4]
  assign RetimeWrapper_1_reset = reset; // @[:@5507.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@5509.4]
  assign RetimeWrapper_1_io_in = _T_226 | io_parentAck; // @[package.scala 94:16:@5508.4]
  assign RetimeWrapper_2_clock = clock; // @[:@5523.4]
  assign RetimeWrapper_2_reset = reset; // @[:@5524.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@5526.4]
  assign RetimeWrapper_2_io_in = allDone & _T_239; // @[package.scala 94:16:@5525.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_225 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_239 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_225 <= 1'h0;
    end else begin
      _T_225 <= _T_222;
    end
    if (reset) begin
      _T_239 <= 1'h0;
    end else begin
      _T_239 <= _T_222;
    end
  end
endmodule
module x505_reg( // @[:@5709.2]
  input         clock, // @[:@5710.4]
  input         reset, // @[:@5711.4]
  output [31:0] io_rPort_0_output_0, // @[:@5712.4]
  input  [31:0] io_wPort_0_data_0, // @[:@5712.4]
  input         io_wPort_0_reset, // @[:@5712.4]
  input         io_wPort_0_en_0 // @[:@5712.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@5728.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 325:32:@5730.4]
  wire [31:0] _T_70; // @[MemPrimitives.scala 325:12:@5731.4]
  assign _T_69 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@5730.4]
  assign _T_70 = io_wPort_0_reset ? 32'h0 : _T_69; // @[MemPrimitives.scala 325:12:@5731.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@5733.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module x516_inr_UnitPipe_sm( // @[:@5941.2]
  input   clock, // @[:@5942.4]
  input   reset, // @[:@5943.4]
  input   io_enable, // @[:@5944.4]
  output  io_done, // @[:@5944.4]
  output  io_doneLatch, // @[:@5944.4]
  input   io_ctrDone, // @[:@5944.4]
  output  io_datapathEn, // @[:@5944.4]
  output  io_ctrInc, // @[:@5944.4]
  input   io_parentAck, // @[:@5944.4]
  input   io_backpressure, // @[:@5944.4]
  input   io_break // @[:@5944.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@5946.4]
  wire  active_reset; // @[Controllers.scala 261:22:@5946.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@5946.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@5946.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@5946.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@5946.4]
  wire  done_clock; // @[Controllers.scala 262:20:@5949.4]
  wire  done_reset; // @[Controllers.scala 262:20:@5949.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@5949.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@5949.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@5949.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@5949.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@5983.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@5983.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@5983.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@5983.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@5983.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6005.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6005.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6005.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6005.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6005.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6017.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6017.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6017.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6017.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6017.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6025.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6025.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6025.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6025.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6025.4]
  wire  _T_80; // @[Controllers.scala 264:48:@5954.4]
  wire  _T_81; // @[Controllers.scala 264:46:@5955.4]
  wire  _T_82; // @[Controllers.scala 264:62:@5956.4]
  wire  _T_100; // @[package.scala 100:49:@5974.4]
  reg  _T_103; // @[package.scala 48:56:@5975.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@5998.4]
  wire  _T_124; // @[package.scala 96:25:@6010.4 package.scala 96:25:@6011.4]
  wire  _T_126; // @[package.scala 100:49:@6012.4]
  reg  _T_129; // @[package.scala 48:56:@6013.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@6035.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@6037.4]
  reg  _T_153; // @[package.scala 48:56:@6038.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@6040.4]
  wire  _T_156; // @[Controllers.scala 292:61:@6041.4]
  wire  _T_157; // @[Controllers.scala 292:24:@6042.4]
  SRFF active ( // @[Controllers.scala 261:22:@5946.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@5949.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@5983.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@6005.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6017.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6025.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@5954.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@5955.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@5956.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@5974.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@5998.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6010.4 package.scala 96:25:@6011.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@6012.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@6037.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@6040.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@6041.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@6042.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@6016.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@6044.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@6001.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@6004.4]
  assign active_clock = clock; // @[:@5947.4]
  assign active_reset = reset; // @[:@5948.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@5959.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@5963.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@5964.4]
  assign done_clock = clock; // @[:@5950.4]
  assign done_reset = reset; // @[:@5951.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@5979.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@5972.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@5973.4]
  assign RetimeWrapper_clock = clock; // @[:@5984.4]
  assign RetimeWrapper_reset = reset; // @[:@5985.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@5987.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@5986.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6006.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6007.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@6009.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@6008.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6018.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6019.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6021.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@6020.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6026.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6027.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6029.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@6028.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1( // @[:@6167.2]
  input         clock, // @[:@6168.4]
  input         reset, // @[:@6169.4]
  output        io_in_x475_fifo_rPort_0_en_0, // @[:@6170.4]
  input  [95:0] io_in_x475_fifo_rPort_0_output_0, // @[:@6170.4]
  input         io_in_x475_fifo_empty, // @[:@6170.4]
  output [31:0] io_in_x507_reg_wPort_0_data_0, // @[:@6170.4]
  output        io_in_x507_reg_wPort_0_reset, // @[:@6170.4]
  output        io_in_x507_reg_wPort_0_en_0, // @[:@6170.4]
  output        io_in_x507_reg_reset, // @[:@6170.4]
  output [31:0] io_in_x505_reg_wPort_0_data_0, // @[:@6170.4]
  output        io_in_x505_reg_wPort_0_reset, // @[:@6170.4]
  output        io_in_x505_reg_wPort_0_en_0, // @[:@6170.4]
  output        io_in_x505_reg_reset, // @[:@6170.4]
  output [31:0] io_in_x506_reg_wPort_0_data_0, // @[:@6170.4]
  output        io_in_x506_reg_wPort_0_reset, // @[:@6170.4]
  output        io_in_x506_reg_wPort_0_en_0, // @[:@6170.4]
  output        io_in_x506_reg_reset, // @[:@6170.4]
  output [63:0] io_in_instrctrs_4_cycs, // @[:@6170.4]
  output [63:0] io_in_instrctrs_4_iters, // @[:@6170.4]
  output [63:0] io_in_instrctrs_4_stalls, // @[:@6170.4]
  output [63:0] io_in_instrctrs_4_idles, // @[:@6170.4]
  input         io_sigsIn_done, // @[:@6170.4]
  input         io_sigsIn_forwardpressure, // @[:@6170.4]
  input         io_sigsIn_datapathEn, // @[:@6170.4]
  input         io_sigsIn_baseEn, // @[:@6170.4]
  input         io_sigsIn_break, // @[:@6170.4]
  input         io_rr // @[:@6170.4]
);
  wire  cycles_x516_inr_UnitPipe_clock; // @[sm_x516_inr_UnitPipe.scala 76:44:@6337.4]
  wire  cycles_x516_inr_UnitPipe_reset; // @[sm_x516_inr_UnitPipe.scala 76:44:@6337.4]
  wire  cycles_x516_inr_UnitPipe_io_enable; // @[sm_x516_inr_UnitPipe.scala 76:44:@6337.4]
  wire [63:0] cycles_x516_inr_UnitPipe_io_count; // @[sm_x516_inr_UnitPipe.scala 76:44:@6337.4]
  wire  iters_x516_inr_UnitPipe_clock; // @[sm_x516_inr_UnitPipe.scala 77:43:@6340.4]
  wire  iters_x516_inr_UnitPipe_reset; // @[sm_x516_inr_UnitPipe.scala 77:43:@6340.4]
  wire  iters_x516_inr_UnitPipe_io_enable; // @[sm_x516_inr_UnitPipe.scala 77:43:@6340.4]
  wire [63:0] iters_x516_inr_UnitPipe_io_count; // @[sm_x516_inr_UnitPipe.scala 77:43:@6340.4]
  wire  stalls_x516_inr_UnitPipe_clock; // @[sm_x516_inr_UnitPipe.scala 80:44:@6349.4]
  wire  stalls_x516_inr_UnitPipe_reset; // @[sm_x516_inr_UnitPipe.scala 80:44:@6349.4]
  wire  stalls_x516_inr_UnitPipe_io_enable; // @[sm_x516_inr_UnitPipe.scala 80:44:@6349.4]
  wire [63:0] stalls_x516_inr_UnitPipe_io_count; // @[sm_x516_inr_UnitPipe.scala 80:44:@6349.4]
  wire  idles_x516_inr_UnitPipe_clock; // @[sm_x516_inr_UnitPipe.scala 81:43:@6352.4]
  wire  idles_x516_inr_UnitPipe_reset; // @[sm_x516_inr_UnitPipe.scala 81:43:@6352.4]
  wire  idles_x516_inr_UnitPipe_io_enable; // @[sm_x516_inr_UnitPipe.scala 81:43:@6352.4]
  wire [63:0] idles_x516_inr_UnitPipe_io_count; // @[sm_x516_inr_UnitPipe.scala 81:43:@6352.4]
  wire  _T_690; // @[package.scala 100:49:@6344.4]
  reg  _T_693; // @[package.scala 48:56:@6345.4]
  reg [31:0] _RAND_0;
  wire  _T_702; // @[sm_x516_inr_UnitPipe.scala 83:67:@6359.4]
  wire  _T_707; // @[sm_x516_inr_UnitPipe.scala 83:63:@6363.4]
  wire  _T_718; // @[implicits.scala 56:10:@6372.4]
  wire  _T_719; // @[sm_x516_inr_UnitPipe.scala 89:120:@6373.4]
  wire  _T_720; // @[sm_x516_inr_UnitPipe.scala 89:117:@6374.4]
  wire  _T_725; // @[implicits.scala 56:10:@6377.4]
  wire  _T_740; // @[sm_x516_inr_UnitPipe.scala 101:133:@6395.4]
  InstrumentationCounter cycles_x516_inr_UnitPipe ( // @[sm_x516_inr_UnitPipe.scala 76:44:@6337.4]
    .clock(cycles_x516_inr_UnitPipe_clock),
    .reset(cycles_x516_inr_UnitPipe_reset),
    .io_enable(cycles_x516_inr_UnitPipe_io_enable),
    .io_count(cycles_x516_inr_UnitPipe_io_count)
  );
  InstrumentationCounter iters_x516_inr_UnitPipe ( // @[sm_x516_inr_UnitPipe.scala 77:43:@6340.4]
    .clock(iters_x516_inr_UnitPipe_clock),
    .reset(iters_x516_inr_UnitPipe_reset),
    .io_enable(iters_x516_inr_UnitPipe_io_enable),
    .io_count(iters_x516_inr_UnitPipe_io_count)
  );
  InstrumentationCounter stalls_x516_inr_UnitPipe ( // @[sm_x516_inr_UnitPipe.scala 80:44:@6349.4]
    .clock(stalls_x516_inr_UnitPipe_clock),
    .reset(stalls_x516_inr_UnitPipe_reset),
    .io_enable(stalls_x516_inr_UnitPipe_io_enable),
    .io_count(stalls_x516_inr_UnitPipe_io_count)
  );
  InstrumentationCounter idles_x516_inr_UnitPipe ( // @[sm_x516_inr_UnitPipe.scala 81:43:@6352.4]
    .clock(idles_x516_inr_UnitPipe_clock),
    .reset(idles_x516_inr_UnitPipe_reset),
    .io_enable(idles_x516_inr_UnitPipe_io_enable),
    .io_count(idles_x516_inr_UnitPipe_io_count)
  );
  assign _T_690 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@6344.4]
  assign _T_702 = ~ io_in_x475_fifo_empty; // @[sm_x516_inr_UnitPipe.scala 83:67:@6359.4]
  assign _T_707 = ~ _T_702; // @[sm_x516_inr_UnitPipe.scala 83:63:@6363.4]
  assign _T_718 = io_rr ? io_sigsIn_forwardpressure : 1'h0; // @[implicits.scala 56:10:@6372.4]
  assign _T_719 = ~ io_sigsIn_break; // @[sm_x516_inr_UnitPipe.scala 89:120:@6373.4]
  assign _T_720 = _T_718 & _T_719; // @[sm_x516_inr_UnitPipe.scala 89:117:@6374.4]
  assign _T_725 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 56:10:@6377.4]
  assign _T_740 = _T_719 & _T_725; // @[sm_x516_inr_UnitPipe.scala 101:133:@6395.4]
  assign io_in_x475_fifo_rPort_0_en_0 = _T_720 & _T_725; // @[MemInterfaceType.scala 110:79:@6382.4]
  assign io_in_x507_reg_wPort_0_data_0 = io_in_x475_fifo_rPort_0_output_0[31:0]; // @[MemInterfaceType.scala 90:56:@6432.4]
  assign io_in_x507_reg_wPort_0_reset = io_in_x507_reg_reset; // @[MemInterfaceType.scala 91:23:@6433.4]
  assign io_in_x507_reg_wPort_0_en_0 = _T_740 & _T_719; // @[MemInterfaceType.scala 93:57:@6434.4]
  assign io_in_x507_reg_reset = 1'h0;
  assign io_in_x505_reg_wPort_0_data_0 = io_in_x475_fifo_rPort_0_output_0[63:32]; // @[MemInterfaceType.scala 90:56:@6400.4]
  assign io_in_x505_reg_wPort_0_reset = io_in_x505_reg_reset; // @[MemInterfaceType.scala 91:23:@6401.4]
  assign io_in_x505_reg_wPort_0_en_0 = _T_740 & _T_719; // @[MemInterfaceType.scala 93:57:@6402.4]
  assign io_in_x505_reg_reset = 1'h0;
  assign io_in_x506_reg_wPort_0_data_0 = io_in_x475_fifo_rPort_0_output_0[95:64]; // @[MemInterfaceType.scala 90:56:@6416.4]
  assign io_in_x506_reg_wPort_0_reset = io_in_x506_reg_reset; // @[MemInterfaceType.scala 91:23:@6417.4]
  assign io_in_x506_reg_wPort_0_en_0 = _T_740 & _T_719; // @[MemInterfaceType.scala 93:57:@6418.4]
  assign io_in_x506_reg_reset = 1'h0;
  assign io_in_instrctrs_4_cycs = cycles_x516_inr_UnitPipe_io_count; // @[Ledger.scala 293:21:@6366.4]
  assign io_in_instrctrs_4_iters = iters_x516_inr_UnitPipe_io_count; // @[Ledger.scala 294:22:@6367.4]
  assign io_in_instrctrs_4_stalls = stalls_x516_inr_UnitPipe_io_count; // @[Ledger.scala 295:23:@6368.4]
  assign io_in_instrctrs_4_idles = idles_x516_inr_UnitPipe_io_count; // @[Ledger.scala 296:22:@6369.4]
  assign cycles_x516_inr_UnitPipe_clock = clock; // @[:@6338.4]
  assign cycles_x516_inr_UnitPipe_reset = reset; // @[:@6339.4]
  assign cycles_x516_inr_UnitPipe_io_enable = io_sigsIn_baseEn; // @[sm_x516_inr_UnitPipe.scala 78:42:@6343.4]
  assign iters_x516_inr_UnitPipe_clock = clock; // @[:@6341.4]
  assign iters_x516_inr_UnitPipe_reset = reset; // @[:@6342.4]
  assign iters_x516_inr_UnitPipe_io_enable = io_sigsIn_done & _T_693; // @[sm_x516_inr_UnitPipe.scala 79:41:@6348.4]
  assign stalls_x516_inr_UnitPipe_clock = clock; // @[:@6350.4]
  assign stalls_x516_inr_UnitPipe_reset = reset; // @[:@6351.4]
  assign stalls_x516_inr_UnitPipe_io_enable = 1'h0; // @[sm_x516_inr_UnitPipe.scala 82:42:@6357.4]
  assign idles_x516_inr_UnitPipe_clock = clock; // @[:@6353.4]
  assign idles_x516_inr_UnitPipe_reset = reset; // @[:@6354.4]
  assign idles_x516_inr_UnitPipe_io_enable = io_sigsIn_baseEn & _T_707; // @[sm_x516_inr_UnitPipe.scala 83:41:@6365.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_693 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_693 <= 1'h0;
    end else begin
      _T_693 <= _T_690;
    end
  end
endmodule
module SingleCounter_3( // @[:@6474.2]
  input         clock, // @[:@6475.4]
  input         reset, // @[:@6476.4]
  input  [31:0] io_setup_stop, // @[:@6477.4]
  input         io_setup_saturate, // @[:@6477.4]
  input         io_input_reset, // @[:@6477.4]
  input         io_input_enable, // @[:@6477.4]
  output [31:0] io_output_count_0, // @[:@6477.4]
  output        io_output_oobs_0, // @[:@6477.4]
  output        io_output_noop, // @[:@6477.4]
  output        io_output_done // @[:@6477.4]
);
  wire  bases_0_clock; // @[Counter.scala 262:53:@6490.4]
  wire  bases_0_reset; // @[Counter.scala 262:53:@6490.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 262:53:@6490.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 262:53:@6490.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 262:53:@6490.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 262:53:@6490.4]
  wire  SRFF_clock; // @[Counter.scala 264:22:@6506.4]
  wire  SRFF_reset; // @[Counter.scala 264:22:@6506.4]
  wire  SRFF_io_input_set; // @[Counter.scala 264:22:@6506.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 264:22:@6506.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 264:22:@6506.4]
  wire  SRFF_io_output; // @[Counter.scala 264:22:@6506.4]
  wire  _T_36; // @[Counter.scala 265:45:@6509.4]
  wire [31:0] _T_48; // @[Counter.scala 288:52:@6534.4]
  wire [32:0] _T_50; // @[Counter.scala 292:33:@6535.4]
  wire [31:0] _T_51; // @[Counter.scala 292:33:@6536.4]
  wire [31:0] _T_52; // @[Counter.scala 292:33:@6537.4]
  wire  _T_56; // @[Counter.scala 294:18:@6539.4]
  wire [31:0] _T_66; // @[Counter.scala 300:115:@6547.4]
  wire [31:0] _T_68; // @[Counter.scala 300:85:@6549.4]
  wire [31:0] _T_69; // @[Counter.scala 300:152:@6550.4]
  wire [31:0] _T_70; // @[Counter.scala 300:74:@6551.4]
  wire  _T_73; // @[Counter.scala 325:102:@6555.4]
  wire  _T_74; // @[Counter.scala 325:130:@6556.4]
  FF bases_0 ( // @[Counter.scala 262:53:@6490.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 264:22:@6506.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 265:45:@6509.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 288:52:@6534.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 292:33:@6535.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 292:33:@6536.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 292:33:@6537.4]
  assign _T_56 = $signed(_T_52) >= $signed(io_setup_stop); // @[Counter.scala 294:18:@6539.4]
  assign _T_66 = $unsigned(_T_48); // @[Counter.scala 300:115:@6547.4]
  assign _T_68 = io_setup_saturate ? _T_66 : 32'h0; // @[Counter.scala 300:85:@6549.4]
  assign _T_69 = $unsigned(_T_52); // @[Counter.scala 300:152:@6550.4]
  assign _T_70 = _T_56 ? _T_68 : _T_69; // @[Counter.scala 300:74:@6551.4]
  assign _T_73 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 325:102:@6555.4]
  assign _T_74 = $signed(_T_48) >= $signed(io_setup_stop); // @[Counter.scala 325:130:@6556.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 305:28:@6554.4]
  assign io_output_oobs_0 = _T_73 | _T_74; // @[Counter.scala 325:60:@6558.4]
  assign io_output_noop = $signed(32'sh0) == $signed(io_setup_stop); // @[Counter.scala 337:40:@6562.4]
  assign io_output_done = io_input_enable & _T_56; // @[Counter.scala 334:20:@6560.4]
  assign bases_0_clock = clock; // @[:@6491.4]
  assign bases_0_reset = reset; // @[:@6492.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_70; // @[Counter.scala 300:31:@6553.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 282:27:@6532.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 285:29:@6533.4]
  assign SRFF_clock = clock; // @[:@6507.4]
  assign SRFF_reset = reset; // @[:@6508.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 265:23:@6511.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 266:25:@6513.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 267:30:@6514.4]
endmodule
module x519_ctrchain( // @[:@6566.2]
  input         clock, // @[:@6567.4]
  input         reset, // @[:@6568.4]
  input  [31:0] io_setup_stops_0, // @[:@6569.4]
  input         io_input_reset, // @[:@6569.4]
  input         io_input_enable, // @[:@6569.4]
  output [31:0] io_output_counts_0, // @[:@6569.4]
  output        io_output_oobs_0, // @[:@6569.4]
  output        io_output_noop, // @[:@6569.4]
  output        io_output_done // @[:@6569.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 514:46:@6571.4]
  wire  ctrs_0_reset; // @[Counter.scala 514:46:@6571.4]
  wire [31:0] ctrs_0_io_setup_stop; // @[Counter.scala 514:46:@6571.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 514:46:@6571.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 514:46:@6571.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 514:46:@6571.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 514:46:@6571.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 514:46:@6571.4]
  wire  ctrs_0_io_output_noop; // @[Counter.scala 514:46:@6571.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 514:46:@6571.4]
  reg  wasDone; // @[Counter.scala 543:24:@6580.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 547:69:@6586.4]
  wire  _T_47; // @[Counter.scala 547:80:@6587.4]
  reg  doneLatch; // @[Counter.scala 551:26:@6592.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 552:48:@6593.4]
  wire  _T_55; // @[Counter.scala 552:19:@6594.4]
  SingleCounter_3 ctrs_0 ( // @[Counter.scala 514:46:@6571.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_stop(ctrs_0_io_setup_stop),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_noop(ctrs_0_io_output_noop),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 547:69:@6586.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 547:80:@6587.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 552:48:@6593.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 552:19:@6594.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 558:32:@6596.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 559:30:@6598.4]
  assign io_output_noop = ctrs_0_io_output_noop; // @[Counter.scala 546:18:@6584.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 547:18:@6589.4]
  assign ctrs_0_clock = clock; // @[:@6572.4]
  assign ctrs_0_reset = reset; // @[:@6573.4]
  assign ctrs_0_io_setup_stop = io_setup_stops_0; // @[Counter.scala 519:23:@6575.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 531:29:@6579.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 521:24:@6577.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 525:33:@6578.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_59( // @[:@6638.2]
  input   clock, // @[:@6639.4]
  input   reset, // @[:@6640.4]
  input   io_flow, // @[:@6641.4]
  input   io_in, // @[:@6641.4]
  output  io_out // @[:@6641.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6643.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6643.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6643.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6643.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6643.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6643.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@6643.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6656.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6655.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6654.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6653.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6652.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6650.4]
endmodule
module x536_inr_Foreach_sm( // @[:@6786.2]
  input   clock, // @[:@6787.4]
  input   reset, // @[:@6788.4]
  input   io_enable, // @[:@6789.4]
  output  io_done, // @[:@6789.4]
  output  io_doneLatch, // @[:@6789.4]
  input   io_ctrDone, // @[:@6789.4]
  output  io_datapathEn, // @[:@6789.4]
  output  io_ctrInc, // @[:@6789.4]
  output  io_ctrRst, // @[:@6789.4]
  input   io_parentAck, // @[:@6789.4]
  input   io_backpressure, // @[:@6789.4]
  input   io_break // @[:@6789.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@6791.4]
  wire  active_reset; // @[Controllers.scala 261:22:@6791.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@6791.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@6791.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@6791.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@6791.4]
  wire  done_clock; // @[Controllers.scala 262:20:@6794.4]
  wire  done_reset; // @[Controllers.scala 262:20:@6794.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@6794.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@6794.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@6794.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@6794.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6828.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6828.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6828.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6828.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6828.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6850.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6850.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6850.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6850.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6850.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6862.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6862.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6862.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6862.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6862.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6870.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6870.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6870.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6870.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6870.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@6886.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@6886.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@6886.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@6886.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@6886.4]
  wire  _T_80; // @[Controllers.scala 264:48:@6799.4]
  wire  _T_81; // @[Controllers.scala 264:46:@6800.4]
  wire  _T_82; // @[Controllers.scala 264:62:@6801.4]
  wire  _T_100; // @[package.scala 100:49:@6819.4]
  reg  _T_103; // @[package.scala 48:56:@6820.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@6833.4 package.scala 96:25:@6834.4]
  wire  _T_110; // @[package.scala 100:49:@6835.4]
  reg  _T_113; // @[package.scala 48:56:@6836.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@6838.4]
  wire  _T_118; // @[Controllers.scala 283:41:@6843.4]
  wire  _T_124; // @[package.scala 96:25:@6855.4 package.scala 96:25:@6856.4]
  wire  _T_126; // @[package.scala 100:49:@6857.4]
  reg  _T_129; // @[package.scala 48:56:@6858.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@6880.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@6882.4]
  reg  _T_153; // @[package.scala 48:56:@6883.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@6891.4 package.scala 96:25:@6892.4]
  wire  _T_158; // @[Controllers.scala 292:61:@6893.4]
  wire  _T_159; // @[Controllers.scala 292:24:@6894.4]
  SRFF active ( // @[Controllers.scala 261:22:@6791.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@6794.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_59 RetimeWrapper ( // @[package.scala 93:22:@6828.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_59 RetimeWrapper_1 ( // @[package.scala 93:22:@6850.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6862.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6870.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@6886.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@6799.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@6800.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@6801.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@6819.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@6833.4 package.scala 96:25:@6834.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@6835.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@6838.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@6843.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6855.4 package.scala 96:25:@6856.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@6857.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@6882.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@6891.4 package.scala 96:25:@6892.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@6893.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@6894.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@6861.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@6896.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@6846.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@6849.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@6841.4]
  assign active_clock = clock; // @[:@6792.4]
  assign active_reset = reset; // @[:@6793.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@6804.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@6808.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@6809.4]
  assign done_clock = clock; // @[:@6795.4]
  assign done_reset = reset; // @[:@6796.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@6824.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@6817.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@6818.4]
  assign RetimeWrapper_clock = clock; // @[:@6829.4]
  assign RetimeWrapper_reset = reset; // @[:@6830.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@6832.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@6831.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6851.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6852.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@6854.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@6853.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6863.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6864.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6866.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@6865.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6871.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6872.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6874.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@6873.4]
  assign RetimeWrapper_4_clock = clock; // @[:@6887.4]
  assign RetimeWrapper_4_reset = reset; // @[:@6888.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@6890.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@6889.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x536_inr_Foreach_kernelx536_inr_Foreach_concrete1( // @[:@7916.2]
  input         clock, // @[:@7917.4]
  input         reset, // @[:@7918.4]
  output [8:0]  io_in_x472_A_sram_1_wPort_0_ofs_0, // @[:@7919.4]
  output [31:0] io_in_x472_A_sram_1_wPort_0_data_0, // @[:@7919.4]
  output        io_in_x472_A_sram_1_wPort_0_en_0, // @[:@7919.4]
  input         io_in_b504, // @[:@7919.4]
  output [8:0]  io_in_x471_A_sram_0_wPort_0_ofs_0, // @[:@7919.4]
  output [31:0] io_in_x471_A_sram_0_wPort_0_data_0, // @[:@7919.4]
  output        io_in_x471_A_sram_0_wPort_0_en_0, // @[:@7919.4]
  output        io_in_x476_ready, // @[:@7919.4]
  input         io_in_x476_valid, // @[:@7919.4]
  input  [31:0] io_in_x476_bits_rdata_0, // @[:@7919.4]
  input  [31:0] io_in_b503_number, // @[:@7919.4]
  input  [31:0] io_in_x505_reg_rPort_0_output_0, // @[:@7919.4]
  output [8:0]  io_in_x473_A_sram_2_wPort_0_ofs_0, // @[:@7919.4]
  output [31:0] io_in_x473_A_sram_2_wPort_0_data_0, // @[:@7919.4]
  output        io_in_x473_A_sram_2_wPort_0_en_0, // @[:@7919.4]
  input  [31:0] io_in_x506_reg_rPort_0_output_0, // @[:@7919.4]
  output [63:0] io_in_instrctrs_5_cycs, // @[:@7919.4]
  output [63:0] io_in_instrctrs_5_iters, // @[:@7919.4]
  output [63:0] io_in_instrctrs_5_stalls, // @[:@7919.4]
  output [63:0] io_in_instrctrs_5_idles, // @[:@7919.4]
  input         io_sigsIn_done, // @[:@7919.4]
  input         io_sigsIn_datapathEn, // @[:@7919.4]
  input         io_sigsIn_baseEn, // @[:@7919.4]
  input         io_sigsIn_break, // @[:@7919.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@7919.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@7919.4]
  input         io_rr // @[:@7919.4]
);
  wire  cycles_x536_inr_Foreach_clock; // @[sm_x536_inr_Foreach.scala 89:43:@8090.4]
  wire  cycles_x536_inr_Foreach_reset; // @[sm_x536_inr_Foreach.scala 89:43:@8090.4]
  wire  cycles_x536_inr_Foreach_io_enable; // @[sm_x536_inr_Foreach.scala 89:43:@8090.4]
  wire [63:0] cycles_x536_inr_Foreach_io_count; // @[sm_x536_inr_Foreach.scala 89:43:@8090.4]
  wire  iters_x536_inr_Foreach_clock; // @[sm_x536_inr_Foreach.scala 90:42:@8093.4]
  wire  iters_x536_inr_Foreach_reset; // @[sm_x536_inr_Foreach.scala 90:42:@8093.4]
  wire  iters_x536_inr_Foreach_io_enable; // @[sm_x536_inr_Foreach.scala 90:42:@8093.4]
  wire [63:0] iters_x536_inr_Foreach_io_count; // @[sm_x536_inr_Foreach.scala 90:42:@8093.4]
  wire  stalls_x536_inr_Foreach_clock; // @[sm_x536_inr_Foreach.scala 93:43:@8102.4]
  wire  stalls_x536_inr_Foreach_reset; // @[sm_x536_inr_Foreach.scala 93:43:@8102.4]
  wire  stalls_x536_inr_Foreach_io_enable; // @[sm_x536_inr_Foreach.scala 93:43:@8102.4]
  wire [63:0] stalls_x536_inr_Foreach_io_count; // @[sm_x536_inr_Foreach.scala 93:43:@8102.4]
  wire  idles_x536_inr_Foreach_clock; // @[sm_x536_inr_Foreach.scala 94:42:@8105.4]
  wire  idles_x536_inr_Foreach_reset; // @[sm_x536_inr_Foreach.scala 94:42:@8105.4]
  wire  idles_x536_inr_Foreach_io_enable; // @[sm_x536_inr_Foreach.scala 94:42:@8105.4]
  wire [63:0] idles_x536_inr_Foreach_io_count; // @[sm_x536_inr_Foreach.scala 94:42:@8105.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@8123.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@8123.4]
  wire  x527_sub_1_clock; // @[Math.scala 191:24:@8174.4]
  wire  x527_sub_1_reset; // @[Math.scala 191:24:@8174.4]
  wire [31:0] x527_sub_1_io_a; // @[Math.scala 191:24:@8174.4]
  wire [31:0] x527_sub_1_io_b; // @[Math.scala 191:24:@8174.4]
  wire  x527_sub_1_io_flow; // @[Math.scala 191:24:@8174.4]
  wire [31:0] x527_sub_1_io_result; // @[Math.scala 191:24:@8174.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@8190.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@8190.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@8190.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@8190.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@8190.4]
  wire  x743_sum_1_clock; // @[Math.scala 150:24:@8206.4]
  wire  x743_sum_1_reset; // @[Math.scala 150:24:@8206.4]
  wire [31:0] x743_sum_1_io_a; // @[Math.scala 150:24:@8206.4]
  wire [31:0] x743_sum_1_io_b; // @[Math.scala 150:24:@8206.4]
  wire  x743_sum_1_io_flow; // @[Math.scala 150:24:@8206.4]
  wire [31:0] x743_sum_1_io_result; // @[Math.scala 150:24:@8206.4]
  wire  x532_sum_1_clock; // @[Math.scala 150:24:@8216.4]
  wire  x532_sum_1_reset; // @[Math.scala 150:24:@8216.4]
  wire [31:0] x532_sum_1_io_a; // @[Math.scala 150:24:@8216.4]
  wire [31:0] x532_sum_1_io_b; // @[Math.scala 150:24:@8216.4]
  wire  x532_sum_1_io_flow; // @[Math.scala 150:24:@8216.4]
  wire [31:0] x532_sum_1_io_result; // @[Math.scala 150:24:@8216.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@8227.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@8227.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@8227.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@8227.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@8227.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@8237.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@8237.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@8237.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@8237.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@8237.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@8247.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@8247.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@8247.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@8247.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@8247.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@8257.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@8257.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@8257.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@8257.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@8257.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@8271.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@8271.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@8271.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@8271.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@8271.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@8297.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@8297.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@8297.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@8297.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@8297.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@8323.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@8323.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@8323.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@8323.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@8323.4]
  wire  _T_782; // @[package.scala 100:49:@8097.4]
  reg  _T_785; // @[package.scala 48:56:@8098.4]
  reg [31:0] _RAND_0;
  wire  _T_792; // @[sm_x536_inr_Foreach.scala 96:62:@8112.4]
  wire  b521; // @[sm_x536_inr_Foreach.scala 99:18:@8131.4]
  wire  _T_806; // @[sm_x536_inr_Foreach.scala 104:119:@8135.4]
  wire [31:0] _T_818; // @[Math.scala 493:37:@8147.4]
  wire [31:0] b520_number; // @[Math.scala 723:22:@8128.4 Math.scala 724:14:@8129.4]
  wire [31:0] _T_819; // @[Math.scala 493:51:@8148.4]
  wire  x523; // @[Math.scala 493:44:@8149.4]
  wire [31:0] _T_839; // @[Math.scala 476:50:@8167.4]
  wire  x525; // @[Math.scala 476:44:@8168.4]
  wire  _T_853; // @[sm_x536_inr_Foreach.scala 121:26:@8184.4]
  wire [32:0] _GEN_0; // @[Math.scala 461:32:@8202.4]
  wire [32:0] _T_869; // @[Math.scala 461:32:@8202.4]
  wire  _T_908; // @[package.scala 96:25:@8276.4 package.scala 96:25:@8277.4]
  wire  _T_910; // @[implicits.scala 56:10:@8278.4]
  wire  _T_911; // @[sm_x536_inr_Foreach.scala 146:118:@8279.4]
  wire  _T_913; // @[sm_x536_inr_Foreach.scala 146:215:@8281.4]
  wire  x767_x526_D2; // @[package.scala 96:25:@8252.4 package.scala 96:25:@8253.4]
  wire  _T_915; // @[sm_x536_inr_Foreach.scala 146:260:@8283.4]
  wire  x768_b521_D2; // @[package.scala 96:25:@8262.4 package.scala 96:25:@8263.4]
  wire  _T_916; // @[sm_x536_inr_Foreach.scala 146:268:@8284.4]
  wire  x765_b504_D2; // @[package.scala 96:25:@8232.4 package.scala 96:25:@8233.4]
  wire  _T_928; // @[package.scala 96:25:@8302.4 package.scala 96:25:@8303.4]
  wire  _T_930; // @[implicits.scala 56:10:@8304.4]
  wire  _T_931; // @[sm_x536_inr_Foreach.scala 151:118:@8305.4]
  wire  _T_933; // @[sm_x536_inr_Foreach.scala 151:215:@8307.4]
  wire  _T_935; // @[sm_x536_inr_Foreach.scala 151:260:@8309.4]
  wire  _T_936; // @[sm_x536_inr_Foreach.scala 151:268:@8310.4]
  wire  _T_948; // @[package.scala 96:25:@8328.4 package.scala 96:25:@8329.4]
  wire  _T_950; // @[implicits.scala 56:10:@8330.4]
  wire  _T_951; // @[sm_x536_inr_Foreach.scala 156:118:@8331.4]
  wire  _T_953; // @[sm_x536_inr_Foreach.scala 156:215:@8333.4]
  wire  _T_955; // @[sm_x536_inr_Foreach.scala 156:260:@8335.4]
  wire  _T_956; // @[sm_x536_inr_Foreach.scala 156:268:@8336.4]
  wire [31:0] x532_sum_number; // @[Math.scala 154:22:@8222.4 Math.scala 155:14:@8223.4]
  InstrumentationCounter cycles_x536_inr_Foreach ( // @[sm_x536_inr_Foreach.scala 89:43:@8090.4]
    .clock(cycles_x536_inr_Foreach_clock),
    .reset(cycles_x536_inr_Foreach_reset),
    .io_enable(cycles_x536_inr_Foreach_io_enable),
    .io_count(cycles_x536_inr_Foreach_io_count)
  );
  InstrumentationCounter iters_x536_inr_Foreach ( // @[sm_x536_inr_Foreach.scala 90:42:@8093.4]
    .clock(iters_x536_inr_Foreach_clock),
    .reset(iters_x536_inr_Foreach_reset),
    .io_enable(iters_x536_inr_Foreach_io_enable),
    .io_count(iters_x536_inr_Foreach_io_count)
  );
  InstrumentationCounter stalls_x536_inr_Foreach ( // @[sm_x536_inr_Foreach.scala 93:43:@8102.4]
    .clock(stalls_x536_inr_Foreach_clock),
    .reset(stalls_x536_inr_Foreach_reset),
    .io_enable(stalls_x536_inr_Foreach_io_enable),
    .io_count(stalls_x536_inr_Foreach_io_count)
  );
  InstrumentationCounter idles_x536_inr_Foreach ( // @[sm_x536_inr_Foreach.scala 94:42:@8105.4]
    .clock(idles_x536_inr_Foreach_clock),
    .reset(idles_x536_inr_Foreach_reset),
    .io_enable(idles_x536_inr_Foreach_io_enable),
    .io_count(idles_x536_inr_Foreach_io_count)
  );
  _ _ ( // @[Math.scala 720:24:@8123.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x485_sub x527_sub_1 ( // @[Math.scala 191:24:@8174.4]
    .clock(x527_sub_1_clock),
    .reset(x527_sub_1_reset),
    .io_a(x527_sub_1_io_a),
    .io_b(x527_sub_1_io_b),
    .io_flow(x527_sub_1_io_flow),
    .io_result(x527_sub_1_io_result)
  );
  RetimeWrapper_32 RetimeWrapper ( // @[package.scala 93:22:@8190.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x739_sum x743_sum_1 ( // @[Math.scala 150:24:@8206.4]
    .clock(x743_sum_1_clock),
    .reset(x743_sum_1_reset),
    .io_a(x743_sum_1_io_a),
    .io_b(x743_sum_1_io_b),
    .io_flow(x743_sum_1_io_flow),
    .io_result(x743_sum_1_io_result)
  );
  x739_sum x532_sum_1 ( // @[Math.scala 150:24:@8216.4]
    .clock(x532_sum_1_clock),
    .reset(x532_sum_1_reset),
    .io_a(x532_sum_1_io_a),
    .io_b(x532_sum_1_io_b),
    .io_flow(x532_sum_1_io_flow),
    .io_result(x532_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@8227.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_2 ( // @[package.scala 93:22:@8237.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@8247.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@8257.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@8271.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@8297.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@8323.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign _T_782 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@8097.4]
  assign _T_792 = ~ io_in_x476_valid; // @[sm_x536_inr_Foreach.scala 96:62:@8112.4]
  assign b521 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x536_inr_Foreach.scala 99:18:@8131.4]
  assign _T_806 = ~ io_sigsIn_break; // @[sm_x536_inr_Foreach.scala 104:119:@8135.4]
  assign _T_818 = $signed(io_in_x505_reg_rPort_0_output_0); // @[Math.scala 493:37:@8147.4]
  assign b520_number = __io_result; // @[Math.scala 723:22:@8128.4 Math.scala 724:14:@8129.4]
  assign _T_819 = $signed(b520_number); // @[Math.scala 493:51:@8148.4]
  assign x523 = $signed(_T_818) <= $signed(_T_819); // @[Math.scala 493:44:@8149.4]
  assign _T_839 = $signed(io_in_x506_reg_rPort_0_output_0); // @[Math.scala 476:50:@8167.4]
  assign x525 = $signed(_T_819) < $signed(_T_839); // @[Math.scala 476:44:@8168.4]
  assign _T_853 = b521 & io_in_b504; // @[sm_x536_inr_Foreach.scala 121:26:@8184.4]
  assign _GEN_0 = {{1'd0}, io_in_b503_number}; // @[Math.scala 461:32:@8202.4]
  assign _T_869 = _GEN_0 << 1; // @[Math.scala 461:32:@8202.4]
  assign _T_908 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@8276.4 package.scala 96:25:@8277.4]
  assign _T_910 = io_rr ? _T_908 : 1'h0; // @[implicits.scala 56:10:@8278.4]
  assign _T_911 = _T_806 & _T_910; // @[sm_x536_inr_Foreach.scala 146:118:@8279.4]
  assign _T_913 = _T_911 & _T_806; // @[sm_x536_inr_Foreach.scala 146:215:@8281.4]
  assign x767_x526_D2 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@8252.4 package.scala 96:25:@8253.4]
  assign _T_915 = _T_913 & x767_x526_D2; // @[sm_x536_inr_Foreach.scala 146:260:@8283.4]
  assign x768_b521_D2 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@8262.4 package.scala 96:25:@8263.4]
  assign _T_916 = _T_915 & x768_b521_D2; // @[sm_x536_inr_Foreach.scala 146:268:@8284.4]
  assign x765_b504_D2 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@8232.4 package.scala 96:25:@8233.4]
  assign _T_928 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@8302.4 package.scala 96:25:@8303.4]
  assign _T_930 = io_rr ? _T_928 : 1'h0; // @[implicits.scala 56:10:@8304.4]
  assign _T_931 = _T_806 & _T_930; // @[sm_x536_inr_Foreach.scala 151:118:@8305.4]
  assign _T_933 = _T_931 & _T_806; // @[sm_x536_inr_Foreach.scala 151:215:@8307.4]
  assign _T_935 = _T_933 & x767_x526_D2; // @[sm_x536_inr_Foreach.scala 151:260:@8309.4]
  assign _T_936 = _T_935 & x768_b521_D2; // @[sm_x536_inr_Foreach.scala 151:268:@8310.4]
  assign _T_948 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@8328.4 package.scala 96:25:@8329.4]
  assign _T_950 = io_rr ? _T_948 : 1'h0; // @[implicits.scala 56:10:@8330.4]
  assign _T_951 = _T_806 & _T_950; // @[sm_x536_inr_Foreach.scala 156:118:@8331.4]
  assign _T_953 = _T_951 & _T_806; // @[sm_x536_inr_Foreach.scala 156:215:@8333.4]
  assign _T_955 = _T_953 & x767_x526_D2; // @[sm_x536_inr_Foreach.scala 156:260:@8335.4]
  assign _T_956 = _T_955 & x768_b521_D2; // @[sm_x536_inr_Foreach.scala 156:268:@8336.4]
  assign x532_sum_number = x532_sum_1_io_result; // @[Math.scala 154:22:@8222.4 Math.scala 155:14:@8223.4]
  assign io_in_x472_A_sram_1_wPort_0_ofs_0 = x532_sum_number[8:0]; // @[MemInterfaceType.scala 89:54:@8287.4]
  assign io_in_x472_A_sram_1_wPort_0_data_0 = RetimeWrapper_2_io_out; // @[MemInterfaceType.scala 90:56:@8288.4]
  assign io_in_x472_A_sram_1_wPort_0_en_0 = _T_916 & x765_b504_D2; // @[MemInterfaceType.scala 93:57:@8290.4]
  assign io_in_x471_A_sram_0_wPort_0_ofs_0 = x532_sum_number[8:0]; // @[MemInterfaceType.scala 89:54:@8313.4]
  assign io_in_x471_A_sram_0_wPort_0_data_0 = RetimeWrapper_2_io_out; // @[MemInterfaceType.scala 90:56:@8314.4]
  assign io_in_x471_A_sram_0_wPort_0_en_0 = _T_936 & x765_b504_D2; // @[MemInterfaceType.scala 93:57:@8316.4]
  assign io_in_x476_ready = _T_853 & io_sigsIn_datapathEn; // @[sm_x536_inr_Foreach.scala 121:18:@8186.4]
  assign io_in_x473_A_sram_2_wPort_0_ofs_0 = x532_sum_number[8:0]; // @[MemInterfaceType.scala 89:54:@8339.4]
  assign io_in_x473_A_sram_2_wPort_0_data_0 = RetimeWrapper_2_io_out; // @[MemInterfaceType.scala 90:56:@8340.4]
  assign io_in_x473_A_sram_2_wPort_0_en_0 = _T_956 & x765_b504_D2; // @[MemInterfaceType.scala 93:57:@8342.4]
  assign io_in_instrctrs_5_cycs = cycles_x536_inr_Foreach_io_count; // @[Ledger.scala 293:21:@8115.4]
  assign io_in_instrctrs_5_iters = iters_x536_inr_Foreach_io_count; // @[Ledger.scala 294:22:@8116.4]
  assign io_in_instrctrs_5_stalls = stalls_x536_inr_Foreach_io_count; // @[Ledger.scala 295:23:@8117.4]
  assign io_in_instrctrs_5_idles = idles_x536_inr_Foreach_io_count; // @[Ledger.scala 296:22:@8118.4]
  assign cycles_x536_inr_Foreach_clock = clock; // @[:@8091.4]
  assign cycles_x536_inr_Foreach_reset = reset; // @[:@8092.4]
  assign cycles_x536_inr_Foreach_io_enable = io_sigsIn_baseEn; // @[sm_x536_inr_Foreach.scala 91:41:@8096.4]
  assign iters_x536_inr_Foreach_clock = clock; // @[:@8094.4]
  assign iters_x536_inr_Foreach_reset = reset; // @[:@8095.4]
  assign iters_x536_inr_Foreach_io_enable = io_sigsIn_done & _T_785; // @[sm_x536_inr_Foreach.scala 92:40:@8101.4]
  assign stalls_x536_inr_Foreach_clock = clock; // @[:@8103.4]
  assign stalls_x536_inr_Foreach_reset = reset; // @[:@8104.4]
  assign stalls_x536_inr_Foreach_io_enable = 1'h0; // @[sm_x536_inr_Foreach.scala 95:41:@8110.4]
  assign idles_x536_inr_Foreach_clock = clock; // @[:@8106.4]
  assign idles_x536_inr_Foreach_reset = reset; // @[:@8107.4]
  assign idles_x536_inr_Foreach_io_enable = io_sigsIn_baseEn & _T_792; // @[sm_x536_inr_Foreach.scala 96:40:@8114.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@8126.4]
  assign x527_sub_1_clock = clock; // @[:@8175.4]
  assign x527_sub_1_reset = reset; // @[:@8176.4]
  assign x527_sub_1_io_a = __io_result; // @[Math.scala 192:17:@8177.4]
  assign x527_sub_1_io_b = io_in_x505_reg_rPort_0_output_0; // @[Math.scala 193:17:@8178.4]
  assign x527_sub_1_io_flow = 1'h1; // @[Math.scala 194:20:@8179.4]
  assign RetimeWrapper_clock = clock; // @[:@8191.4]
  assign RetimeWrapper_reset = reset; // @[:@8192.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@8194.4]
  assign RetimeWrapper_io_in = io_in_x476_bits_rdata_0; // @[package.scala 94:16:@8193.4]
  assign x743_sum_1_clock = clock; // @[:@8207.4]
  assign x743_sum_1_reset = reset; // @[:@8208.4]
  assign x743_sum_1_io_a = _T_869[31:0]; // @[Math.scala 151:17:@8209.4]
  assign x743_sum_1_io_b = io_in_b503_number; // @[Math.scala 152:17:@8210.4]
  assign x743_sum_1_io_flow = 1'h1; // @[Math.scala 153:20:@8211.4]
  assign x532_sum_1_clock = clock; // @[:@8217.4]
  assign x532_sum_1_reset = reset; // @[:@8218.4]
  assign x532_sum_1_io_a = x743_sum_1_io_result; // @[Math.scala 151:17:@8219.4]
  assign x532_sum_1_io_b = x527_sub_1_io_result; // @[Math.scala 152:17:@8220.4]
  assign x532_sum_1_io_flow = 1'h1; // @[Math.scala 153:20:@8221.4]
  assign RetimeWrapper_1_clock = clock; // @[:@8228.4]
  assign RetimeWrapper_1_reset = reset; // @[:@8229.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@8231.4]
  assign RetimeWrapper_1_io_in = io_in_b504; // @[package.scala 94:16:@8230.4]
  assign RetimeWrapper_2_clock = clock; // @[:@8238.4]
  assign RetimeWrapper_2_reset = reset; // @[:@8239.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@8241.4]
  assign RetimeWrapper_2_io_in = RetimeWrapper_io_out; // @[package.scala 94:16:@8240.4]
  assign RetimeWrapper_3_clock = clock; // @[:@8248.4]
  assign RetimeWrapper_3_reset = reset; // @[:@8249.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@8251.4]
  assign RetimeWrapper_3_io_in = x523 & x525; // @[package.scala 94:16:@8250.4]
  assign RetimeWrapper_4_clock = clock; // @[:@8258.4]
  assign RetimeWrapper_4_reset = reset; // @[:@8259.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@8261.4]
  assign RetimeWrapper_4_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@8260.4]
  assign RetimeWrapper_5_clock = clock; // @[:@8272.4]
  assign RetimeWrapper_5_reset = reset; // @[:@8273.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@8275.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@8274.4]
  assign RetimeWrapper_6_clock = clock; // @[:@8298.4]
  assign RetimeWrapper_6_reset = reset; // @[:@8299.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@8301.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@8300.4]
  assign RetimeWrapper_7_clock = clock; // @[:@8324.4]
  assign RetimeWrapper_7_reset = reset; // @[:@8325.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@8327.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@8326.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_785 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_785 <= 1'h0;
    end else begin
      _T_785 <= _T_782;
    end
  end
endmodule
module x537_outr_Foreach_kernelx537_outr_Foreach_concrete1( // @[:@8344.2]
  input         clock, // @[:@8345.4]
  input         reset, // @[:@8346.4]
  output [8:0]  io_in_x472_A_sram_1_wPort_0_ofs_0, // @[:@8347.4]
  output [31:0] io_in_x472_A_sram_1_wPort_0_data_0, // @[:@8347.4]
  output        io_in_x472_A_sram_1_wPort_0_en_0, // @[:@8347.4]
  output        io_in_x475_fifo_rPort_0_en_0, // @[:@8347.4]
  input  [95:0] io_in_x475_fifo_rPort_0_output_0, // @[:@8347.4]
  input         io_in_x475_fifo_empty, // @[:@8347.4]
  output [8:0]  io_in_x471_A_sram_0_wPort_0_ofs_0, // @[:@8347.4]
  output [31:0] io_in_x471_A_sram_0_wPort_0_data_0, // @[:@8347.4]
  output        io_in_x471_A_sram_0_wPort_0_en_0, // @[:@8347.4]
  output        io_in_x476_ready, // @[:@8347.4]
  input         io_in_x476_valid, // @[:@8347.4]
  input  [31:0] io_in_x476_bits_rdata_0, // @[:@8347.4]
  output [8:0]  io_in_x473_A_sram_2_wPort_0_ofs_0, // @[:@8347.4]
  output [31:0] io_in_x473_A_sram_2_wPort_0_data_0, // @[:@8347.4]
  output        io_in_x473_A_sram_2_wPort_0_en_0, // @[:@8347.4]
  output [63:0] io_in_instrctrs_3_cycs, // @[:@8347.4]
  output [63:0] io_in_instrctrs_3_iters, // @[:@8347.4]
  output [63:0] io_in_instrctrs_4_cycs, // @[:@8347.4]
  output [63:0] io_in_instrctrs_4_iters, // @[:@8347.4]
  output [63:0] io_in_instrctrs_4_stalls, // @[:@8347.4]
  output [63:0] io_in_instrctrs_4_idles, // @[:@8347.4]
  output [63:0] io_in_instrctrs_5_cycs, // @[:@8347.4]
  output [63:0] io_in_instrctrs_5_iters, // @[:@8347.4]
  output [63:0] io_in_instrctrs_5_stalls, // @[:@8347.4]
  output [63:0] io_in_instrctrs_5_idles, // @[:@8347.4]
  input         io_sigsIn_done, // @[:@8347.4]
  input         io_sigsIn_baseEn, // @[:@8347.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@8347.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@8347.4]
  input         io_sigsIn_smChildAcks_0, // @[:@8347.4]
  input         io_sigsIn_smChildAcks_1, // @[:@8347.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@8347.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@8347.4]
  output        io_sigsOut_smDoneIn_0, // @[:@8347.4]
  output        io_sigsOut_smDoneIn_1, // @[:@8347.4]
  output        io_sigsOut_smMaskIn_0, // @[:@8347.4]
  output        io_sigsOut_smMaskIn_1, // @[:@8347.4]
  input         io_rr // @[:@8347.4]
);
  wire  cycles_x537_outr_Foreach_clock; // @[sm_x537_outr_Foreach.scala 76:44:@8516.4]
  wire  cycles_x537_outr_Foreach_reset; // @[sm_x537_outr_Foreach.scala 76:44:@8516.4]
  wire  cycles_x537_outr_Foreach_io_enable; // @[sm_x537_outr_Foreach.scala 76:44:@8516.4]
  wire [63:0] cycles_x537_outr_Foreach_io_count; // @[sm_x537_outr_Foreach.scala 76:44:@8516.4]
  wire  iters_x537_outr_Foreach_clock; // @[sm_x537_outr_Foreach.scala 77:43:@8519.4]
  wire  iters_x537_outr_Foreach_reset; // @[sm_x537_outr_Foreach.scala 77:43:@8519.4]
  wire  iters_x537_outr_Foreach_io_enable; // @[sm_x537_outr_Foreach.scala 77:43:@8519.4]
  wire [63:0] iters_x537_outr_Foreach_io_count; // @[sm_x537_outr_Foreach.scala 77:43:@8519.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@8536.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@8536.4]
  wire  x505_reg_clock; // @[m_x505_reg.scala 27:22:@8545.4]
  wire  x505_reg_reset; // @[m_x505_reg.scala 27:22:@8545.4]
  wire [31:0] x505_reg_io_rPort_0_output_0; // @[m_x505_reg.scala 27:22:@8545.4]
  wire [31:0] x505_reg_io_wPort_0_data_0; // @[m_x505_reg.scala 27:22:@8545.4]
  wire  x505_reg_io_wPort_0_reset; // @[m_x505_reg.scala 27:22:@8545.4]
  wire  x505_reg_io_wPort_0_en_0; // @[m_x505_reg.scala 27:22:@8545.4]
  wire  x506_reg_clock; // @[m_x506_reg.scala 27:22:@8562.4]
  wire  x506_reg_reset; // @[m_x506_reg.scala 27:22:@8562.4]
  wire [31:0] x506_reg_io_rPort_0_output_0; // @[m_x506_reg.scala 27:22:@8562.4]
  wire [31:0] x506_reg_io_wPort_0_data_0; // @[m_x506_reg.scala 27:22:@8562.4]
  wire  x506_reg_io_wPort_0_reset; // @[m_x506_reg.scala 27:22:@8562.4]
  wire  x506_reg_io_wPort_0_en_0; // @[m_x506_reg.scala 27:22:@8562.4]
  wire  x507_reg_clock; // @[m_x507_reg.scala 27:22:@8579.4]
  wire  x507_reg_reset; // @[m_x507_reg.scala 27:22:@8579.4]
  wire [31:0] x507_reg_io_rPort_0_output_0; // @[m_x507_reg.scala 27:22:@8579.4]
  wire [31:0] x507_reg_io_wPort_0_data_0; // @[m_x507_reg.scala 27:22:@8579.4]
  wire  x507_reg_io_wPort_0_reset; // @[m_x507_reg.scala 27:22:@8579.4]
  wire  x507_reg_io_wPort_0_en_0; // @[m_x507_reg.scala 27:22:@8579.4]
  wire  x516_inr_UnitPipe_sm_clock; // @[sm_x516_inr_UnitPipe.scala 34:18:@8632.4]
  wire  x516_inr_UnitPipe_sm_reset; // @[sm_x516_inr_UnitPipe.scala 34:18:@8632.4]
  wire  x516_inr_UnitPipe_sm_io_enable; // @[sm_x516_inr_UnitPipe.scala 34:18:@8632.4]
  wire  x516_inr_UnitPipe_sm_io_done; // @[sm_x516_inr_UnitPipe.scala 34:18:@8632.4]
  wire  x516_inr_UnitPipe_sm_io_doneLatch; // @[sm_x516_inr_UnitPipe.scala 34:18:@8632.4]
  wire  x516_inr_UnitPipe_sm_io_ctrDone; // @[sm_x516_inr_UnitPipe.scala 34:18:@8632.4]
  wire  x516_inr_UnitPipe_sm_io_datapathEn; // @[sm_x516_inr_UnitPipe.scala 34:18:@8632.4]
  wire  x516_inr_UnitPipe_sm_io_ctrInc; // @[sm_x516_inr_UnitPipe.scala 34:18:@8632.4]
  wire  x516_inr_UnitPipe_sm_io_parentAck; // @[sm_x516_inr_UnitPipe.scala 34:18:@8632.4]
  wire  x516_inr_UnitPipe_sm_io_backpressure; // @[sm_x516_inr_UnitPipe.scala 34:18:@8632.4]
  wire  x516_inr_UnitPipe_sm_io_break; // @[sm_x516_inr_UnitPipe.scala 34:18:@8632.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@8694.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@8694.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@8694.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@8694.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@8694.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@8702.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@8702.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@8702.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@8702.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@8702.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_clock; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_reset; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x475_fifo_rPort_0_en_0; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire [95:0] x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x475_fifo_rPort_0_output_0; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x475_fifo_empty; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire [31:0] x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_data_0; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_reset; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_en_0; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_reset; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire [31:0] x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_data_0; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_reset; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_en_0; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_reset; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire [31:0] x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_data_0; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_reset; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_en_0; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_reset; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire [63:0] x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_instrctrs_4_cycs; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire [63:0] x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_instrctrs_4_iters; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire [63:0] x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_instrctrs_4_stalls; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire [63:0] x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_instrctrs_4_idles; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_done; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_forwardpressure; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_baseEn; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_break; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_rr; // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
  wire  x519_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@9000.4]
  wire  x519_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@9000.4]
  wire [31:0] x519_ctrchain_io_setup_stops_0; // @[SpatialBlocks.scala 37:22:@9000.4]
  wire  x519_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@9000.4]
  wire  x519_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@9000.4]
  wire [31:0] x519_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@9000.4]
  wire  x519_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@9000.4]
  wire  x519_ctrchain_io_output_noop; // @[SpatialBlocks.scala 37:22:@9000.4]
  wire  x519_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@9000.4]
  wire  x536_inr_Foreach_sm_clock; // @[sm_x536_inr_Foreach.scala 35:18:@9055.4]
  wire  x536_inr_Foreach_sm_reset; // @[sm_x536_inr_Foreach.scala 35:18:@9055.4]
  wire  x536_inr_Foreach_sm_io_enable; // @[sm_x536_inr_Foreach.scala 35:18:@9055.4]
  wire  x536_inr_Foreach_sm_io_done; // @[sm_x536_inr_Foreach.scala 35:18:@9055.4]
  wire  x536_inr_Foreach_sm_io_doneLatch; // @[sm_x536_inr_Foreach.scala 35:18:@9055.4]
  wire  x536_inr_Foreach_sm_io_ctrDone; // @[sm_x536_inr_Foreach.scala 35:18:@9055.4]
  wire  x536_inr_Foreach_sm_io_datapathEn; // @[sm_x536_inr_Foreach.scala 35:18:@9055.4]
  wire  x536_inr_Foreach_sm_io_ctrInc; // @[sm_x536_inr_Foreach.scala 35:18:@9055.4]
  wire  x536_inr_Foreach_sm_io_ctrRst; // @[sm_x536_inr_Foreach.scala 35:18:@9055.4]
  wire  x536_inr_Foreach_sm_io_parentAck; // @[sm_x536_inr_Foreach.scala 35:18:@9055.4]
  wire  x536_inr_Foreach_sm_io_backpressure; // @[sm_x536_inr_Foreach.scala 35:18:@9055.4]
  wire  x536_inr_Foreach_sm_io_break; // @[sm_x536_inr_Foreach.scala 35:18:@9055.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@9084.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@9084.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@9084.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@9084.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@9084.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@9124.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@9124.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@9124.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@9124.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@9124.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@9132.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@9132.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@9132.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@9132.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@9132.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_clock; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_reset; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire [8:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire [31:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_data_0; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_en_0; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_b504; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire [8:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire [31:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_data_0; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_en_0; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x476_ready; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x476_valid; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire [31:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x476_bits_rdata_0; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire [31:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_b503_number; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire [31:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x505_reg_rPort_0_output_0; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire [8:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire [31:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_data_0; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_en_0; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire [31:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x506_reg_rPort_0_output_0; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire [63:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_instrctrs_5_cycs; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire [63:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_instrctrs_5_iters; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire [63:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_instrctrs_5_stalls; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire [63:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_instrctrs_5_idles; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_done; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire [31:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_rr; // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
  wire  _T_712; // @[package.scala 100:49:@8523.4]
  reg  _T_715; // @[package.scala 48:56:@8524.4]
  reg [31:0] _RAND_0;
  wire  b504; // @[sm_x537_outr_Foreach.scala 82:18:@8544.4]
  wire  _T_787; // @[package.scala 100:49:@8660.4]
  reg  _T_790; // @[package.scala 48:56:@8661.4]
  reg [31:0] _RAND_1;
  wire  _T_798; // @[sm_x537_outr_Foreach.scala 89:46:@8668.4]
  wire  x516_inr_UnitPipe_mySignalsIn_forwardpressure; // @[sm_x537_outr_Foreach.scala 89:115:@8672.4]
  wire  _T_811; // @[package.scala 96:25:@8699.4 package.scala 96:25:@8700.4]
  wire  _T_817; // @[package.scala 96:25:@8707.4 package.scala 96:25:@8708.4]
  wire  _T_820; // @[SpatialBlocks.scala 137:99:@8710.4]
  wire  x516_inr_UnitPipe_mySignalsIn_baseEn; // @[SpatialBlocks.scala 137:96:@8711.4]
  wire [31:0] x734_rd_x507_number; // @[sm_x537_outr_Foreach.scala 95:30:@8986.4 sm_x537_outr_Foreach.scala 100:202:@8999.4]
  wire  _T_908; // @[package.scala 96:25:@9089.4 package.scala 96:25:@9090.4]
  wire  x536_inr_Foreach_mySignalsIn_forwardpressure; // @[sm_x537_outr_Foreach.scala 108:68:@9096.4]
  wire  _T_917; // @[sm_x537_outr_Foreach.scala 111:32:@9100.4]
  wire  x536_inr_Foreach_mySignalsIn_mask; // @[sm_x537_outr_Foreach.scala 111:74:@9101.4]
  wire  _T_923; // @[package.scala 96:25:@9129.4 package.scala 96:25:@9130.4]
  wire  _T_929; // @[package.scala 96:25:@9137.4 package.scala 96:25:@9138.4]
  wire  _T_932; // @[SpatialBlocks.scala 137:99:@9140.4]
  wire  x536_inr_Foreach_mySignalsIn_baseEn; // @[SpatialBlocks.scala 137:96:@9141.4]
  wire  _T_934; // @[SpatialBlocks.scala 156:36:@9149.4]
  wire  _T_935; // @[SpatialBlocks.scala 156:78:@9150.4]
  wire  _T_942; // @[SpatialBlocks.scala 158:58:@9162.4]
  InstrumentationCounter cycles_x537_outr_Foreach ( // @[sm_x537_outr_Foreach.scala 76:44:@8516.4]
    .clock(cycles_x537_outr_Foreach_clock),
    .reset(cycles_x537_outr_Foreach_reset),
    .io_enable(cycles_x537_outr_Foreach_io_enable),
    .io_count(cycles_x537_outr_Foreach_io_count)
  );
  InstrumentationCounter iters_x537_outr_Foreach ( // @[sm_x537_outr_Foreach.scala 77:43:@8519.4]
    .clock(iters_x537_outr_Foreach_clock),
    .reset(iters_x537_outr_Foreach_reset),
    .io_enable(iters_x537_outr_Foreach_io_enable),
    .io_count(iters_x537_outr_Foreach_io_count)
  );
  _ _ ( // @[Math.scala 720:24:@8536.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x505_reg x505_reg ( // @[m_x505_reg.scala 27:22:@8545.4]
    .clock(x505_reg_clock),
    .reset(x505_reg_reset),
    .io_rPort_0_output_0(x505_reg_io_rPort_0_output_0),
    .io_wPort_0_data_0(x505_reg_io_wPort_0_data_0),
    .io_wPort_0_reset(x505_reg_io_wPort_0_reset),
    .io_wPort_0_en_0(x505_reg_io_wPort_0_en_0)
  );
  x505_reg x506_reg ( // @[m_x506_reg.scala 27:22:@8562.4]
    .clock(x506_reg_clock),
    .reset(x506_reg_reset),
    .io_rPort_0_output_0(x506_reg_io_rPort_0_output_0),
    .io_wPort_0_data_0(x506_reg_io_wPort_0_data_0),
    .io_wPort_0_reset(x506_reg_io_wPort_0_reset),
    .io_wPort_0_en_0(x506_reg_io_wPort_0_en_0)
  );
  x505_reg x507_reg ( // @[m_x507_reg.scala 27:22:@8579.4]
    .clock(x507_reg_clock),
    .reset(x507_reg_reset),
    .io_rPort_0_output_0(x507_reg_io_rPort_0_output_0),
    .io_wPort_0_data_0(x507_reg_io_wPort_0_data_0),
    .io_wPort_0_reset(x507_reg_io_wPort_0_reset),
    .io_wPort_0_en_0(x507_reg_io_wPort_0_en_0)
  );
  x516_inr_UnitPipe_sm x516_inr_UnitPipe_sm ( // @[sm_x516_inr_UnitPipe.scala 34:18:@8632.4]
    .clock(x516_inr_UnitPipe_sm_clock),
    .reset(x516_inr_UnitPipe_sm_reset),
    .io_enable(x516_inr_UnitPipe_sm_io_enable),
    .io_done(x516_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x516_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x516_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x516_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x516_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x516_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x516_inr_UnitPipe_sm_io_backpressure),
    .io_break(x516_inr_UnitPipe_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@8694.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@8702.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1 x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1 ( // @[sm_x516_inr_UnitPipe.scala 117:24:@8731.4]
    .clock(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_clock),
    .reset(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_reset),
    .io_in_x475_fifo_rPort_0_en_0(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x475_fifo_rPort_0_en_0),
    .io_in_x475_fifo_rPort_0_output_0(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x475_fifo_rPort_0_output_0),
    .io_in_x475_fifo_empty(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x475_fifo_empty),
    .io_in_x507_reg_wPort_0_data_0(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_data_0),
    .io_in_x507_reg_wPort_0_reset(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_reset),
    .io_in_x507_reg_wPort_0_en_0(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_en_0),
    .io_in_x507_reg_reset(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_reset),
    .io_in_x505_reg_wPort_0_data_0(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_data_0),
    .io_in_x505_reg_wPort_0_reset(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_reset),
    .io_in_x505_reg_wPort_0_en_0(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_en_0),
    .io_in_x505_reg_reset(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_reset),
    .io_in_x506_reg_wPort_0_data_0(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_data_0),
    .io_in_x506_reg_wPort_0_reset(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_reset),
    .io_in_x506_reg_wPort_0_en_0(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_en_0),
    .io_in_x506_reg_reset(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_reset),
    .io_in_instrctrs_4_cycs(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_instrctrs_4_cycs),
    .io_in_instrctrs_4_iters(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_instrctrs_4_iters),
    .io_in_instrctrs_4_stalls(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_instrctrs_4_stalls),
    .io_in_instrctrs_4_idles(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_instrctrs_4_idles),
    .io_sigsIn_done(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_done),
    .io_sigsIn_forwardpressure(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_forwardpressure),
    .io_sigsIn_datapathEn(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_break),
    .io_rr(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_rr)
  );
  x519_ctrchain x519_ctrchain ( // @[SpatialBlocks.scala 37:22:@9000.4]
    .clock(x519_ctrchain_clock),
    .reset(x519_ctrchain_reset),
    .io_setup_stops_0(x519_ctrchain_io_setup_stops_0),
    .io_input_reset(x519_ctrchain_io_input_reset),
    .io_input_enable(x519_ctrchain_io_input_enable),
    .io_output_counts_0(x519_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x519_ctrchain_io_output_oobs_0),
    .io_output_noop(x519_ctrchain_io_output_noop),
    .io_output_done(x519_ctrchain_io_output_done)
  );
  x536_inr_Foreach_sm x536_inr_Foreach_sm ( // @[sm_x536_inr_Foreach.scala 35:18:@9055.4]
    .clock(x536_inr_Foreach_sm_clock),
    .reset(x536_inr_Foreach_sm_reset),
    .io_enable(x536_inr_Foreach_sm_io_enable),
    .io_done(x536_inr_Foreach_sm_io_done),
    .io_doneLatch(x536_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x536_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x536_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x536_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x536_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x536_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x536_inr_Foreach_sm_io_backpressure),
    .io_break(x536_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@9084.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@9124.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@9132.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1 x536_inr_Foreach_kernelx536_inr_Foreach_concrete1 ( // @[sm_x536_inr_Foreach.scala 158:24:@9166.4]
    .clock(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_clock),
    .reset(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_reset),
    .io_in_x472_A_sram_1_wPort_0_ofs_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0),
    .io_in_x472_A_sram_1_wPort_0_data_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_data_0),
    .io_in_x472_A_sram_1_wPort_0_en_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_en_0),
    .io_in_b504(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_b504),
    .io_in_x471_A_sram_0_wPort_0_ofs_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0),
    .io_in_x471_A_sram_0_wPort_0_data_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_data_0),
    .io_in_x471_A_sram_0_wPort_0_en_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_en_0),
    .io_in_x476_ready(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x476_ready),
    .io_in_x476_valid(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x476_valid),
    .io_in_x476_bits_rdata_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x476_bits_rdata_0),
    .io_in_b503_number(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_b503_number),
    .io_in_x505_reg_rPort_0_output_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x505_reg_rPort_0_output_0),
    .io_in_x473_A_sram_2_wPort_0_ofs_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0),
    .io_in_x473_A_sram_2_wPort_0_data_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_data_0),
    .io_in_x473_A_sram_2_wPort_0_en_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_en_0),
    .io_in_x506_reg_rPort_0_output_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x506_reg_rPort_0_output_0),
    .io_in_instrctrs_5_cycs(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_instrctrs_5_cycs),
    .io_in_instrctrs_5_iters(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_instrctrs_5_iters),
    .io_in_instrctrs_5_stalls(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_instrctrs_5_stalls),
    .io_in_instrctrs_5_idles(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_instrctrs_5_idles),
    .io_sigsIn_done(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_datapathEn(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_rr)
  );
  assign _T_712 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@8523.4]
  assign b504 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x537_outr_Foreach.scala 82:18:@8544.4]
  assign _T_787 = x516_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@8660.4]
  assign _T_798 = ~ io_in_x475_fifo_empty; // @[sm_x537_outr_Foreach.scala 89:46:@8668.4]
  assign x516_inr_UnitPipe_mySignalsIn_forwardpressure = _T_798 | x516_inr_UnitPipe_sm_io_doneLatch; // @[sm_x537_outr_Foreach.scala 89:115:@8672.4]
  assign _T_811 = RetimeWrapper_io_out; // @[package.scala 96:25:@8699.4 package.scala 96:25:@8700.4]
  assign _T_817 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@8707.4 package.scala 96:25:@8708.4]
  assign _T_820 = ~ _T_817; // @[SpatialBlocks.scala 137:99:@8710.4]
  assign x516_inr_UnitPipe_mySignalsIn_baseEn = _T_811 & _T_820; // @[SpatialBlocks.scala 137:96:@8711.4]
  assign x734_rd_x507_number = x507_reg_io_rPort_0_output_0; // @[sm_x537_outr_Foreach.scala 95:30:@8986.4 sm_x537_outr_Foreach.scala 100:202:@8999.4]
  assign _T_908 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@9089.4 package.scala 96:25:@9090.4]
  assign x536_inr_Foreach_mySignalsIn_forwardpressure = io_in_x476_valid | x536_inr_Foreach_sm_io_doneLatch; // @[sm_x537_outr_Foreach.scala 108:68:@9096.4]
  assign _T_917 = ~ x519_ctrchain_io_output_noop; // @[sm_x537_outr_Foreach.scala 111:32:@9100.4]
  assign x536_inr_Foreach_mySignalsIn_mask = _T_917 & b504; // @[sm_x537_outr_Foreach.scala 111:74:@9101.4]
  assign _T_923 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@9129.4 package.scala 96:25:@9130.4]
  assign _T_929 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@9137.4 package.scala 96:25:@9138.4]
  assign _T_932 = ~ _T_929; // @[SpatialBlocks.scala 137:99:@9140.4]
  assign x536_inr_Foreach_mySignalsIn_baseEn = _T_923 & _T_932; // @[SpatialBlocks.scala 137:96:@9141.4]
  assign _T_934 = x536_inr_Foreach_sm_io_datapathEn & x536_inr_Foreach_mySignalsIn_mask; // @[SpatialBlocks.scala 156:36:@9149.4]
  assign _T_935 = ~ x536_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 156:78:@9150.4]
  assign _T_942 = x536_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 158:58:@9162.4]
  assign io_in_x472_A_sram_1_wPort_0_ofs_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@9368.4]
  assign io_in_x472_A_sram_1_wPort_0_data_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@9367.4]
  assign io_in_x472_A_sram_1_wPort_0_en_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@9363.4]
  assign io_in_x475_fifo_rPort_0_en_0 = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x475_fifo_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@8931.4]
  assign io_in_x471_A_sram_0_wPort_0_ofs_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@9376.4]
  assign io_in_x471_A_sram_0_wPort_0_data_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@9375.4]
  assign io_in_x471_A_sram_0_wPort_0_en_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@9371.4]
  assign io_in_x476_ready = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x476_ready; // @[sm_x536_inr_Foreach.scala 67:23:@9380.4]
  assign io_in_x473_A_sram_2_wPort_0_ofs_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@9392.4]
  assign io_in_x473_A_sram_2_wPort_0_data_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@9391.4]
  assign io_in_x473_A_sram_2_wPort_0_en_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@9387.4]
  assign io_in_instrctrs_3_cycs = cycles_x537_outr_Foreach_io_count; // @[Ledger.scala 293:21:@8528.4]
  assign io_in_instrctrs_3_iters = iters_x537_outr_Foreach_io_count; // @[Ledger.scala 294:22:@8529.4]
  assign io_in_instrctrs_4_cycs = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_instrctrs_4_cycs; // @[Ledger.scala 302:78:@8958.4]
  assign io_in_instrctrs_4_iters = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_instrctrs_4_iters; // @[Ledger.scala 302:78:@8957.4]
  assign io_in_instrctrs_4_stalls = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_instrctrs_4_stalls; // @[Ledger.scala 302:78:@8956.4]
  assign io_in_instrctrs_4_idles = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_instrctrs_4_idles; // @[Ledger.scala 302:78:@8955.4]
  assign io_in_instrctrs_5_cycs = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_instrctrs_5_cycs; // @[Ledger.scala 302:78:@9402.4]
  assign io_in_instrctrs_5_iters = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_instrctrs_5_iters; // @[Ledger.scala 302:78:@9401.4]
  assign io_in_instrctrs_5_stalls = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_instrctrs_5_stalls; // @[Ledger.scala 302:78:@9400.4]
  assign io_in_instrctrs_5_idles = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_instrctrs_5_idles; // @[Ledger.scala 302:78:@9399.4]
  assign io_sigsOut_smDoneIn_0 = x516_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 155:56:@8717.4]
  assign io_sigsOut_smDoneIn_1 = x536_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@9147.4]
  assign io_sigsOut_smMaskIn_0 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[SpatialBlocks.scala 155:86:@8718.4]
  assign io_sigsOut_smMaskIn_1 = _T_917 & b504; // @[SpatialBlocks.scala 155:86:@9148.4]
  assign cycles_x537_outr_Foreach_clock = clock; // @[:@8517.4]
  assign cycles_x537_outr_Foreach_reset = reset; // @[:@8518.4]
  assign cycles_x537_outr_Foreach_io_enable = io_sigsIn_baseEn; // @[sm_x537_outr_Foreach.scala 78:42:@8522.4]
  assign iters_x537_outr_Foreach_clock = clock; // @[:@8520.4]
  assign iters_x537_outr_Foreach_reset = reset; // @[:@8521.4]
  assign iters_x537_outr_Foreach_io_enable = io_sigsIn_done & _T_715; // @[sm_x537_outr_Foreach.scala 79:41:@8527.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@8539.4]
  assign x505_reg_clock = clock; // @[:@8546.4]
  assign x505_reg_reset = reset; // @[:@8547.4]
  assign x505_reg_io_wPort_0_data_0 = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@8945.4]
  assign x505_reg_io_wPort_0_reset = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_reset; // @[MemInterfaceType.scala 67:44:@8944.4]
  assign x505_reg_io_wPort_0_en_0 = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@8941.4]
  assign x506_reg_clock = clock; // @[:@8563.4]
  assign x506_reg_reset = reset; // @[:@8564.4]
  assign x506_reg_io_wPort_0_data_0 = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@8952.4]
  assign x506_reg_io_wPort_0_reset = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_reset; // @[MemInterfaceType.scala 67:44:@8951.4]
  assign x506_reg_io_wPort_0_en_0 = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@8948.4]
  assign x507_reg_clock = clock; // @[:@8580.4]
  assign x507_reg_reset = reset; // @[:@8581.4]
  assign x507_reg_io_wPort_0_data_0 = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@8938.4]
  assign x507_reg_io_wPort_0_reset = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_reset; // @[MemInterfaceType.scala 67:44:@8937.4]
  assign x507_reg_io_wPort_0_en_0 = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@8934.4]
  assign x516_inr_UnitPipe_sm_clock = clock; // @[:@8633.4]
  assign x516_inr_UnitPipe_sm_reset = reset; // @[:@8634.4]
  assign x516_inr_UnitPipe_sm_io_enable = x516_inr_UnitPipe_mySignalsIn_baseEn & x516_inr_UnitPipe_mySignalsIn_forwardpressure; // @[SpatialBlocks.scala 139:18:@8714.4]
  assign x516_inr_UnitPipe_sm_io_ctrDone = x516_inr_UnitPipe_sm_io_ctrInc & _T_790; // @[sm_x537_outr_Foreach.scala 87:39:@8664.4]
  assign x516_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@8716.4]
  assign x516_inr_UnitPipe_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@8688.4]
  assign x516_inr_UnitPipe_sm_io_break = 1'h0; // @[sm_x537_outr_Foreach.scala 91:37:@8675.4]
  assign RetimeWrapper_clock = clock; // @[:@8695.4]
  assign RetimeWrapper_reset = reset; // @[:@8696.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@8698.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@8697.4]
  assign RetimeWrapper_1_clock = clock; // @[:@8703.4]
  assign RetimeWrapper_1_reset = reset; // @[:@8704.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@8706.4]
  assign RetimeWrapper_1_io_in = x516_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@8705.4]
  assign x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_clock = clock; // @[:@8732.4]
  assign x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_reset = reset; // @[:@8733.4]
  assign x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x475_fifo_rPort_0_output_0 = io_in_x475_fifo_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@8929.4]
  assign x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x475_fifo_empty = io_in_x475_fifo_empty; // @[MemInterfaceType.scala 161:16:@8925.4]
  assign x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_done = x516_inr_UnitPipe_sm_io_done; // @[sm_x516_inr_UnitPipe.scala 123:22:@8978.4]
  assign x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_forwardpressure = _T_798 | x516_inr_UnitPipe_sm_io_doneLatch; // @[sm_x516_inr_UnitPipe.scala 123:22:@8972.4]
  assign x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x516_inr_UnitPipe_sm_io_datapathEn & b504; // @[sm_x516_inr_UnitPipe.scala 123:22:@8971.4]
  assign x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_baseEn = _T_811 & _T_820; // @[sm_x516_inr_UnitPipe.scala 123:22:@8970.4]
  assign x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_break = x516_inr_UnitPipe_sm_io_break; // @[sm_x516_inr_UnitPipe.scala 123:22:@8969.4]
  assign x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x516_inr_UnitPipe.scala 122:18:@8959.4]
  assign x519_ctrchain_clock = clock; // @[:@9001.4]
  assign x519_ctrchain_reset = reset; // @[:@9002.4]
  assign x519_ctrchain_io_setup_stops_0 = $signed(x734_rd_x507_number); // @[SpatialBlocks.scala 40:87:@9016.4]
  assign x519_ctrchain_io_input_reset = x536_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@9165.4]
  assign x519_ctrchain_io_input_enable = _T_942 & x536_inr_Foreach_mySignalsIn_forwardpressure; // @[SpatialBlocks.scala 158:42:@9164.4]
  assign x536_inr_Foreach_sm_clock = clock; // @[:@9056.4]
  assign x536_inr_Foreach_sm_reset = reset; // @[:@9057.4]
  assign x536_inr_Foreach_sm_io_enable = x536_inr_Foreach_mySignalsIn_baseEn & x536_inr_Foreach_mySignalsIn_forwardpressure; // @[SpatialBlocks.scala 139:18:@9144.4]
  assign x536_inr_Foreach_sm_io_ctrDone = io_rr ? _T_908 : 1'h0; // @[sm_x537_outr_Foreach.scala 106:38:@9092.4]
  assign x536_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 141:21:@9146.4]
  assign x536_inr_Foreach_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@9118.4]
  assign x536_inr_Foreach_sm_io_break = 1'h0; // @[sm_x537_outr_Foreach.scala 110:36:@9099.4]
  assign RetimeWrapper_2_clock = clock; // @[:@9085.4]
  assign RetimeWrapper_2_reset = reset; // @[:@9086.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@9088.4]
  assign RetimeWrapper_2_io_in = x519_ctrchain_io_output_done; // @[package.scala 94:16:@9087.4]
  assign RetimeWrapper_3_clock = clock; // @[:@9125.4]
  assign RetimeWrapper_3_reset = reset; // @[:@9126.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@9128.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@9127.4]
  assign RetimeWrapper_4_clock = clock; // @[:@9133.4]
  assign RetimeWrapper_4_reset = reset; // @[:@9134.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@9136.4]
  assign RetimeWrapper_4_io_in = x536_inr_Foreach_sm_io_done; // @[package.scala 94:16:@9135.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_clock = clock; // @[:@9167.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_reset = reset; // @[:@9168.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_b504 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x536_inr_Foreach.scala 65:23:@9370.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x476_valid = io_in_x476_valid; // @[sm_x536_inr_Foreach.scala 67:23:@9379.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x476_bits_rdata_0 = io_in_x476_bits_rdata_0; // @[sm_x536_inr_Foreach.scala 67:23:@9378.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_b503_number = __io_result; // @[sm_x536_inr_Foreach.scala 68:23:@9381.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x505_reg_rPort_0_output_0 = x505_reg_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@9382.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x506_reg_rPort_0_output_0 = x506_reg_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@9394.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_done = x536_inr_Foreach_sm_io_done; // @[sm_x536_inr_Foreach.scala 164:22:@9422.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_934 & _T_935; // @[sm_x536_inr_Foreach.scala 164:22:@9415.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_baseEn = _T_923 & _T_932; // @[sm_x536_inr_Foreach.scala 164:22:@9414.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_break = x536_inr_Foreach_sm_io_break; // @[sm_x536_inr_Foreach.scala 164:22:@9413.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x519_ctrchain_io_output_counts_0; // @[sm_x536_inr_Foreach.scala 164:22:@9408.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x519_ctrchain_io_output_oobs_0; // @[sm_x536_inr_Foreach.scala 164:22:@9407.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x536_inr_Foreach.scala 163:18:@9403.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_715 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_790 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_715 <= 1'h0;
    end else begin
      _T_715 <= _T_712;
    end
    if (reset) begin
      _T_790 <= 1'h0;
    end else begin
      _T_790 <= _T_787;
    end
  end
endmodule
module x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1( // @[:@9431.2]
  input         clock, // @[:@9432.4]
  input         reset, // @[:@9433.4]
  input  [63:0] io_in_x468_A_dram_number, // @[:@9434.4]
  output [8:0]  io_in_x472_A_sram_1_wPort_0_ofs_0, // @[:@9434.4]
  output [31:0] io_in_x472_A_sram_1_wPort_0_data_0, // @[:@9434.4]
  output        io_in_x472_A_sram_1_wPort_0_en_0, // @[:@9434.4]
  output [8:0]  io_in_x471_A_sram_0_wPort_0_ofs_0, // @[:@9434.4]
  output [31:0] io_in_x471_A_sram_0_wPort_0_data_0, // @[:@9434.4]
  output        io_in_x471_A_sram_0_wPort_0_en_0, // @[:@9434.4]
  output        io_in_x476_ready, // @[:@9434.4]
  input         io_in_x476_valid, // @[:@9434.4]
  input  [31:0] io_in_x476_bits_rdata_0, // @[:@9434.4]
  output [8:0]  io_in_x473_A_sram_2_wPort_0_ofs_0, // @[:@9434.4]
  output [31:0] io_in_x473_A_sram_2_wPort_0_data_0, // @[:@9434.4]
  output        io_in_x473_A_sram_2_wPort_0_en_0, // @[:@9434.4]
  input         io_in_x474_ready, // @[:@9434.4]
  output        io_in_x474_valid, // @[:@9434.4]
  output [63:0] io_in_x474_bits_addr, // @[:@9434.4]
  output [31:0] io_in_x474_bits_size, // @[:@9434.4]
  output [63:0] io_in_instrctrs_1_cycs, // @[:@9434.4]
  output [63:0] io_in_instrctrs_1_iters, // @[:@9434.4]
  output [63:0] io_in_instrctrs_2_cycs, // @[:@9434.4]
  output [63:0] io_in_instrctrs_2_iters, // @[:@9434.4]
  output [63:0] io_in_instrctrs_2_stalls, // @[:@9434.4]
  output [63:0] io_in_instrctrs_2_idles, // @[:@9434.4]
  output [63:0] io_in_instrctrs_3_cycs, // @[:@9434.4]
  output [63:0] io_in_instrctrs_3_iters, // @[:@9434.4]
  output [63:0] io_in_instrctrs_4_cycs, // @[:@9434.4]
  output [63:0] io_in_instrctrs_4_iters, // @[:@9434.4]
  output [63:0] io_in_instrctrs_4_stalls, // @[:@9434.4]
  output [63:0] io_in_instrctrs_4_idles, // @[:@9434.4]
  output [63:0] io_in_instrctrs_5_cycs, // @[:@9434.4]
  output [63:0] io_in_instrctrs_5_iters, // @[:@9434.4]
  output [63:0] io_in_instrctrs_5_stalls, // @[:@9434.4]
  output [63:0] io_in_instrctrs_5_idles, // @[:@9434.4]
  input         io_sigsIn_done, // @[:@9434.4]
  input         io_sigsIn_baseEn, // @[:@9434.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@9434.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@9434.4]
  input         io_sigsIn_smChildAcks_0, // @[:@9434.4]
  input         io_sigsIn_smChildAcks_1, // @[:@9434.4]
  output        io_sigsOut_smDoneIn_0, // @[:@9434.4]
  output        io_sigsOut_smDoneIn_1, // @[:@9434.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@9434.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@9434.4]
  input         io_rr // @[:@9434.4]
);
  wire  cycles_x538_outr_UnitPipe_DenseTransfer_clock; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 81:59:@9583.4]
  wire  cycles_x538_outr_UnitPipe_DenseTransfer_reset; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 81:59:@9583.4]
  wire  cycles_x538_outr_UnitPipe_DenseTransfer_io_enable; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 81:59:@9583.4]
  wire [63:0] cycles_x538_outr_UnitPipe_DenseTransfer_io_count; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 81:59:@9583.4]
  wire  iters_x538_outr_UnitPipe_DenseTransfer_clock; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 82:58:@9586.4]
  wire  iters_x538_outr_UnitPipe_DenseTransfer_reset; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 82:58:@9586.4]
  wire  iters_x538_outr_UnitPipe_DenseTransfer_io_enable; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 82:58:@9586.4]
  wire [63:0] iters_x538_outr_UnitPipe_DenseTransfer_io_count; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 82:58:@9586.4]
  wire  x475_fifo_clock; // @[m_x475_fifo.scala 27:22:@9599.4]
  wire  x475_fifo_reset; // @[m_x475_fifo.scala 27:22:@9599.4]
  wire  x475_fifo_io_rPort_0_en_0; // @[m_x475_fifo.scala 27:22:@9599.4]
  wire [95:0] x475_fifo_io_rPort_0_output_0; // @[m_x475_fifo.scala 27:22:@9599.4]
  wire [95:0] x475_fifo_io_wPort_0_data_0; // @[m_x475_fifo.scala 27:22:@9599.4]
  wire  x475_fifo_io_wPort_0_en_0; // @[m_x475_fifo.scala 27:22:@9599.4]
  wire  x475_fifo_io_full; // @[m_x475_fifo.scala 27:22:@9599.4]
  wire  x475_fifo_io_empty; // @[m_x475_fifo.scala 27:22:@9599.4]
  wire  x475_fifo_io_active_0_in; // @[m_x475_fifo.scala 27:22:@9599.4]
  wire  x475_fifo_io_active_0_out; // @[m_x475_fifo.scala 27:22:@9599.4]
  wire  x478_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@9625.4]
  wire  x478_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@9625.4]
  wire  x478_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@9625.4]
  wire  x478_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@9625.4]
  wire [8:0] x478_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@9625.4]
  wire  x478_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@9625.4]
  wire  x478_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@9625.4]
  wire  x499_inr_Foreach_sm_clock; // @[sm_x499_inr_Foreach.scala 34:18:@9678.4]
  wire  x499_inr_Foreach_sm_reset; // @[sm_x499_inr_Foreach.scala 34:18:@9678.4]
  wire  x499_inr_Foreach_sm_io_enable; // @[sm_x499_inr_Foreach.scala 34:18:@9678.4]
  wire  x499_inr_Foreach_sm_io_done; // @[sm_x499_inr_Foreach.scala 34:18:@9678.4]
  wire  x499_inr_Foreach_sm_io_doneLatch; // @[sm_x499_inr_Foreach.scala 34:18:@9678.4]
  wire  x499_inr_Foreach_sm_io_rst; // @[sm_x499_inr_Foreach.scala 34:18:@9678.4]
  wire  x499_inr_Foreach_sm_io_ctrDone; // @[sm_x499_inr_Foreach.scala 34:18:@9678.4]
  wire  x499_inr_Foreach_sm_io_datapathEn; // @[sm_x499_inr_Foreach.scala 34:18:@9678.4]
  wire  x499_inr_Foreach_sm_io_ctrInc; // @[sm_x499_inr_Foreach.scala 34:18:@9678.4]
  wire  x499_inr_Foreach_sm_io_ctrRst; // @[sm_x499_inr_Foreach.scala 34:18:@9678.4]
  wire  x499_inr_Foreach_sm_io_parentAck; // @[sm_x499_inr_Foreach.scala 34:18:@9678.4]
  wire  x499_inr_Foreach_sm_io_backpressure; // @[sm_x499_inr_Foreach.scala 34:18:@9678.4]
  wire  x499_inr_Foreach_sm_io_break; // @[sm_x499_inr_Foreach.scala 34:18:@9678.4]
  wire  x499_inr_Foreach_iiCtr_clock; // @[sm_x499_inr_Foreach.scala 35:21:@9703.4]
  wire  x499_inr_Foreach_iiCtr_reset; // @[sm_x499_inr_Foreach.scala 35:21:@9703.4]
  wire  x499_inr_Foreach_iiCtr_io_input_enable; // @[sm_x499_inr_Foreach.scala 35:21:@9703.4]
  wire  x499_inr_Foreach_iiCtr_io_input_reset; // @[sm_x499_inr_Foreach.scala 35:21:@9703.4]
  wire  x499_inr_Foreach_iiCtr_io_output_issue; // @[sm_x499_inr_Foreach.scala 35:21:@9703.4]
  wire  x499_inr_Foreach_iiCtr_io_output_done; // @[sm_x499_inr_Foreach.scala 35:21:@9703.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@9707.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@9707.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@9707.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@9707.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@9707.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@9716.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@9716.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@9716.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@9716.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@9716.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@9759.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@9759.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@9759.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@9759.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@9759.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@9767.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@9767.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@9767.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@9767.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@9767.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_clock; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_reset; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire [63:0] x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x468_A_dram_number; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire [95:0] x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_wPort_0_data_0; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_wPort_0_en_0; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_full; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_active_0_in; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_active_0_out; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_ready; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_valid; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire [63:0] x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_bits_addr; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire [31:0] x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_bits_size; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire [63:0] x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_instrctrs_2_cycs; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire [63:0] x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_instrctrs_2_iters; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire [63:0] x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_instrctrs_2_stalls; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire [63:0] x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_instrctrs_2_idles; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_done; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_iiIssue; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire [31:0] x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_rr; // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
  wire  x502_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@10007.4]
  wire  x502_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@10007.4]
  wire  x502_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@10007.4]
  wire  x502_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@10007.4]
  wire [8:0] x502_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@10007.4]
  wire  x502_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@10007.4]
  wire  x502_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@10007.4]
  wire  x537_outr_Foreach_sm_clock; // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
  wire  x537_outr_Foreach_sm_reset; // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
  wire  x537_outr_Foreach_sm_io_enable; // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
  wire  x537_outr_Foreach_sm_io_done; // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
  wire  x537_outr_Foreach_sm_io_ctrDone; // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
  wire  x537_outr_Foreach_sm_io_ctrInc; // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
  wire  x537_outr_Foreach_sm_io_ctrRst; // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
  wire  x537_outr_Foreach_sm_io_parentAck; // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
  wire  x537_outr_Foreach_sm_io_doneIn_0; // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
  wire  x537_outr_Foreach_sm_io_doneIn_1; // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
  wire  x537_outr_Foreach_sm_io_maskIn_0; // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
  wire  x537_outr_Foreach_sm_io_maskIn_1; // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
  wire  x537_outr_Foreach_sm_io_enableOut_0; // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
  wire  x537_outr_Foreach_sm_io_enableOut_1; // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
  wire  x537_outr_Foreach_sm_io_childAck_0; // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
  wire  x537_outr_Foreach_sm_io_childAck_1; // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@10099.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@10099.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@10099.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@10099.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@10099.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@10144.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@10144.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@10144.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@10144.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@10144.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@10152.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@10152.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@10152.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@10152.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@10152.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_clock; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_reset; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [8:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [31:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_data_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_en_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_rPort_0_en_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [95:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_rPort_0_output_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_empty; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [8:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [31:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_data_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_en_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_ready; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_valid; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [31:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_bits_rdata_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [8:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [31:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_data_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_en_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [63:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_3_cycs; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [63:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_3_iters; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [63:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_4_cycs; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [63:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_4_iters; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [63:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_4_stalls; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [63:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_4_idles; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [63:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_5_cycs; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [63:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_5_iters; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [63:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_5_stalls; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [63:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_5_idles; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_done; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire [31:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_rr; // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
  wire  _T_546; // @[package.scala 100:49:@9590.4]
  reg  _T_549; // @[package.scala 48:56:@9591.4]
  reg [31:0] _RAND_0;
  wire  _T_616; // @[package.scala 96:25:@9712.4 package.scala 96:25:@9713.4]
  wire  _T_622; // @[package.scala 96:25:@9721.4 package.scala 96:25:@9722.4]
  wire  _T_625; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 93:41:@9724.4]
  wire  _T_626; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 93:68:@9725.4]
  wire  _T_627; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 93:66:@9726.4]
  wire  _T_628; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 93:96:@9727.4]
  wire  _T_642; // @[package.scala 96:25:@9764.4 package.scala 96:25:@9765.4]
  wire  _T_648; // @[package.scala 96:25:@9772.4 package.scala 96:25:@9773.4]
  wire  _T_651; // @[SpatialBlocks.scala 137:99:@9775.4]
  wire  _T_653; // @[SpatialBlocks.scala 156:36:@9784.4]
  wire  _T_654; // @[SpatialBlocks.scala 156:78:@9785.4]
  wire  x499_inr_Foreach_mySignalsIn_iiDone; // @[SpatialBlocks.scala 157:126:@9792.4]
  wire  _T_725; // @[package.scala 96:25:@10104.4 package.scala 96:25:@10105.4]
  wire  _T_742; // @[package.scala 96:25:@10149.4 package.scala 96:25:@10150.4]
  wire  _T_748; // @[package.scala 96:25:@10157.4 package.scala 96:25:@10158.4]
  wire  _T_751; // @[SpatialBlocks.scala 137:99:@10160.4]
  InstrumentationCounter cycles_x538_outr_UnitPipe_DenseTransfer ( // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 81:59:@9583.4]
    .clock(cycles_x538_outr_UnitPipe_DenseTransfer_clock),
    .reset(cycles_x538_outr_UnitPipe_DenseTransfer_reset),
    .io_enable(cycles_x538_outr_UnitPipe_DenseTransfer_io_enable),
    .io_count(cycles_x538_outr_UnitPipe_DenseTransfer_io_count)
  );
  InstrumentationCounter iters_x538_outr_UnitPipe_DenseTransfer ( // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 82:58:@9586.4]
    .clock(iters_x538_outr_UnitPipe_DenseTransfer_clock),
    .reset(iters_x538_outr_UnitPipe_DenseTransfer_reset),
    .io_enable(iters_x538_outr_UnitPipe_DenseTransfer_io_enable),
    .io_count(iters_x538_outr_UnitPipe_DenseTransfer_io_count)
  );
  x475_fifo x475_fifo ( // @[m_x475_fifo.scala 27:22:@9599.4]
    .clock(x475_fifo_clock),
    .reset(x475_fifo_reset),
    .io_rPort_0_en_0(x475_fifo_io_rPort_0_en_0),
    .io_rPort_0_output_0(x475_fifo_io_rPort_0_output_0),
    .io_wPort_0_data_0(x475_fifo_io_wPort_0_data_0),
    .io_wPort_0_en_0(x475_fifo_io_wPort_0_en_0),
    .io_full(x475_fifo_io_full),
    .io_empty(x475_fifo_io_empty),
    .io_active_0_in(x475_fifo_io_active_0_in),
    .io_active_0_out(x475_fifo_io_active_0_out)
  );
  x478_ctrchain x478_ctrchain ( // @[SpatialBlocks.scala 37:22:@9625.4]
    .clock(x478_ctrchain_clock),
    .reset(x478_ctrchain_reset),
    .io_input_reset(x478_ctrchain_io_input_reset),
    .io_input_enable(x478_ctrchain_io_input_enable),
    .io_output_counts_0(x478_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x478_ctrchain_io_output_oobs_0),
    .io_output_done(x478_ctrchain_io_output_done)
  );
  x499_inr_Foreach_sm x499_inr_Foreach_sm ( // @[sm_x499_inr_Foreach.scala 34:18:@9678.4]
    .clock(x499_inr_Foreach_sm_clock),
    .reset(x499_inr_Foreach_sm_reset),
    .io_enable(x499_inr_Foreach_sm_io_enable),
    .io_done(x499_inr_Foreach_sm_io_done),
    .io_doneLatch(x499_inr_Foreach_sm_io_doneLatch),
    .io_rst(x499_inr_Foreach_sm_io_rst),
    .io_ctrDone(x499_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x499_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x499_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x499_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x499_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x499_inr_Foreach_sm_io_backpressure),
    .io_break(x499_inr_Foreach_sm_io_break)
  );
  x499_inr_Foreach_iiCtr x499_inr_Foreach_iiCtr ( // @[sm_x499_inr_Foreach.scala 35:21:@9703.4]
    .clock(x499_inr_Foreach_iiCtr_clock),
    .reset(x499_inr_Foreach_iiCtr_reset),
    .io_input_enable(x499_inr_Foreach_iiCtr_io_input_enable),
    .io_input_reset(x499_inr_Foreach_iiCtr_io_input_reset),
    .io_output_issue(x499_inr_Foreach_iiCtr_io_output_issue),
    .io_output_done(x499_inr_Foreach_iiCtr_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@9707.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@9716.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@9759.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@9767.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1 x499_inr_Foreach_kernelx499_inr_Foreach_concrete1 ( // @[sm_x499_inr_Foreach.scala 135:24:@9802.4]
    .clock(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_clock),
    .reset(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_reset),
    .io_in_x468_A_dram_number(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x468_A_dram_number),
    .io_in_x475_fifo_wPort_0_data_0(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_wPort_0_data_0),
    .io_in_x475_fifo_wPort_0_en_0(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_wPort_0_en_0),
    .io_in_x475_fifo_full(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_full),
    .io_in_x475_fifo_active_0_in(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_active_0_in),
    .io_in_x475_fifo_active_0_out(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_active_0_out),
    .io_in_x474_ready(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_ready),
    .io_in_x474_valid(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_valid),
    .io_in_x474_bits_addr(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_bits_addr),
    .io_in_x474_bits_size(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_bits_size),
    .io_in_instrctrs_2_cycs(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_instrctrs_2_cycs),
    .io_in_instrctrs_2_iters(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_instrctrs_2_iters),
    .io_in_instrctrs_2_stalls(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_instrctrs_2_stalls),
    .io_in_instrctrs_2_idles(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_instrctrs_2_idles),
    .io_sigsIn_done(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_iiIssue(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_iiIssue),
    .io_sigsIn_backpressure(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_rr)
  );
  x478_ctrchain x502_ctrchain ( // @[SpatialBlocks.scala 37:22:@10007.4]
    .clock(x502_ctrchain_clock),
    .reset(x502_ctrchain_reset),
    .io_input_reset(x502_ctrchain_io_input_reset),
    .io_input_enable(x502_ctrchain_io_input_enable),
    .io_output_counts_0(x502_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x502_ctrchain_io_output_oobs_0),
    .io_output_done(x502_ctrchain_io_output_done)
  );
  x537_outr_Foreach_sm x537_outr_Foreach_sm ( // @[sm_x537_outr_Foreach.scala 34:18:@10065.4]
    .clock(x537_outr_Foreach_sm_clock),
    .reset(x537_outr_Foreach_sm_reset),
    .io_enable(x537_outr_Foreach_sm_io_enable),
    .io_done(x537_outr_Foreach_sm_io_done),
    .io_ctrDone(x537_outr_Foreach_sm_io_ctrDone),
    .io_ctrInc(x537_outr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x537_outr_Foreach_sm_io_ctrRst),
    .io_parentAck(x537_outr_Foreach_sm_io_parentAck),
    .io_doneIn_0(x537_outr_Foreach_sm_io_doneIn_0),
    .io_doneIn_1(x537_outr_Foreach_sm_io_doneIn_1),
    .io_maskIn_0(x537_outr_Foreach_sm_io_maskIn_0),
    .io_maskIn_1(x537_outr_Foreach_sm_io_maskIn_1),
    .io_enableOut_0(x537_outr_Foreach_sm_io_enableOut_0),
    .io_enableOut_1(x537_outr_Foreach_sm_io_enableOut_1),
    .io_childAck_0(x537_outr_Foreach_sm_io_childAck_0),
    .io_childAck_1(x537_outr_Foreach_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@10099.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@10144.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@10152.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1 x537_outr_Foreach_kernelx537_outr_Foreach_concrete1 ( // @[sm_x537_outr_Foreach.scala 115:24:@10187.4]
    .clock(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_clock),
    .reset(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_reset),
    .io_in_x472_A_sram_1_wPort_0_ofs_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0),
    .io_in_x472_A_sram_1_wPort_0_data_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_data_0),
    .io_in_x472_A_sram_1_wPort_0_en_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_en_0),
    .io_in_x475_fifo_rPort_0_en_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_rPort_0_en_0),
    .io_in_x475_fifo_rPort_0_output_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_rPort_0_output_0),
    .io_in_x475_fifo_empty(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_empty),
    .io_in_x471_A_sram_0_wPort_0_ofs_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0),
    .io_in_x471_A_sram_0_wPort_0_data_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_data_0),
    .io_in_x471_A_sram_0_wPort_0_en_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_en_0),
    .io_in_x476_ready(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_ready),
    .io_in_x476_valid(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_valid),
    .io_in_x476_bits_rdata_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_bits_rdata_0),
    .io_in_x473_A_sram_2_wPort_0_ofs_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0),
    .io_in_x473_A_sram_2_wPort_0_data_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_data_0),
    .io_in_x473_A_sram_2_wPort_0_en_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_en_0),
    .io_in_instrctrs_3_cycs(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_3_cycs),
    .io_in_instrctrs_3_iters(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_3_iters),
    .io_in_instrctrs_4_cycs(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_4_cycs),
    .io_in_instrctrs_4_iters(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_4_iters),
    .io_in_instrctrs_4_stalls(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_4_stalls),
    .io_in_instrctrs_4_idles(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_4_idles),
    .io_in_instrctrs_5_cycs(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_5_cycs),
    .io_in_instrctrs_5_iters(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_5_iters),
    .io_in_instrctrs_5_stalls(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_5_stalls),
    .io_in_instrctrs_5_idles(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_5_idles),
    .io_sigsIn_done(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smEnableOuts_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsOut_smDoneIn_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smMaskIn_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0),
    .io_sigsOut_smMaskIn_1(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1),
    .io_rr(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_rr)
  );
  assign _T_546 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@9590.4]
  assign _T_616 = RetimeWrapper_io_out; // @[package.scala 96:25:@9712.4 package.scala 96:25:@9713.4]
  assign _T_622 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@9721.4 package.scala 96:25:@9722.4]
  assign _T_625 = ~ _T_622; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 93:41:@9724.4]
  assign _T_626 = ~ x475_fifo_io_active_0_out; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 93:68:@9725.4]
  assign _T_627 = _T_625 | _T_626; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 93:66:@9726.4]
  assign _T_628 = _T_627 & io_in_x474_ready; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 93:96:@9727.4]
  assign _T_642 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@9764.4 package.scala 96:25:@9765.4]
  assign _T_648 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@9772.4 package.scala 96:25:@9773.4]
  assign _T_651 = ~ _T_648; // @[SpatialBlocks.scala 137:99:@9775.4]
  assign _T_653 = x499_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 156:36:@9784.4]
  assign _T_654 = ~ x499_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 156:78:@9785.4]
  assign x499_inr_Foreach_mySignalsIn_iiDone = x499_inr_Foreach_iiCtr_io_output_done; // @[SpatialBlocks.scala 157:126:@9792.4]
  assign _T_725 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@10104.4 package.scala 96:25:@10105.4]
  assign _T_742 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@10149.4 package.scala 96:25:@10150.4]
  assign _T_748 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@10157.4 package.scala 96:25:@10158.4]
  assign _T_751 = ~ _T_748; // @[SpatialBlocks.scala 137:99:@10160.4]
  assign io_in_x472_A_sram_1_wPort_0_ofs_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@10388.4]
  assign io_in_x472_A_sram_1_wPort_0_data_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@10387.4]
  assign io_in_x472_A_sram_1_wPort_0_en_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@10383.4]
  assign io_in_x471_A_sram_0_wPort_0_ofs_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@10408.4]
  assign io_in_x471_A_sram_0_wPort_0_data_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@10407.4]
  assign io_in_x471_A_sram_0_wPort_0_en_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@10403.4]
  assign io_in_x476_ready = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_ready; // @[sm_x537_outr_Foreach.scala 60:23:@10412.4]
  assign io_in_x473_A_sram_2_wPort_0_ofs_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@10418.4]
  assign io_in_x473_A_sram_2_wPort_0_data_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@10417.4]
  assign io_in_x473_A_sram_2_wPort_0_en_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@10413.4]
  assign io_in_x474_valid = x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_valid; // @[sm_x499_inr_Foreach.scala 55:23:@9974.4]
  assign io_in_x474_bits_addr = x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_bits_addr; // @[sm_x499_inr_Foreach.scala 55:23:@9973.4]
  assign io_in_x474_bits_size = x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_bits_size; // @[sm_x499_inr_Foreach.scala 55:23:@9972.4]
  assign io_in_instrctrs_1_cycs = cycles_x538_outr_UnitPipe_DenseTransfer_io_count; // @[Ledger.scala 293:21:@9595.4]
  assign io_in_instrctrs_1_iters = iters_x538_outr_UnitPipe_DenseTransfer_io_count; // @[Ledger.scala 294:22:@9596.4]
  assign io_in_instrctrs_2_cycs = x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_instrctrs_2_cycs; // @[Ledger.scala 302:78:@9979.4]
  assign io_in_instrctrs_2_iters = x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_instrctrs_2_iters; // @[Ledger.scala 302:78:@9978.4]
  assign io_in_instrctrs_2_stalls = x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_instrctrs_2_stalls; // @[Ledger.scala 302:78:@9977.4]
  assign io_in_instrctrs_2_idles = x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_instrctrs_2_idles; // @[Ledger.scala 302:78:@9976.4]
  assign io_in_instrctrs_3_cycs = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_3_cycs; // @[Ledger.scala 302:78:@10423.4]
  assign io_in_instrctrs_3_iters = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_3_iters; // @[Ledger.scala 302:78:@10422.4]
  assign io_in_instrctrs_4_cycs = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_4_cycs; // @[Ledger.scala 302:78:@10427.4]
  assign io_in_instrctrs_4_iters = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_4_iters; // @[Ledger.scala 302:78:@10426.4]
  assign io_in_instrctrs_4_stalls = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_4_stalls; // @[Ledger.scala 302:78:@10425.4]
  assign io_in_instrctrs_4_idles = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_4_idles; // @[Ledger.scala 302:78:@10424.4]
  assign io_in_instrctrs_5_cycs = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_5_cycs; // @[Ledger.scala 302:78:@10431.4]
  assign io_in_instrctrs_5_iters = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_5_iters; // @[Ledger.scala 302:78:@10430.4]
  assign io_in_instrctrs_5_stalls = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_5_stalls; // @[Ledger.scala 302:78:@10429.4]
  assign io_in_instrctrs_5_idles = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_instrctrs_5_idles; // @[Ledger.scala 302:78:@10428.4]
  assign io_sigsOut_smDoneIn_0 = x499_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@9782.4]
  assign io_sigsOut_smDoneIn_1 = x537_outr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@10167.4]
  assign io_sigsOut_smCtrCopyDone_0 = x499_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 170:140:@9801.4]
  assign io_sigsOut_smCtrCopyDone_1 = x537_outr_Foreach_sm_io_done; // @[SpatialBlocks.scala 170:140:@10186.4]
  assign cycles_x538_outr_UnitPipe_DenseTransfer_clock = clock; // @[:@9584.4]
  assign cycles_x538_outr_UnitPipe_DenseTransfer_reset = reset; // @[:@9585.4]
  assign cycles_x538_outr_UnitPipe_DenseTransfer_io_enable = io_sigsIn_baseEn; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 83:57:@9589.4]
  assign iters_x538_outr_UnitPipe_DenseTransfer_clock = clock; // @[:@9587.4]
  assign iters_x538_outr_UnitPipe_DenseTransfer_reset = reset; // @[:@9588.4]
  assign iters_x538_outr_UnitPipe_DenseTransfer_io_enable = io_sigsIn_done & _T_549; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 84:56:@9594.4]
  assign x475_fifo_clock = clock; // @[:@9600.4]
  assign x475_fifo_reset = reset; // @[:@9601.4]
  assign x475_fifo_io_rPort_0_en_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@10400.4]
  assign x475_fifo_io_wPort_0_data_0 = x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@9969.4]
  assign x475_fifo_io_wPort_0_en_0 = x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@9965.4]
  assign x475_fifo_io_active_0_in = x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_active_0_in; // @[MemInterfaceType.scala 167:86:@9964.4]
  assign x478_ctrchain_clock = clock; // @[:@9626.4]
  assign x478_ctrchain_reset = reset; // @[:@9627.4]
  assign x478_ctrchain_io_input_reset = x499_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@9800.4]
  assign x478_ctrchain_io_input_enable = x499_inr_Foreach_sm_io_ctrInc & x499_inr_Foreach_mySignalsIn_iiDone; // @[SpatialBlocks.scala 158:42:@9799.4]
  assign x499_inr_Foreach_sm_clock = clock; // @[:@9679.4]
  assign x499_inr_Foreach_sm_reset = reset; // @[:@9680.4]
  assign x499_inr_Foreach_sm_io_enable = _T_642 & _T_651; // @[SpatialBlocks.scala 139:18:@9779.4]
  assign x499_inr_Foreach_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 133:15:@9754.4]
  assign x499_inr_Foreach_sm_io_ctrDone = io_rr ? _T_616 : 1'h0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 92:38:@9715.4]
  assign x499_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@9781.4]
  assign x499_inr_Foreach_sm_io_backpressure = _T_628 | x499_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 132:24:@9753.4]
  assign x499_inr_Foreach_sm_io_break = 1'h0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 96:36:@9734.4]
  assign x499_inr_Foreach_iiCtr_clock = clock; // @[:@9704.4]
  assign x499_inr_Foreach_iiCtr_reset = reset; // @[:@9705.4]
  assign x499_inr_Foreach_iiCtr_io_input_enable = _T_653 & _T_654; // @[SpatialBlocks.scala 157:27:@9788.4]
  assign x499_inr_Foreach_iiCtr_io_input_reset = x499_inr_Foreach_sm_io_rst | x499_inr_Foreach_sm_io_parentAck; // @[SpatialBlocks.scala 157:63:@9790.4]
  assign RetimeWrapper_clock = clock; // @[:@9708.4]
  assign RetimeWrapper_reset = reset; // @[:@9709.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@9711.4]
  assign RetimeWrapper_io_in = x478_ctrchain_io_output_done; // @[package.scala 94:16:@9710.4]
  assign RetimeWrapper_1_clock = clock; // @[:@9717.4]
  assign RetimeWrapper_1_reset = reset; // @[:@9718.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@9720.4]
  assign RetimeWrapper_1_io_in = x475_fifo_io_full; // @[package.scala 94:16:@9719.4]
  assign RetimeWrapper_2_clock = clock; // @[:@9760.4]
  assign RetimeWrapper_2_reset = reset; // @[:@9761.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@9763.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@9762.4]
  assign RetimeWrapper_3_clock = clock; // @[:@9768.4]
  assign RetimeWrapper_3_reset = reset; // @[:@9769.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@9771.4]
  assign RetimeWrapper_3_io_in = x499_inr_Foreach_sm_io_done; // @[package.scala 94:16:@9770.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_clock = clock; // @[:@9803.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_reset = reset; // @[:@9804.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x468_A_dram_number = io_in_x468_A_dram_number; // @[sm_x499_inr_Foreach.scala 53:30:@9956.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_full = x475_fifo_io_full; // @[MemInterfaceType.scala 159:15:@9959.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_active_0_out = x475_fifo_io_active_0_out; // @[MemInterfaceType.scala 158:75:@9957.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_ready = io_in_x474_ready; // @[sm_x499_inr_Foreach.scala 55:23:@9975.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_done = x499_inr_Foreach_sm_io_done; // @[sm_x499_inr_Foreach.scala 141:22:@9999.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_iiIssue = x499_inr_Foreach_iiCtr_io_output_issue; // @[sm_x499_inr_Foreach.scala 141:22:@9996.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_628 | x499_inr_Foreach_sm_io_doneLatch; // @[sm_x499_inr_Foreach.scala 141:22:@9994.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_653 & _T_654; // @[sm_x499_inr_Foreach.scala 141:22:@9992.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_baseEn = _T_642 & _T_651; // @[sm_x499_inr_Foreach.scala 141:22:@9991.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_break = x499_inr_Foreach_sm_io_break; // @[sm_x499_inr_Foreach.scala 141:22:@9990.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{23{x478_ctrchain_io_output_counts_0[8]}},x478_ctrchain_io_output_counts_0}; // @[sm_x499_inr_Foreach.scala 141:22:@9985.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x478_ctrchain_io_output_oobs_0; // @[sm_x499_inr_Foreach.scala 141:22:@9984.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x499_inr_Foreach.scala 140:18:@9980.4]
  assign x502_ctrchain_clock = clock; // @[:@10008.4]
  assign x502_ctrchain_reset = reset; // @[:@10009.4]
  assign x502_ctrchain_io_input_reset = x537_outr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@10185.4]
  assign x502_ctrchain_io_input_enable = x537_outr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 158:42:@10184.4]
  assign x537_outr_Foreach_sm_clock = clock; // @[:@10066.4]
  assign x537_outr_Foreach_sm_reset = reset; // @[:@10067.4]
  assign x537_outr_Foreach_sm_io_enable = _T_742 & _T_751; // @[SpatialBlocks.scala 139:18:@10164.4]
  assign x537_outr_Foreach_sm_io_ctrDone = io_rr ? _T_725 : 1'h0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 105:39:@10107.4]
  assign x537_outr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 141:21:@10166.4]
  assign x537_outr_Foreach_sm_io_doneIn_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@10134.4]
  assign x537_outr_Foreach_sm_io_doneIn_1 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:72:@10135.4]
  assign x537_outr_Foreach_sm_io_maskIn_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0; // @[SpatialBlocks.scala 131:72:@10136.4]
  assign x537_outr_Foreach_sm_io_maskIn_1 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1; // @[SpatialBlocks.scala 131:72:@10137.4]
  assign RetimeWrapper_4_clock = clock; // @[:@10100.4]
  assign RetimeWrapper_4_reset = reset; // @[:@10101.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@10103.4]
  assign RetimeWrapper_4_io_in = x502_ctrchain_io_output_done; // @[package.scala 94:16:@10102.4]
  assign RetimeWrapper_5_clock = clock; // @[:@10145.4]
  assign RetimeWrapper_5_reset = reset; // @[:@10146.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@10148.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@10147.4]
  assign RetimeWrapper_6_clock = clock; // @[:@10153.4]
  assign RetimeWrapper_6_reset = reset; // @[:@10154.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@10156.4]
  assign RetimeWrapper_6_io_in = x537_outr_Foreach_sm_io_done; // @[package.scala 94:16:@10155.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_clock = clock; // @[:@10188.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_reset = reset; // @[:@10189.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_rPort_0_output_0 = x475_fifo_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@10398.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_empty = x475_fifo_io_empty; // @[MemInterfaceType.scala 161:16:@10394.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_valid = io_in_x476_valid; // @[sm_x537_outr_Foreach.scala 60:23:@10411.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_bits_rdata_0 = io_in_x476_bits_rdata_0; // @[sm_x537_outr_Foreach.scala 60:23:@10410.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_done = x537_outr_Foreach_sm_io_done; // @[sm_x537_outr_Foreach.scala 121:22:@10454.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_baseEn = _T_742 & _T_751; // @[sm_x537_outr_Foreach.scala 121:22:@10446.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0 = x537_outr_Foreach_sm_io_enableOut_0; // @[sm_x537_outr_Foreach.scala 121:22:@10442.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1 = x537_outr_Foreach_sm_io_enableOut_1; // @[sm_x537_outr_Foreach.scala 121:22:@10443.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0 = x537_outr_Foreach_sm_io_childAck_0; // @[sm_x537_outr_Foreach.scala 121:22:@10438.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1 = x537_outr_Foreach_sm_io_childAck_1; // @[sm_x537_outr_Foreach.scala 121:22:@10439.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{23{x502_ctrchain_io_output_counts_0[8]}},x502_ctrchain_io_output_counts_0}; // @[sm_x537_outr_Foreach.scala 121:22:@10437.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x502_ctrchain_io_output_oobs_0; // @[sm_x537_outr_Foreach.scala 121:22:@10436.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_rr = io_rr; // @[sm_x537_outr_Foreach.scala 120:18:@10432.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_549 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_549 <= 1'h0;
    end else begin
      _T_549 <= _T_546;
    end
  end
endmodule
module x668_outr_Foreach_sm( // @[:@11104.2]
  input   clock, // @[:@11105.4]
  input   reset, // @[:@11106.4]
  input   io_enable, // @[:@11107.4]
  output  io_done, // @[:@11107.4]
  input   io_ctrDone, // @[:@11107.4]
  output  io_ctrInc, // @[:@11107.4]
  output  io_ctrRst, // @[:@11107.4]
  input   io_parentAck, // @[:@11107.4]
  input   io_doneIn_0, // @[:@11107.4]
  input   io_doneIn_1, // @[:@11107.4]
  input   io_maskIn_0, // @[:@11107.4]
  input   io_maskIn_1, // @[:@11107.4]
  output  io_enableOut_0, // @[:@11107.4]
  output  io_enableOut_1, // @[:@11107.4]
  output  io_childAck_0, // @[:@11107.4]
  output  io_childAck_1 // @[:@11107.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@11110.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@11110.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@11110.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@11110.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@11110.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@11110.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@11113.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@11113.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@11113.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@11113.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@11113.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@11113.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@11116.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@11116.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@11116.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@11116.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@11116.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@11116.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@11119.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@11119.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@11119.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@11119.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@11119.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@11119.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@11148.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@11148.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@11148.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@11148.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@11148.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@11148.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@11151.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@11151.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@11151.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@11151.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@11151.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@11151.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@11192.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@11192.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@11192.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@11192.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@11192.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@11218.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@11218.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@11218.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@11218.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@11218.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@11238.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@11238.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@11238.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@11238.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@11238.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@11287.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@11287.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@11287.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@11287.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@11287.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@11304.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@11304.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@11304.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@11304.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@11304.4]
  wire  allDone; // @[Controllers.scala 80:47:@11122.4]
  wire  _T_128; // @[Controllers.scala 102:95:@11178.4]
  wire  _T_127; // @[Controllers.scala 101:55:@11177.4]
  wire  _T_132; // @[package.scala 96:25:@11184.4 package.scala 96:25:@11185.4]
  wire  _T_135; // @[Controllers.scala 102:142:@11187.4]
  wire  _T_136; // @[Controllers.scala 102:138:@11188.4]
  wire  _T_137; // @[Controllers.scala 102:123:@11189.4]
  wire  _T_138; // @[Controllers.scala 102:112:@11190.4]
  wire  _T_139; // @[Controllers.scala 102:95:@11191.4]
  wire  _T_143; // @[package.scala 96:25:@11197.4 package.scala 96:25:@11198.4]
  wire  _T_146; // @[Controllers.scala 102:142:@11200.4]
  wire  _T_147; // @[Controllers.scala 102:138:@11201.4]
  wire  _T_148; // @[Controllers.scala 102:123:@11202.4]
  wire  _T_149; // @[Controllers.scala 102:112:@11203.4]
  wire  synchronize; // @[Controllers.scala 102:164:@11204.4]
  wire  _T_152; // @[Controllers.scala 105:33:@11206.4]
  wire  _T_154; // @[Controllers.scala 105:54:@11207.4]
  wire  _T_155; // @[Controllers.scala 105:52:@11208.4]
  wire  _T_161; // @[Controllers.scala 107:51:@11215.4]
  wire  _T_164; // @[Controllers.scala 107:64:@11217.4]
  wire  _T_168; // @[package.scala 96:25:@11223.4 package.scala 96:25:@11224.4]
  wire  _T_172; // @[Controllers.scala 107:89:@11226.4]
  wire  _T_173; // @[Controllers.scala 107:86:@11227.4]
  wire  _T_174; // @[Controllers.scala 107:108:@11228.4]
  wire  _T_189; // @[Controllers.scala 114:49:@11246.4]
  wire  _T_192; // @[Controllers.scala 115:57:@11250.4]
  wire  _T_203; // @[Controllers.scala 213:68:@11265.4]
  wire  _T_204; // @[Controllers.scala 213:92:@11266.4]
  wire  _T_205; // @[Controllers.scala 213:90:@11267.4]
  wire  _T_206; // @[Controllers.scala 213:115:@11268.4]
  wire  _T_207; // @[Controllers.scala 213:132:@11269.4]
  wire  _T_208; // @[Controllers.scala 213:130:@11270.4]
  wire  _T_209; // @[Controllers.scala 213:156:@11271.4]
  wire  _T_211; // @[Controllers.scala 213:68:@11274.4]
  wire  _T_212; // @[Controllers.scala 213:92:@11275.4]
  wire  _T_213; // @[Controllers.scala 213:90:@11276.4]
  wire  _T_214; // @[Controllers.scala 213:115:@11277.4]
  wire  _T_220; // @[package.scala 100:49:@11282.4]
  reg  _T_223; // @[package.scala 48:56:@11283.4]
  reg [31:0] _RAND_0;
  wire  _T_224; // @[package.scala 100:41:@11285.4]
  reg  _T_237; // @[package.scala 48:56:@11301.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@11110.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@11113.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@11116.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@11119.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@11148.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@11151.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@11179.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@11192.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@11218.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@11238.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@11287.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@11304.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@11122.4]
  assign _T_128 = active_0_io_output == iterDone_0_io_output; // @[Controllers.scala 102:95:@11178.4]
  assign _T_127 = iterDone_0_io_output | iterDone_1_io_output; // @[Controllers.scala 101:55:@11177.4]
  assign _T_132 = RetimeWrapper_io_out; // @[package.scala 96:25:@11184.4 package.scala 96:25:@11185.4]
  assign _T_135 = ~ _T_132; // @[Controllers.scala 102:142:@11187.4]
  assign _T_136 = active_0_io_output == _T_135; // @[Controllers.scala 102:138:@11188.4]
  assign _T_137 = _T_127 & _T_136; // @[Controllers.scala 102:123:@11189.4]
  assign _T_138 = _T_128 | _T_137; // @[Controllers.scala 102:112:@11190.4]
  assign _T_139 = active_1_io_output == iterDone_1_io_output; // @[Controllers.scala 102:95:@11191.4]
  assign _T_143 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@11197.4 package.scala 96:25:@11198.4]
  assign _T_146 = ~ _T_143; // @[Controllers.scala 102:142:@11200.4]
  assign _T_147 = active_1_io_output == _T_146; // @[Controllers.scala 102:138:@11201.4]
  assign _T_148 = _T_127 & _T_147; // @[Controllers.scala 102:123:@11202.4]
  assign _T_149 = _T_139 | _T_148; // @[Controllers.scala 102:112:@11203.4]
  assign synchronize = _T_138 & _T_149; // @[Controllers.scala 102:164:@11204.4]
  assign _T_152 = done_0_io_output == 1'h0; // @[Controllers.scala 105:33:@11206.4]
  assign _T_154 = io_ctrDone == 1'h0; // @[Controllers.scala 105:54:@11207.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 105:52:@11208.4]
  assign _T_161 = synchronize == 1'h0; // @[Controllers.scala 107:51:@11215.4]
  assign _T_164 = _T_161 & _T_152; // @[Controllers.scala 107:64:@11217.4]
  assign _T_168 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@11223.4 package.scala 96:25:@11224.4]
  assign _T_172 = _T_168 == 1'h0; // @[Controllers.scala 107:89:@11226.4]
  assign _T_173 = _T_164 & _T_172; // @[Controllers.scala 107:86:@11227.4]
  assign _T_174 = _T_173 & io_enable; // @[Controllers.scala 107:108:@11228.4]
  assign _T_189 = synchronize & active_0_io_output; // @[Controllers.scala 114:49:@11246.4]
  assign _T_192 = done_0_io_output & synchronize; // @[Controllers.scala 115:57:@11250.4]
  assign _T_203 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@11265.4]
  assign _T_204 = ~ iterDone_0_io_output; // @[Controllers.scala 213:92:@11266.4]
  assign _T_205 = _T_203 & _T_204; // @[Controllers.scala 213:90:@11267.4]
  assign _T_206 = _T_205 & io_maskIn_0; // @[Controllers.scala 213:115:@11268.4]
  assign _T_207 = ~ allDone; // @[Controllers.scala 213:132:@11269.4]
  assign _T_208 = _T_206 & _T_207; // @[Controllers.scala 213:130:@11270.4]
  assign _T_209 = ~ io_ctrDone; // @[Controllers.scala 213:156:@11271.4]
  assign _T_211 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@11274.4]
  assign _T_212 = ~ iterDone_1_io_output; // @[Controllers.scala 213:92:@11275.4]
  assign _T_213 = _T_211 & _T_212; // @[Controllers.scala 213:90:@11276.4]
  assign _T_214 = _T_213 & io_maskIn_1; // @[Controllers.scala 213:115:@11277.4]
  assign _T_220 = allDone == 1'h0; // @[package.scala 100:49:@11282.4]
  assign _T_224 = allDone & _T_223; // @[package.scala 100:41:@11285.4]
  assign io_done = RetimeWrapper_5_io_out; // @[Controllers.scala 245:13:@11311.4]
  assign io_ctrInc = iterDone_0_io_output & synchronize; // @[Controllers.scala 98:17:@11176.4]
  assign io_ctrRst = RetimeWrapper_4_io_out; // @[Controllers.scala 215:13:@11294.4]
  assign io_enableOut_0 = _T_208 & _T_209; // @[Controllers.scala 213:55:@11273.4]
  assign io_enableOut_1 = _T_214 & _T_207; // @[Controllers.scala 213:55:@11281.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@11262.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@11264.4]
  assign active_0_clock = clock; // @[:@11111.4]
  assign active_0_reset = reset; // @[:@11112.4]
  assign active_0_io_input_set = _T_155 & io_enable; // @[Controllers.scala 105:30:@11211.4]
  assign active_0_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 106:32:@11214.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@11125.4]
  assign active_1_clock = clock; // @[:@11114.4]
  assign active_1_reset = reset; // @[:@11115.4]
  assign active_1_io_input_set = _T_189 & io_enable; // @[Controllers.scala 114:32:@11249.4]
  assign active_1_io_input_reset = _T_192 | io_parentAck; // @[Controllers.scala 115:34:@11253.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@11126.4]
  assign done_0_clock = clock; // @[:@11117.4]
  assign done_0_reset = reset; // @[:@11118.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 108:28:@11236.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@11137.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@11127.4]
  assign done_1_clock = clock; // @[:@11120.4]
  assign done_1_reset = reset; // @[:@11121.4]
  assign done_1_io_input_set = done_0_io_output & synchronize; // @[Controllers.scala 117:30:@11260.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@11146.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@11128.4]
  assign iterDone_0_clock = clock; // @[:@11149.4]
  assign iterDone_0_reset = reset; // @[:@11150.4]
  assign iterDone_0_io_input_set = io_doneIn_0 | _T_174; // @[Controllers.scala 107:32:@11232.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@11164.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@11154.4]
  assign iterDone_1_clock = clock; // @[:@11152.4]
  assign iterDone_1_reset = reset; // @[:@11153.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 116:34:@11255.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@11173.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@11155.4]
  assign RetimeWrapper_clock = clock; // @[:@11180.4]
  assign RetimeWrapper_reset = reset; // @[:@11181.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@11183.4]
  assign RetimeWrapper_io_in = io_maskIn_0; // @[package.scala 94:16:@11182.4]
  assign RetimeWrapper_1_clock = clock; // @[:@11193.4]
  assign RetimeWrapper_1_reset = reset; // @[:@11194.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@11196.4]
  assign RetimeWrapper_1_io_in = io_maskIn_1; // @[package.scala 94:16:@11195.4]
  assign RetimeWrapper_2_clock = clock; // @[:@11219.4]
  assign RetimeWrapper_2_reset = reset; // @[:@11220.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@11222.4]
  assign RetimeWrapper_2_io_in = io_maskIn_0; // @[package.scala 94:16:@11221.4]
  assign RetimeWrapper_3_clock = clock; // @[:@11239.4]
  assign RetimeWrapper_3_reset = reset; // @[:@11240.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@11242.4]
  assign RetimeWrapper_3_io_in = synchronize & iterDone_0_io_output; // @[package.scala 94:16:@11241.4]
  assign RetimeWrapper_4_clock = clock; // @[:@11288.4]
  assign RetimeWrapper_4_reset = reset; // @[:@11289.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@11291.4]
  assign RetimeWrapper_4_io_in = _T_224 | io_parentAck; // @[package.scala 94:16:@11290.4]
  assign RetimeWrapper_5_clock = clock; // @[:@11305.4]
  assign RetimeWrapper_5_reset = reset; // @[:@11306.4]
  assign RetimeWrapper_5_io_flow = io_enable; // @[package.scala 95:18:@11308.4]
  assign RetimeWrapper_5_io_in = allDone & _T_237; // @[package.scala 94:16:@11307.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_223 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_237 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_223 <= 1'h0;
    end else begin
      _T_223 <= _T_220;
    end
    if (reset) begin
      _T_237 <= 1'h0;
    end else begin
      _T_237 <= _T_220;
    end
  end
endmodule
module RetimeWrapper_97( // @[:@11811.2]
  input         clock, // @[:@11812.4]
  input         reset, // @[:@11813.4]
  input         io_flow, // @[:@11814.4]
  input  [31:0] io_in, // @[:@11814.4]
  output [31:0] io_out // @[:@11814.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@11816.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@11816.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@11816.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@11816.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@11816.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@11816.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@11816.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@11829.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@11828.4]
  assign sr_init = 32'h1; // @[RetimeShiftRegister.scala 19:16:@11827.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@11826.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@11825.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@11823.4]
endmodule
module NBufCtr( // @[:@11831.2]
  input         clock, // @[:@11832.4]
  input         reset, // @[:@11833.4]
  input         io_input_countUp, // @[:@11834.4]
  input         io_input_enable, // @[:@11834.4]
  output [31:0] io_output_count // @[:@11834.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@11871.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@11871.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@11871.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@11871.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@11871.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@11876.4 package.scala 96:25:@11877.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@11837.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@11838.4]
  wire  _T_21; // @[Counter.scala 49:55:@11839.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@11840.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@11841.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@11842.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@11843.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@11844.4]
  wire  _T_33; // @[Counter.scala 51:52:@11848.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@11849.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@11850.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@11851.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@11852.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@11853.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@11854.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@11855.4]
  wire  _T_45; // @[Counter.scala 52:70:@11856.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@11858.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@11859.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@11860.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@11861.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@11862.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@11863.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@11866.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@11867.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@11869.4]
  RetimeWrapper_97 RetimeWrapper ( // @[package.scala 93:22:@11871.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@11876.4 package.scala 96:25:@11877.4]
  assign _T_18 = {{1'd0}, _T_66}; // @[Counter.scala 49:32:@11837.4]
  assign _T_19 = _T_18[31:0]; // @[Counter.scala 49:32:@11838.4]
  assign _T_21 = _T_19 >= 32'h2; // @[Counter.scala 49:55:@11839.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@11840.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh2); // @[Counter.scala 49:91:@11841.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh2); // @[Counter.scala 49:91:@11842.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@11843.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@11844.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@11848.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@11849.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@11850.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@11851.4]
  assign _T_39 = _T_33 ? 32'h1 : _T_38; // @[Counter.scala 51:47:@11852.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@11853.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@11854.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@11855.4]
  assign _T_45 = _T_43 >= 32'h2; // @[Counter.scala 52:70:@11856.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 52:121:@11858.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 52:121:@11859.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@11860.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@11861.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@11862.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@11863.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@11866.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@11867.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@11869.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@11879.4]
  assign RetimeWrapper_clock = clock; // @[:@11872.4]
  assign RetimeWrapper_reset = reset; // @[:@11873.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@11875.4]
  assign RetimeWrapper_io_in = reset ? 32'h1 : _T_62; // @[package.scala 94:16:@11874.4]
endmodule
module NBufCtr_2( // @[:@11995.2]
  input         clock, // @[:@11996.4]
  input         reset, // @[:@11997.4]
  input         io_input_countUp, // @[:@11998.4]
  input         io_input_enable, // @[:@11998.4]
  output [31:0] io_output_count // @[:@11998.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@12035.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@12035.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@12035.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@12035.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@12035.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@12040.4 package.scala 96:25:@12041.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@12001.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@12002.4]
  wire  _T_21; // @[Counter.scala 49:55:@12003.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@12004.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@12005.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@12006.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@12007.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@12008.4]
  wire  _T_33; // @[Counter.scala 51:52:@12012.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@12013.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@12014.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@12015.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@12016.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@12017.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@12026.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@12027.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@12030.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@12031.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@12033.4]
  RetimeWrapper_97 RetimeWrapper ( // @[package.scala 93:22:@12035.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@12040.4 package.scala 96:25:@12041.4]
  assign _T_18 = _T_66 + 32'h1; // @[Counter.scala 49:32:@12001.4]
  assign _T_19 = _T_66 + 32'h1; // @[Counter.scala 49:32:@12002.4]
  assign _T_21 = _T_19 >= 32'h2; // @[Counter.scala 49:55:@12003.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@12004.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 49:91:@12005.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 49:91:@12006.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@12007.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@12008.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@12012.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@12013.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@12014.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@12015.4]
  assign _T_39 = _T_33 ? 32'h1 : _T_38; // @[Counter.scala 51:47:@12016.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@12017.4]
  assign _T_53 = {{1'd0}, _T_27}; // @[Counter.scala 52:107:@12026.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@12027.4]
  assign _T_58 = _T_21 ? _T_54 : _T_19; // @[Counter.scala 52:45:@12030.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@12031.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@12033.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@12043.4]
  assign RetimeWrapper_clock = clock; // @[:@12036.4]
  assign RetimeWrapper_reset = reset; // @[:@12037.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@12039.4]
  assign RetimeWrapper_io_in = reset ? 32'h1 : _T_62; // @[package.scala 94:16:@12038.4]
endmodule
module NBufController( // @[:@12045.2]
  input        clock, // @[:@12046.4]
  input        reset, // @[:@12047.4]
  input        io_sEn_0, // @[:@12048.4]
  input        io_sEn_1, // @[:@12048.4]
  input        io_sDone_0, // @[:@12048.4]
  input        io_sDone_1, // @[:@12048.4]
  output [2:0] io_statesInW_0, // @[:@12048.4]
  output [2:0] io_statesInR_1 // @[:@12048.4]
);
  wire  sEn_latch_0_clock; // @[NBuffers.scala 21:52:@12050.4]
  wire  sEn_latch_0_reset; // @[NBuffers.scala 21:52:@12050.4]
  wire  sEn_latch_0_io_input_set; // @[NBuffers.scala 21:52:@12050.4]
  wire  sEn_latch_0_io_input_reset; // @[NBuffers.scala 21:52:@12050.4]
  wire  sEn_latch_0_io_input_asyn_reset; // @[NBuffers.scala 21:52:@12050.4]
  wire  sEn_latch_0_io_output; // @[NBuffers.scala 21:52:@12050.4]
  wire  sEn_latch_1_clock; // @[NBuffers.scala 21:52:@12053.4]
  wire  sEn_latch_1_reset; // @[NBuffers.scala 21:52:@12053.4]
  wire  sEn_latch_1_io_input_set; // @[NBuffers.scala 21:52:@12053.4]
  wire  sEn_latch_1_io_input_reset; // @[NBuffers.scala 21:52:@12053.4]
  wire  sEn_latch_1_io_input_asyn_reset; // @[NBuffers.scala 21:52:@12053.4]
  wire  sEn_latch_1_io_output; // @[NBuffers.scala 21:52:@12053.4]
  wire  sDone_latch_0_clock; // @[NBuffers.scala 22:54:@12056.4]
  wire  sDone_latch_0_reset; // @[NBuffers.scala 22:54:@12056.4]
  wire  sDone_latch_0_io_input_set; // @[NBuffers.scala 22:54:@12056.4]
  wire  sDone_latch_0_io_input_reset; // @[NBuffers.scala 22:54:@12056.4]
  wire  sDone_latch_0_io_input_asyn_reset; // @[NBuffers.scala 22:54:@12056.4]
  wire  sDone_latch_0_io_output; // @[NBuffers.scala 22:54:@12056.4]
  wire  sDone_latch_1_clock; // @[NBuffers.scala 22:54:@12059.4]
  wire  sDone_latch_1_reset; // @[NBuffers.scala 22:54:@12059.4]
  wire  sDone_latch_1_io_input_set; // @[NBuffers.scala 22:54:@12059.4]
  wire  sDone_latch_1_io_input_reset; // @[NBuffers.scala 22:54:@12059.4]
  wire  sDone_latch_1_io_input_asyn_reset; // @[NBuffers.scala 22:54:@12059.4]
  wire  sDone_latch_1_io_output; // @[NBuffers.scala 22:54:@12059.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@12066.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@12066.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@12066.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@12066.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@12066.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@12074.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@12074.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@12074.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@12074.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@12074.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@12083.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@12083.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@12083.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@12083.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@12083.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@12091.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@12091.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@12091.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@12091.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@12091.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@12102.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@12102.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@12102.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@12102.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@12102.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@12110.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@12110.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@12110.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@12110.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@12110.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@12119.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@12119.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@12119.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@12119.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@12119.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@12127.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@12127.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@12127.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@12127.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@12127.4]
  wire  NBufCtr_clock; // @[NBuffers.scala 40:19:@12148.4]
  wire  NBufCtr_reset; // @[NBuffers.scala 40:19:@12148.4]
  wire  NBufCtr_io_input_countUp; // @[NBuffers.scala 40:19:@12148.4]
  wire  NBufCtr_io_input_enable; // @[NBuffers.scala 40:19:@12148.4]
  wire [31:0] NBufCtr_io_output_count; // @[NBuffers.scala 40:19:@12148.4]
  wire  statesInR_0_clock; // @[NBuffers.scala 50:19:@12159.4]
  wire  statesInR_0_reset; // @[NBuffers.scala 50:19:@12159.4]
  wire  statesInR_0_io_input_countUp; // @[NBuffers.scala 50:19:@12159.4]
  wire  statesInR_0_io_input_enable; // @[NBuffers.scala 50:19:@12159.4]
  wire [31:0] statesInR_0_io_output_count; // @[NBuffers.scala 50:19:@12159.4]
  wire  statesInR_1_clock; // @[NBuffers.scala 50:19:@12170.4]
  wire  statesInR_1_reset; // @[NBuffers.scala 50:19:@12170.4]
  wire  statesInR_1_io_input_countUp; // @[NBuffers.scala 50:19:@12170.4]
  wire  statesInR_1_io_input_enable; // @[NBuffers.scala 50:19:@12170.4]
  wire [31:0] statesInR_1_io_output_count; // @[NBuffers.scala 50:19:@12170.4]
  wire  _T_33; // @[NBuffers.scala 26:46:@12063.4]
  wire  _T_48; // @[NBuffers.scala 26:46:@12099.4]
  wire  anyEnabled; // @[NBuffers.scala 33:64:@12135.4]
  wire  _T_62; // @[NBuffers.scala 34:124:@12136.4]
  wire  _T_63; // @[NBuffers.scala 34:104:@12137.4]
  wire  _T_64; // @[NBuffers.scala 34:124:@12138.4]
  wire  _T_65; // @[NBuffers.scala 34:104:@12139.4]
  wire  _T_66; // @[NBuffers.scala 34:150:@12140.4]
  wire  _T_67; // @[NBuffers.scala 34:154:@12141.4]
  wire  _T_69; // @[package.scala 100:49:@12142.4]
  reg  _T_72; // @[package.scala 48:56:@12143.4]
  reg [31:0] _RAND_0;
  SRFF sEn_latch_0 ( // @[NBuffers.scala 21:52:@12050.4]
    .clock(sEn_latch_0_clock),
    .reset(sEn_latch_0_reset),
    .io_input_set(sEn_latch_0_io_input_set),
    .io_input_reset(sEn_latch_0_io_input_reset),
    .io_input_asyn_reset(sEn_latch_0_io_input_asyn_reset),
    .io_output(sEn_latch_0_io_output)
  );
  SRFF sEn_latch_1 ( // @[NBuffers.scala 21:52:@12053.4]
    .clock(sEn_latch_1_clock),
    .reset(sEn_latch_1_reset),
    .io_input_set(sEn_latch_1_io_input_set),
    .io_input_reset(sEn_latch_1_io_input_reset),
    .io_input_asyn_reset(sEn_latch_1_io_input_asyn_reset),
    .io_output(sEn_latch_1_io_output)
  );
  SRFF sDone_latch_0 ( // @[NBuffers.scala 22:54:@12056.4]
    .clock(sDone_latch_0_clock),
    .reset(sDone_latch_0_reset),
    .io_input_set(sDone_latch_0_io_input_set),
    .io_input_reset(sDone_latch_0_io_input_reset),
    .io_input_asyn_reset(sDone_latch_0_io_input_asyn_reset),
    .io_output(sDone_latch_0_io_output)
  );
  SRFF sDone_latch_1 ( // @[NBuffers.scala 22:54:@12059.4]
    .clock(sDone_latch_1_clock),
    .reset(sDone_latch_1_reset),
    .io_input_set(sDone_latch_1_io_input_set),
    .io_input_reset(sDone_latch_1_io_input_reset),
    .io_input_asyn_reset(sDone_latch_1_io_input_asyn_reset),
    .io_output(sDone_latch_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@12066.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@12074.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@12083.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@12091.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@12102.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@12110.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@12119.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@12127.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  NBufCtr NBufCtr ( // @[NBuffers.scala 40:19:@12148.4]
    .clock(NBufCtr_clock),
    .reset(NBufCtr_reset),
    .io_input_countUp(NBufCtr_io_input_countUp),
    .io_input_enable(NBufCtr_io_input_enable),
    .io_output_count(NBufCtr_io_output_count)
  );
  NBufCtr statesInR_0 ( // @[NBuffers.scala 50:19:@12159.4]
    .clock(statesInR_0_clock),
    .reset(statesInR_0_reset),
    .io_input_countUp(statesInR_0_io_input_countUp),
    .io_input_enable(statesInR_0_io_input_enable),
    .io_output_count(statesInR_0_io_output_count)
  );
  NBufCtr_2 statesInR_1 ( // @[NBuffers.scala 50:19:@12170.4]
    .clock(statesInR_1_clock),
    .reset(statesInR_1_reset),
    .io_input_countUp(statesInR_1_io_input_countUp),
    .io_input_enable(statesInR_1_io_input_enable),
    .io_output_count(statesInR_1_io_output_count)
  );
  assign _T_33 = io_sDone_0 == 1'h0; // @[NBuffers.scala 26:46:@12063.4]
  assign _T_48 = io_sDone_1 == 1'h0; // @[NBuffers.scala 26:46:@12099.4]
  assign anyEnabled = sEn_latch_0_io_output | sEn_latch_1_io_output; // @[NBuffers.scala 33:64:@12135.4]
  assign _T_62 = sDone_latch_0_io_output | io_sDone_0; // @[NBuffers.scala 34:124:@12136.4]
  assign _T_63 = sEn_latch_0_io_output == _T_62; // @[NBuffers.scala 34:104:@12137.4]
  assign _T_64 = sDone_latch_1_io_output | io_sDone_1; // @[NBuffers.scala 34:124:@12138.4]
  assign _T_65 = sEn_latch_1_io_output == _T_64; // @[NBuffers.scala 34:104:@12139.4]
  assign _T_66 = _T_63 & _T_65; // @[NBuffers.scala 34:150:@12140.4]
  assign _T_67 = _T_66 & anyEnabled; // @[NBuffers.scala 34:154:@12141.4]
  assign _T_69 = _T_67 == 1'h0; // @[package.scala 100:49:@12142.4]
  assign io_statesInW_0 = NBufCtr_io_output_count[2:0]; // @[NBuffers.scala 44:21:@12158.4]
  assign io_statesInR_1 = statesInR_1_io_output_count[2:0]; // @[NBuffers.scala 54:21:@12180.4]
  assign sEn_latch_0_clock = clock; // @[:@12051.4]
  assign sEn_latch_0_reset = reset; // @[:@12052.4]
  assign sEn_latch_0_io_input_set = io_sEn_0 & _T_33; // @[NBuffers.scala 26:31:@12065.4]
  assign sEn_latch_0_io_input_reset = RetimeWrapper_io_out; // @[NBuffers.scala 27:33:@12073.4]
  assign sEn_latch_0_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[NBuffers.scala 28:38:@12081.4]
  assign sEn_latch_1_clock = clock; // @[:@12054.4]
  assign sEn_latch_1_reset = reset; // @[:@12055.4]
  assign sEn_latch_1_io_input_set = io_sEn_1 & _T_48; // @[NBuffers.scala 26:31:@12101.4]
  assign sEn_latch_1_io_input_reset = RetimeWrapper_4_io_out; // @[NBuffers.scala 27:33:@12109.4]
  assign sEn_latch_1_io_input_asyn_reset = RetimeWrapper_5_io_out; // @[NBuffers.scala 28:38:@12117.4]
  assign sDone_latch_0_clock = clock; // @[:@12057.4]
  assign sDone_latch_0_reset = reset; // @[:@12058.4]
  assign sDone_latch_0_io_input_set = io_sDone_0; // @[NBuffers.scala 29:33:@12082.4]
  assign sDone_latch_0_io_input_reset = RetimeWrapper_2_io_out; // @[NBuffers.scala 30:35:@12090.4]
  assign sDone_latch_0_io_input_asyn_reset = RetimeWrapper_3_io_out; // @[NBuffers.scala 31:40:@12098.4]
  assign sDone_latch_1_clock = clock; // @[:@12060.4]
  assign sDone_latch_1_reset = reset; // @[:@12061.4]
  assign sDone_latch_1_io_input_set = io_sDone_1; // @[NBuffers.scala 29:33:@12118.4]
  assign sDone_latch_1_io_input_reset = RetimeWrapper_6_io_out; // @[NBuffers.scala 30:35:@12126.4]
  assign sDone_latch_1_io_input_asyn_reset = RetimeWrapper_7_io_out; // @[NBuffers.scala 31:40:@12134.4]
  assign RetimeWrapper_clock = clock; // @[:@12067.4]
  assign RetimeWrapper_reset = reset; // @[:@12068.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@12070.4]
  assign RetimeWrapper_io_in = _T_67 & _T_72; // @[package.scala 94:16:@12069.4]
  assign RetimeWrapper_1_clock = clock; // @[:@12075.4]
  assign RetimeWrapper_1_reset = reset; // @[:@12076.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@12078.4]
  assign RetimeWrapper_1_io_in = reset; // @[package.scala 94:16:@12077.4]
  assign RetimeWrapper_2_clock = clock; // @[:@12084.4]
  assign RetimeWrapper_2_reset = reset; // @[:@12085.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@12087.4]
  assign RetimeWrapper_2_io_in = _T_67 & _T_72; // @[package.scala 94:16:@12086.4]
  assign RetimeWrapper_3_clock = clock; // @[:@12092.4]
  assign RetimeWrapper_3_reset = reset; // @[:@12093.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@12095.4]
  assign RetimeWrapper_3_io_in = reset; // @[package.scala 94:16:@12094.4]
  assign RetimeWrapper_4_clock = clock; // @[:@12103.4]
  assign RetimeWrapper_4_reset = reset; // @[:@12104.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@12106.4]
  assign RetimeWrapper_4_io_in = _T_67 & _T_72; // @[package.scala 94:16:@12105.4]
  assign RetimeWrapper_5_clock = clock; // @[:@12111.4]
  assign RetimeWrapper_5_reset = reset; // @[:@12112.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@12114.4]
  assign RetimeWrapper_5_io_in = reset; // @[package.scala 94:16:@12113.4]
  assign RetimeWrapper_6_clock = clock; // @[:@12120.4]
  assign RetimeWrapper_6_reset = reset; // @[:@12121.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@12123.4]
  assign RetimeWrapper_6_io_in = _T_67 & _T_72; // @[package.scala 94:16:@12122.4]
  assign RetimeWrapper_7_clock = clock; // @[:@12128.4]
  assign RetimeWrapper_7_reset = reset; // @[:@12129.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@12131.4]
  assign RetimeWrapper_7_io_in = reset; // @[package.scala 94:16:@12130.4]
  assign NBufCtr_clock = clock; // @[:@12149.4]
  assign NBufCtr_reset = reset; // @[:@12150.4]
  assign NBufCtr_io_input_countUp = 1'h0; // @[NBuffers.scala 43:24:@12157.4]
  assign NBufCtr_io_input_enable = _T_67 & _T_72; // @[NBuffers.scala 42:23:@12156.4]
  assign statesInR_0_clock = clock; // @[:@12160.4]
  assign statesInR_0_reset = reset; // @[:@12161.4]
  assign statesInR_0_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@12168.4]
  assign statesInR_0_io_input_enable = _T_67 & _T_72; // @[NBuffers.scala 52:23:@12167.4]
  assign statesInR_1_clock = clock; // @[:@12171.4]
  assign statesInR_1_reset = reset; // @[:@12172.4]
  assign statesInR_1_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@12179.4]
  assign statesInR_1_io_input_enable = _T_67 & _T_72; // @[NBuffers.scala 52:23:@12178.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_72 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_72 <= 1'h0;
    end else begin
      _T_72 <= _T_69;
    end
  end
endmodule
module NBuf( // @[:@12232.2]
  input         clock, // @[:@12233.4]
  input         reset, // @[:@12234.4]
  output [31:0] io_rPort_0_output_0, // @[:@12235.4]
  input  [31:0] io_wPort_0_data_0, // @[:@12235.4]
  input         io_wPort_0_reset, // @[:@12235.4]
  input         io_wPort_0_en_0, // @[:@12235.4]
  input         io_sEn_0, // @[:@12235.4]
  input         io_sEn_1, // @[:@12235.4]
  input         io_sDone_0, // @[:@12235.4]
  input         io_sDone_1 // @[:@12235.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@12243.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@12243.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@12243.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@12243.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@12243.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@12243.4]
  wire [2:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@12243.4]
  wire [2:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@12243.4]
  wire  FF_clock; // @[NBuffers.scala 146:23:@12250.4]
  wire  FF_reset; // @[NBuffers.scala 146:23:@12250.4]
  wire [31:0] FF_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@12250.4]
  wire [31:0] FF_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@12250.4]
  wire  FF_io_wPort_0_reset; // @[NBuffers.scala 146:23:@12250.4]
  wire  FF_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@12250.4]
  wire  FF_1_clock; // @[NBuffers.scala 146:23:@12266.4]
  wire  FF_1_reset; // @[NBuffers.scala 146:23:@12266.4]
  wire [31:0] FF_1_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@12266.4]
  wire [31:0] FF_1_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@12266.4]
  wire  FF_1_io_wPort_0_reset; // @[NBuffers.scala 146:23:@12266.4]
  wire  FF_1_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@12266.4]
  wire  _T_106; // @[NBuffers.scala 153:105:@12284.4]
  wire  _T_110; // @[NBuffers.scala 157:92:@12294.4]
  wire  _T_113; // @[NBuffers.scala 153:105:@12300.4]
  wire  _T_117; // @[NBuffers.scala 157:92:@12310.4]
  wire [31:0] _T_125; // @[Mux.scala 19:72:@12318.4]
  wire [31:0] _T_127; // @[Mux.scala 19:72:@12319.4]
  NBufController ctrl ( // @[NBuffers.scala 83:20:@12243.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1)
  );
  FF FF ( // @[NBuffers.scala 146:23:@12250.4]
    .clock(FF_clock),
    .reset(FF_reset),
    .io_rPort_0_output_0(FF_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_io_wPort_0_en_0)
  );
  FF FF_1 ( // @[NBuffers.scala 146:23:@12266.4]
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_rPort_0_output_0(FF_1_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_1_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_1_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_1_io_wPort_0_en_0)
  );
  assign _T_106 = ctrl_io_statesInW_0 == 3'h0; // @[NBuffers.scala 153:105:@12284.4]
  assign _T_110 = ctrl_io_statesInR_1 == 3'h0; // @[NBuffers.scala 157:92:@12294.4]
  assign _T_113 = ctrl_io_statesInW_0 == 3'h1; // @[NBuffers.scala 153:105:@12300.4]
  assign _T_117 = ctrl_io_statesInR_1 == 3'h1; // @[NBuffers.scala 157:92:@12310.4]
  assign _T_125 = _T_110 ? FF_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@12318.4]
  assign _T_127 = _T_117 ? FF_1_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@12319.4]
  assign io_rPort_0_output_0 = _T_125 | _T_127; // @[NBuffers.scala 163:66:@12323.4]
  assign ctrl_clock = clock; // @[:@12244.4]
  assign ctrl_reset = reset; // @[:@12245.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@12246.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@12248.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@12247.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@12249.4]
  assign FF_clock = clock; // @[:@12251.4]
  assign FF_reset = reset; // @[:@12252.4]
  assign FF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@12287.4]
  assign FF_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@12288.4]
  assign FF_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_106; // @[MemPrimitives.scala 37:29:@12293.4]
  assign FF_1_clock = clock; // @[:@12267.4]
  assign FF_1_reset = reset; // @[:@12268.4]
  assign FF_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@12303.4]
  assign FF_1_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@12304.4]
  assign FF_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_113; // @[MemPrimitives.scala 37:29:@12309.4]
endmodule
module b542_chain( // @[:@12325.2]
  input         clock, // @[:@12326.4]
  input         reset, // @[:@12327.4]
  output [31:0] io_rPort_0_output_0, // @[:@12328.4]
  input  [31:0] io_wPort_0_data_0, // @[:@12328.4]
  input         io_wPort_0_reset, // @[:@12328.4]
  input         io_wPort_0_en_0, // @[:@12328.4]
  input         io_sEn_0, // @[:@12328.4]
  input         io_sEn_1, // @[:@12328.4]
  input         io_sDone_0, // @[:@12328.4]
  input         io_sDone_1 // @[:@12328.4]
);
  wire  nbufFF_clock; // @[NBuffers.scala 298:22:@12336.4]
  wire  nbufFF_reset; // @[NBuffers.scala 298:22:@12336.4]
  wire [31:0] nbufFF_io_rPort_0_output_0; // @[NBuffers.scala 298:22:@12336.4]
  wire [31:0] nbufFF_io_wPort_0_data_0; // @[NBuffers.scala 298:22:@12336.4]
  wire  nbufFF_io_wPort_0_reset; // @[NBuffers.scala 298:22:@12336.4]
  wire  nbufFF_io_wPort_0_en_0; // @[NBuffers.scala 298:22:@12336.4]
  wire  nbufFF_io_sEn_0; // @[NBuffers.scala 298:22:@12336.4]
  wire  nbufFF_io_sEn_1; // @[NBuffers.scala 298:22:@12336.4]
  wire  nbufFF_io_sDone_0; // @[NBuffers.scala 298:22:@12336.4]
  wire  nbufFF_io_sDone_1; // @[NBuffers.scala 298:22:@12336.4]
  NBuf nbufFF ( // @[NBuffers.scala 298:22:@12336.4]
    .clock(nbufFF_clock),
    .reset(nbufFF_reset),
    .io_rPort_0_output_0(nbufFF_io_rPort_0_output_0),
    .io_wPort_0_data_0(nbufFF_io_wPort_0_data_0),
    .io_wPort_0_reset(nbufFF_io_wPort_0_reset),
    .io_wPort_0_en_0(nbufFF_io_wPort_0_en_0),
    .io_sEn_0(nbufFF_io_sEn_0),
    .io_sEn_1(nbufFF_io_sEn_1),
    .io_sDone_0(nbufFF_io_sDone_0),
    .io_sDone_1(nbufFF_io_sDone_1)
  );
  assign io_rPort_0_output_0 = nbufFF_io_rPort_0_output_0; // @[NBuffers.scala 299:6:@12358.4]
  assign nbufFF_clock = clock; // @[:@12337.4]
  assign nbufFF_reset = reset; // @[:@12338.4]
  assign nbufFF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[NBuffers.scala 299:6:@12355.4]
  assign nbufFF_io_wPort_0_reset = io_wPort_0_reset; // @[NBuffers.scala 299:6:@12354.4]
  assign nbufFF_io_wPort_0_en_0 = io_wPort_0_en_0; // @[NBuffers.scala 299:6:@12351.4]
  assign nbufFF_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 299:6:@12341.4]
  assign nbufFF_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 299:6:@12342.4]
  assign nbufFF_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 299:6:@12339.4]
  assign nbufFF_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 299:6:@12340.4]
endmodule
module FF_9( // @[:@13128.2]
  input   clock, // @[:@13129.4]
  input   reset, // @[:@13130.4]
  output  io_rPort_0_output_0, // @[:@13131.4]
  input   io_wPort_0_data_0, // @[:@13131.4]
  input   io_wPort_0_reset, // @[:@13131.4]
  input   io_wPort_0_en_0 // @[:@13131.4]
);
  reg  ff; // @[MemPrimitives.scala 321:19:@13146.4]
  reg [31:0] _RAND_0;
  wire  _T_68; // @[MemPrimitives.scala 325:32:@13148.4]
  wire  _T_69; // @[MemPrimitives.scala 325:12:@13149.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@13148.4]
  assign _T_69 = io_wPort_0_reset ? 1'h0 : _T_68; // @[MemPrimitives.scala 325:12:@13149.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@13151.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 1'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 1'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module NBuf_1( // @[:@13178.2]
  input   clock, // @[:@13179.4]
  input   reset, // @[:@13180.4]
  output  io_rPort_0_output_0, // @[:@13181.4]
  input   io_wPort_0_data_0, // @[:@13181.4]
  input   io_wPort_0_reset, // @[:@13181.4]
  input   io_wPort_0_en_0, // @[:@13181.4]
  input   io_sEn_0, // @[:@13181.4]
  input   io_sEn_1, // @[:@13181.4]
  input   io_sDone_0, // @[:@13181.4]
  input   io_sDone_1 // @[:@13181.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@13189.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@13189.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@13189.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@13189.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@13189.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@13189.4]
  wire [2:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@13189.4]
  wire [2:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@13189.4]
  wire  FF_clock; // @[NBuffers.scala 146:23:@13196.4]
  wire  FF_reset; // @[NBuffers.scala 146:23:@13196.4]
  wire  FF_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@13196.4]
  wire  FF_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@13196.4]
  wire  FF_io_wPort_0_reset; // @[NBuffers.scala 146:23:@13196.4]
  wire  FF_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@13196.4]
  wire  FF_1_clock; // @[NBuffers.scala 146:23:@13212.4]
  wire  FF_1_reset; // @[NBuffers.scala 146:23:@13212.4]
  wire  FF_1_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@13212.4]
  wire  FF_1_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@13212.4]
  wire  FF_1_io_wPort_0_reset; // @[NBuffers.scala 146:23:@13212.4]
  wire  FF_1_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@13212.4]
  wire  _T_106; // @[NBuffers.scala 153:105:@13230.4]
  wire  _T_110; // @[NBuffers.scala 157:92:@13240.4]
  wire  _T_113; // @[NBuffers.scala 153:105:@13246.4]
  wire  _T_117; // @[NBuffers.scala 157:92:@13256.4]
  wire  _T_125; // @[Mux.scala 19:72:@13264.4]
  wire  _T_127; // @[Mux.scala 19:72:@13265.4]
  NBufController ctrl ( // @[NBuffers.scala 83:20:@13189.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1)
  );
  FF_9 FF ( // @[NBuffers.scala 146:23:@13196.4]
    .clock(FF_clock),
    .reset(FF_reset),
    .io_rPort_0_output_0(FF_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_io_wPort_0_en_0)
  );
  FF_9 FF_1 ( // @[NBuffers.scala 146:23:@13212.4]
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_rPort_0_output_0(FF_1_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_1_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_1_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_1_io_wPort_0_en_0)
  );
  assign _T_106 = ctrl_io_statesInW_0 == 3'h0; // @[NBuffers.scala 153:105:@13230.4]
  assign _T_110 = ctrl_io_statesInR_1 == 3'h0; // @[NBuffers.scala 157:92:@13240.4]
  assign _T_113 = ctrl_io_statesInW_0 == 3'h1; // @[NBuffers.scala 153:105:@13246.4]
  assign _T_117 = ctrl_io_statesInR_1 == 3'h1; // @[NBuffers.scala 157:92:@13256.4]
  assign _T_125 = _T_110 ? FF_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@13264.4]
  assign _T_127 = _T_117 ? FF_1_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@13265.4]
  assign io_rPort_0_output_0 = _T_125 | _T_127; // @[NBuffers.scala 163:66:@13269.4]
  assign ctrl_clock = clock; // @[:@13190.4]
  assign ctrl_reset = reset; // @[:@13191.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@13192.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@13194.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@13193.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@13195.4]
  assign FF_clock = clock; // @[:@13197.4]
  assign FF_reset = reset; // @[:@13198.4]
  assign FF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@13233.4]
  assign FF_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@13234.4]
  assign FF_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_106; // @[MemPrimitives.scala 37:29:@13239.4]
  assign FF_1_clock = clock; // @[:@13213.4]
  assign FF_1_reset = reset; // @[:@13214.4]
  assign FF_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@13249.4]
  assign FF_1_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@13250.4]
  assign FF_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_113; // @[MemPrimitives.scala 37:29:@13255.4]
endmodule
module b543_chain( // @[:@13271.2]
  input   clock, // @[:@13272.4]
  input   reset, // @[:@13273.4]
  output  io_rPort_0_output_0, // @[:@13274.4]
  input   io_wPort_0_data_0, // @[:@13274.4]
  input   io_wPort_0_reset, // @[:@13274.4]
  input   io_wPort_0_en_0, // @[:@13274.4]
  input   io_sEn_0, // @[:@13274.4]
  input   io_sEn_1, // @[:@13274.4]
  input   io_sDone_0, // @[:@13274.4]
  input   io_sDone_1 // @[:@13274.4]
);
  wire  nbufFF_clock; // @[NBuffers.scala 298:22:@13282.4]
  wire  nbufFF_reset; // @[NBuffers.scala 298:22:@13282.4]
  wire  nbufFF_io_rPort_0_output_0; // @[NBuffers.scala 298:22:@13282.4]
  wire  nbufFF_io_wPort_0_data_0; // @[NBuffers.scala 298:22:@13282.4]
  wire  nbufFF_io_wPort_0_reset; // @[NBuffers.scala 298:22:@13282.4]
  wire  nbufFF_io_wPort_0_en_0; // @[NBuffers.scala 298:22:@13282.4]
  wire  nbufFF_io_sEn_0; // @[NBuffers.scala 298:22:@13282.4]
  wire  nbufFF_io_sEn_1; // @[NBuffers.scala 298:22:@13282.4]
  wire  nbufFF_io_sDone_0; // @[NBuffers.scala 298:22:@13282.4]
  wire  nbufFF_io_sDone_1; // @[NBuffers.scala 298:22:@13282.4]
  NBuf_1 nbufFF ( // @[NBuffers.scala 298:22:@13282.4]
    .clock(nbufFF_clock),
    .reset(nbufFF_reset),
    .io_rPort_0_output_0(nbufFF_io_rPort_0_output_0),
    .io_wPort_0_data_0(nbufFF_io_wPort_0_data_0),
    .io_wPort_0_reset(nbufFF_io_wPort_0_reset),
    .io_wPort_0_en_0(nbufFF_io_wPort_0_en_0),
    .io_sEn_0(nbufFF_io_sEn_0),
    .io_sEn_1(nbufFF_io_sEn_1),
    .io_sDone_0(nbufFF_io_sDone_0),
    .io_sDone_1(nbufFF_io_sDone_1)
  );
  assign io_rPort_0_output_0 = nbufFF_io_rPort_0_output_0; // @[NBuffers.scala 299:6:@13304.4]
  assign nbufFF_clock = clock; // @[:@13283.4]
  assign nbufFF_reset = reset; // @[:@13284.4]
  assign nbufFF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[NBuffers.scala 299:6:@13301.4]
  assign nbufFF_io_wPort_0_reset = io_wPort_0_reset; // @[NBuffers.scala 299:6:@13300.4]
  assign nbufFF_io_wPort_0_en_0 = io_wPort_0_en_0; // @[NBuffers.scala 299:6:@13297.4]
  assign nbufFF_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 299:6:@13287.4]
  assign nbufFF_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 299:6:@13288.4]
  assign nbufFF_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 299:6:@13285.4]
  assign nbufFF_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 299:6:@13286.4]
endmodule
module SRAM_4( // @[:@13358.2]
  input         clock, // @[:@13359.4]
  input  [1:0]  io_raddr, // @[:@13361.4]
  input         io_wen, // @[:@13361.4]
  input  [1:0]  io_waddr, // @[:@13361.4]
  input  [31:0] io_wdata, // @[:@13361.4]
  output [31:0] io_rdata, // @[:@13361.4]
  input         io_backpressure // @[:@13361.4]
);
  wire [31:0] SRAMVerilogSim_rdata; // @[SRAM.scala 187:23:@13363.4]
  wire [31:0] SRAMVerilogSim_wdata; // @[SRAM.scala 187:23:@13363.4]
  wire  SRAMVerilogSim_backpressure; // @[SRAM.scala 187:23:@13363.4]
  wire  SRAMVerilogSim_wen; // @[SRAM.scala 187:23:@13363.4]
  wire  SRAMVerilogSim_waddrEn; // @[SRAM.scala 187:23:@13363.4]
  wire  SRAMVerilogSim_raddrEn; // @[SRAM.scala 187:23:@13363.4]
  wire [1:0] SRAMVerilogSim_waddr; // @[SRAM.scala 187:23:@13363.4]
  wire [1:0] SRAMVerilogSim_raddr; // @[SRAM.scala 187:23:@13363.4]
  wire  SRAMVerilogSim_clk; // @[SRAM.scala 187:23:@13363.4]
  SRAMVerilogSim #(.DWIDTH(32), .WORDS(3), .AWIDTH(2)) SRAMVerilogSim ( // @[SRAM.scala 187:23:@13363.4]
    .rdata(SRAMVerilogSim_rdata),
    .wdata(SRAMVerilogSim_wdata),
    .backpressure(SRAMVerilogSim_backpressure),
    .wen(SRAMVerilogSim_wen),
    .waddrEn(SRAMVerilogSim_waddrEn),
    .raddrEn(SRAMVerilogSim_raddrEn),
    .waddr(SRAMVerilogSim_waddr),
    .raddr(SRAMVerilogSim_raddr),
    .clk(SRAMVerilogSim_clk)
  );
  assign io_rdata = SRAMVerilogSim_rdata; // @[SRAM.scala 197:16:@13383.4]
  assign SRAMVerilogSim_wdata = io_wdata; // @[SRAM.scala 192:20:@13377.4]
  assign SRAMVerilogSim_backpressure = io_backpressure; // @[SRAM.scala 193:27:@13378.4]
  assign SRAMVerilogSim_wen = io_wen; // @[SRAM.scala 190:18:@13375.4]
  assign SRAMVerilogSim_waddrEn = 1'h1; // @[SRAM.scala 195:22:@13380.4]
  assign SRAMVerilogSim_raddrEn = 1'h1; // @[SRAM.scala 194:22:@13379.4]
  assign SRAMVerilogSim_waddr = io_waddr; // @[SRAM.scala 191:20:@13376.4]
  assign SRAMVerilogSim_raddr = io_raddr; // @[SRAM.scala 189:20:@13374.4]
  assign SRAMVerilogSim_clk = clock; // @[SRAM.scala 188:18:@13373.4]
endmodule
module RetimeWrapper_113( // @[:@13397.2]
  input        clock, // @[:@13398.4]
  input        reset, // @[:@13399.4]
  input        io_flow, // @[:@13400.4]
  input  [1:0] io_in, // @[:@13400.4]
  output [1:0] io_out // @[:@13400.4]
);
  wire [1:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@13402.4]
  wire [1:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@13402.4]
  wire [1:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@13402.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@13402.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@13402.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@13402.4]
  RetimeShiftRegister #(.WIDTH(2), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@13402.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@13415.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@13414.4]
  assign sr_init = 2'h0; // @[RetimeShiftRegister.scala 19:16:@13413.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@13412.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@13411.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@13409.4]
endmodule
module Mem1D_5( // @[:@13417.2]
  input         clock, // @[:@13418.4]
  input         reset, // @[:@13419.4]
  input  [1:0]  io_r_ofs_0, // @[:@13420.4]
  input         io_r_backpressure, // @[:@13420.4]
  input  [1:0]  io_w_ofs_0, // @[:@13420.4]
  input  [31:0] io_w_data_0, // @[:@13420.4]
  input         io_w_en_0, // @[:@13420.4]
  output [31:0] io_output // @[:@13420.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 753:21:@13424.4]
  wire [1:0] SRAM_io_raddr; // @[MemPrimitives.scala 753:21:@13424.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 753:21:@13424.4]
  wire [1:0] SRAM_io_waddr; // @[MemPrimitives.scala 753:21:@13424.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 753:21:@13424.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 753:21:@13424.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 753:21:@13424.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@13427.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@13427.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@13427.4]
  wire [1:0] RetimeWrapper_io_in; // @[package.scala 93:22:@13427.4]
  wire [1:0] RetimeWrapper_io_out; // @[package.scala 93:22:@13427.4]
  SRAM_4 SRAM ( // @[MemPrimitives.scala 753:21:@13424.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_113 RetimeWrapper ( // @[package.scala 93:22:@13427.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 760:17:@13440.4]
  assign SRAM_clock = clock; // @[:@13425.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 754:37:@13434.4]
  assign SRAM_io_wen = io_w_en_0; // @[MemPrimitives.scala 757:22:@13437.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 756:22:@13435.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 758:22:@13438.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 759:30:@13439.4]
  assign RetimeWrapper_clock = clock; // @[:@13428.4]
  assign RetimeWrapper_reset = reset; // @[:@13429.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@13431.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@13430.4]
endmodule
module x544_accum_0( // @[:@13481.2]
  input         clock, // @[:@13482.4]
  input         reset, // @[:@13483.4]
  input  [1:0]  io_rPort_0_ofs_0, // @[:@13484.4]
  input         io_rPort_0_en_0, // @[:@13484.4]
  output [31:0] io_rPort_0_output_0, // @[:@13484.4]
  input  [1:0]  io_wPort_0_ofs_0, // @[:@13484.4]
  input  [31:0] io_wPort_0_data_0, // @[:@13484.4]
  input         io_wPort_0_en_0 // @[:@13484.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@13499.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@13499.4]
  wire [1:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13499.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13499.4]
  wire [1:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13499.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@13499.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@13499.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@13499.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@13525.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@13525.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@13539.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@13539.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@13539.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@13539.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@13539.4]
  wire [34:0] _T_70; // @[Cat.scala 30:58:@13517.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@13529.4]
  wire [3:0] _T_78; // @[Cat.scala 30:58:@13531.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@13499.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@13525.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@13539.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_70 = {io_wPort_0_en_0,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13517.4]
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@13529.4]
  assign _T_78 = {_T_76,1'h1,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13531.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@13546.4]
  assign Mem1D_clock = clock; // @[:@13500.4]
  assign Mem1D_reset = reset; // @[:@13501.4]
  assign Mem1D_io_r_ofs_0 = _T_78[1:0]; // @[MemPrimitives.scala 131:28:@13535.4]
  assign Mem1D_io_r_backpressure = _T_78[2]; // @[MemPrimitives.scala 132:32:@13536.4]
  assign Mem1D_io_w_ofs_0 = _T_70[1:0]; // @[MemPrimitives.scala 94:28:@13521.4]
  assign Mem1D_io_w_data_0 = _T_70[33:2]; // @[MemPrimitives.scala 95:29:@13522.4]
  assign Mem1D_io_w_en_0 = _T_70[34]; // @[MemPrimitives.scala 96:27:@13523.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@13528.4]
  assign RetimeWrapper_clock = clock; // @[:@13540.4]
  assign RetimeWrapper_reset = reset; // @[:@13541.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@13543.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@13542.4]
endmodule
module x545_accum_1( // @[:@14651.2]
  input         clock, // @[:@14652.4]
  input         reset, // @[:@14653.4]
  input  [1:0]  io_rPort_0_ofs_0, // @[:@14654.4]
  input         io_rPort_0_en_0, // @[:@14654.4]
  output [31:0] io_rPort_0_output_0, // @[:@14654.4]
  input  [1:0]  io_wPort_0_ofs_0, // @[:@14654.4]
  input  [31:0] io_wPort_0_data_0, // @[:@14654.4]
  input         io_wPort_0_en_0, // @[:@14654.4]
  input         io_sEn_0, // @[:@14654.4]
  input         io_sEn_1, // @[:@14654.4]
  input         io_sDone_0, // @[:@14654.4]
  input         io_sDone_1 // @[:@14654.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@14663.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@14663.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@14663.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@14663.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@14663.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@14663.4]
  wire [2:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@14663.4]
  wire [2:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@14663.4]
  wire  SRAM_clock; // @[NBuffers.scala 94:23:@14670.4]
  wire  SRAM_reset; // @[NBuffers.scala 94:23:@14670.4]
  wire [1:0] SRAM_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@14670.4]
  wire  SRAM_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@14670.4]
  wire [31:0] SRAM_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@14670.4]
  wire [1:0] SRAM_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@14670.4]
  wire [31:0] SRAM_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@14670.4]
  wire  SRAM_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@14670.4]
  wire  SRAM_1_clock; // @[NBuffers.scala 94:23:@14686.4]
  wire  SRAM_1_reset; // @[NBuffers.scala 94:23:@14686.4]
  wire [1:0] SRAM_1_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@14686.4]
  wire  SRAM_1_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@14686.4]
  wire [31:0] SRAM_1_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@14686.4]
  wire [1:0] SRAM_1_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@14686.4]
  wire [31:0] SRAM_1_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@14686.4]
  wire  SRAM_1_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@14686.4]
  wire  _T_110; // @[NBuffers.scala 104:105:@14702.4]
  wire  _T_114; // @[NBuffers.scala 108:92:@14712.4]
  wire  _T_117; // @[NBuffers.scala 104:105:@14718.4]
  wire  _T_121; // @[NBuffers.scala 108:92:@14728.4]
  wire [31:0] _T_129; // @[Mux.scala 19:72:@14736.4]
  wire [31:0] _T_131; // @[Mux.scala 19:72:@14737.4]
  NBufController ctrl ( // @[NBuffers.scala 83:20:@14663.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1)
  );
  x544_accum_0 SRAM ( // @[NBuffers.scala 94:23:@14670.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_rPort_0_ofs_0(SRAM_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_io_rPort_0_en_0),
    .io_rPort_0_output_0(SRAM_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(SRAM_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_io_wPort_0_en_0)
  );
  x544_accum_0 SRAM_1 ( // @[NBuffers.scala 94:23:@14686.4]
    .clock(SRAM_1_clock),
    .reset(SRAM_1_reset),
    .io_rPort_0_ofs_0(SRAM_1_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_1_io_rPort_0_en_0),
    .io_rPort_0_output_0(SRAM_1_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(SRAM_1_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_1_io_wPort_0_en_0)
  );
  assign _T_110 = ctrl_io_statesInW_0 == 3'h0; // @[NBuffers.scala 104:105:@14702.4]
  assign _T_114 = ctrl_io_statesInR_1 == 3'h0; // @[NBuffers.scala 108:92:@14712.4]
  assign _T_117 = ctrl_io_statesInW_0 == 3'h1; // @[NBuffers.scala 104:105:@14718.4]
  assign _T_121 = ctrl_io_statesInR_1 == 3'h1; // @[NBuffers.scala 108:92:@14728.4]
  assign _T_129 = _T_114 ? SRAM_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@14736.4]
  assign _T_131 = _T_121 ? SRAM_1_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@14737.4]
  assign io_rPort_0_output_0 = _T_129 | _T_131; // @[NBuffers.scala 115:66:@14741.4]
  assign ctrl_clock = clock; // @[:@14664.4]
  assign ctrl_reset = reset; // @[:@14665.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@14666.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@14668.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@14667.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@14669.4]
  assign SRAM_clock = clock; // @[:@14671.4]
  assign SRAM_reset = reset; // @[:@14672.4]
  assign SRAM_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@14714.4]
  assign SRAM_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_114; // @[MemPrimitives.scala 43:33:@14716.4]
  assign SRAM_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@14704.4]
  assign SRAM_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@14705.4]
  assign SRAM_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_110; // @[MemPrimitives.scala 37:29:@14711.4]
  assign SRAM_1_clock = clock; // @[:@14687.4]
  assign SRAM_1_reset = reset; // @[:@14688.4]
  assign SRAM_1_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@14730.4]
  assign SRAM_1_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_121; // @[MemPrimitives.scala 43:33:@14732.4]
  assign SRAM_1_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@14720.4]
  assign SRAM_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@14721.4]
  assign SRAM_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_117; // @[MemPrimitives.scala 37:29:@14727.4]
endmodule
module FF_12( // @[:@14906.2]
  input        clock, // @[:@14907.4]
  input        reset, // @[:@14908.4]
  output [3:0] io_rPort_0_output_0, // @[:@14909.4]
  input  [3:0] io_wPort_0_data_0, // @[:@14909.4]
  input        io_wPort_0_reset, // @[:@14909.4]
  input        io_wPort_0_en_0 // @[:@14909.4]
);
  reg [3:0] ff; // @[MemPrimitives.scala 321:19:@14924.4]
  reg [31:0] _RAND_0;
  wire [3:0] _T_68; // @[MemPrimitives.scala 325:32:@14926.4]
  wire [3:0] _T_69; // @[MemPrimitives.scala 325:12:@14927.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@14926.4]
  assign _T_69 = io_wPort_0_reset ? 4'h0 : _T_68; // @[MemPrimitives.scala 325:12:@14927.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@14929.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 4'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 4'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_6( // @[:@14944.2]
  input        clock, // @[:@14945.4]
  input        reset, // @[:@14946.4]
  input        io_setup_saturate, // @[:@14947.4]
  input        io_input_reset, // @[:@14947.4]
  input        io_input_enable, // @[:@14947.4]
  output [3:0] io_output_count_0, // @[:@14947.4]
  output       io_output_oobs_0, // @[:@14947.4]
  output       io_output_done // @[:@14947.4]
);
  wire  bases_0_clock; // @[Counter.scala 262:53:@14960.4]
  wire  bases_0_reset; // @[Counter.scala 262:53:@14960.4]
  wire [3:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 262:53:@14960.4]
  wire [3:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 262:53:@14960.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 262:53:@14960.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 262:53:@14960.4]
  wire  SRFF_clock; // @[Counter.scala 264:22:@14976.4]
  wire  SRFF_reset; // @[Counter.scala 264:22:@14976.4]
  wire  SRFF_io_input_set; // @[Counter.scala 264:22:@14976.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 264:22:@14976.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 264:22:@14976.4]
  wire  SRFF_io_output; // @[Counter.scala 264:22:@14976.4]
  wire  _T_36; // @[Counter.scala 265:45:@14979.4]
  wire [3:0] _T_48; // @[Counter.scala 288:52:@15004.4]
  wire [4:0] _T_50; // @[Counter.scala 292:33:@15005.4]
  wire [3:0] _T_51; // @[Counter.scala 292:33:@15006.4]
  wire [3:0] _T_52; // @[Counter.scala 292:33:@15007.4]
  wire  _T_57; // @[Counter.scala 294:18:@15009.4]
  wire [3:0] _T_68; // @[Counter.scala 300:115:@15017.4]
  wire [3:0] _T_70; // @[Counter.scala 300:85:@15019.4]
  wire [3:0] _T_71; // @[Counter.scala 300:152:@15020.4]
  wire [3:0] _T_72; // @[Counter.scala 300:74:@15021.4]
  wire  _T_75; // @[Counter.scala 323:102:@15025.4]
  wire  _T_77; // @[Counter.scala 323:130:@15026.4]
  FF_12 bases_0 ( // @[Counter.scala 262:53:@14960.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 264:22:@14976.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 265:45:@14979.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 288:52:@15004.4]
  assign _T_50 = $signed(_T_48) + $signed(4'sh1); // @[Counter.scala 292:33:@15005.4]
  assign _T_51 = $signed(_T_48) + $signed(4'sh1); // @[Counter.scala 292:33:@15006.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 292:33:@15007.4]
  assign _T_57 = $signed(_T_52) >= $signed(4'sh3); // @[Counter.scala 294:18:@15009.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 300:115:@15017.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 4'h0; // @[Counter.scala 300:85:@15019.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 300:152:@15020.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 300:74:@15021.4]
  assign _T_75 = $signed(_T_48) < $signed(4'sh0); // @[Counter.scala 323:102:@15025.4]
  assign _T_77 = $signed(_T_48) >= $signed(4'sh3); // @[Counter.scala 323:130:@15026.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 305:28:@15024.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 323:60:@15028.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 334:20:@15030.4]
  assign bases_0_clock = clock; // @[:@14961.4]
  assign bases_0_reset = reset; // @[:@14962.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 4'h0 : _T_72; // @[Counter.scala 300:31:@15023.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 282:27:@15002.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 285:29:@15003.4]
  assign SRFF_clock = clock; // @[:@14977.4]
  assign SRFF_reset = reset; // @[:@14978.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 265:23:@14981.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 266:25:@14983.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 267:30:@14984.4]
endmodule
module x549_ctrchain( // @[:@15035.2]
  input        clock, // @[:@15036.4]
  input        reset, // @[:@15037.4]
  input        io_input_reset, // @[:@15038.4]
  input        io_input_enable, // @[:@15038.4]
  output [3:0] io_output_counts_0, // @[:@15038.4]
  output       io_output_oobs_0, // @[:@15038.4]
  output       io_output_done // @[:@15038.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 514:46:@15040.4]
  wire  ctrs_0_reset; // @[Counter.scala 514:46:@15040.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 514:46:@15040.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 514:46:@15040.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 514:46:@15040.4]
  wire [3:0] ctrs_0_io_output_count_0; // @[Counter.scala 514:46:@15040.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 514:46:@15040.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 514:46:@15040.4]
  reg  wasDone; // @[Counter.scala 543:24:@15049.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 547:69:@15055.4]
  wire  _T_47; // @[Counter.scala 547:80:@15056.4]
  reg  doneLatch; // @[Counter.scala 551:26:@15061.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 552:48:@15062.4]
  wire  _T_55; // @[Counter.scala 552:19:@15063.4]
  SingleCounter_6 ctrs_0 ( // @[Counter.scala 514:46:@15040.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 547:69:@15055.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 547:80:@15056.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 552:48:@15062.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 552:19:@15063.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 558:32:@15065.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 559:30:@15067.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 547:18:@15058.4]
  assign ctrs_0_clock = clock; // @[:@15041.4]
  assign ctrs_0_reset = reset; // @[:@15042.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 531:29:@15048.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 521:24:@15046.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 525:33:@15047.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x653_outr_Reduce_sm( // @[:@15854.2]
  input   clock, // @[:@15855.4]
  input   reset, // @[:@15856.4]
  input   io_enable, // @[:@15857.4]
  output  io_done, // @[:@15857.4]
  input   io_ctrDone, // @[:@15857.4]
  output  io_ctrInc, // @[:@15857.4]
  output  io_ctrRst, // @[:@15857.4]
  input   io_parentAck, // @[:@15857.4]
  input   io_backpressure, // @[:@15857.4]
  input   io_doneIn_0, // @[:@15857.4]
  input   io_doneIn_1, // @[:@15857.4]
  input   io_doneIn_2, // @[:@15857.4]
  input   io_doneIn_3, // @[:@15857.4]
  input   io_doneIn_4, // @[:@15857.4]
  input   io_doneIn_5, // @[:@15857.4]
  input   io_doneIn_6, // @[:@15857.4]
  input   io_maskIn_0, // @[:@15857.4]
  input   io_maskIn_1, // @[:@15857.4]
  input   io_maskIn_2, // @[:@15857.4]
  input   io_maskIn_4, // @[:@15857.4]
  input   io_maskIn_5, // @[:@15857.4]
  output  io_enableOut_0, // @[:@15857.4]
  output  io_enableOut_1, // @[:@15857.4]
  output  io_enableOut_2, // @[:@15857.4]
  output  io_enableOut_3, // @[:@15857.4]
  output  io_enableOut_4, // @[:@15857.4]
  output  io_enableOut_5, // @[:@15857.4]
  output  io_enableOut_6, // @[:@15857.4]
  output  io_childAck_0, // @[:@15857.4]
  output  io_childAck_1, // @[:@15857.4]
  output  io_childAck_2, // @[:@15857.4]
  output  io_childAck_3, // @[:@15857.4]
  output  io_childAck_4, // @[:@15857.4]
  output  io_childAck_5, // @[:@15857.4]
  output  io_childAck_6 // @[:@15857.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@15860.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@15860.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@15860.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@15860.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@15860.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@15860.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@15863.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@15863.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@15863.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@15863.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@15863.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@15863.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@15866.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@15866.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@15866.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@15866.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@15866.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@15866.4]
  wire  active_3_clock; // @[Controllers.scala 76:50:@15869.4]
  wire  active_3_reset; // @[Controllers.scala 76:50:@15869.4]
  wire  active_3_io_input_set; // @[Controllers.scala 76:50:@15869.4]
  wire  active_3_io_input_reset; // @[Controllers.scala 76:50:@15869.4]
  wire  active_3_io_input_asyn_reset; // @[Controllers.scala 76:50:@15869.4]
  wire  active_3_io_output; // @[Controllers.scala 76:50:@15869.4]
  wire  active_4_clock; // @[Controllers.scala 76:50:@15872.4]
  wire  active_4_reset; // @[Controllers.scala 76:50:@15872.4]
  wire  active_4_io_input_set; // @[Controllers.scala 76:50:@15872.4]
  wire  active_4_io_input_reset; // @[Controllers.scala 76:50:@15872.4]
  wire  active_4_io_input_asyn_reset; // @[Controllers.scala 76:50:@15872.4]
  wire  active_4_io_output; // @[Controllers.scala 76:50:@15872.4]
  wire  active_5_clock; // @[Controllers.scala 76:50:@15875.4]
  wire  active_5_reset; // @[Controllers.scala 76:50:@15875.4]
  wire  active_5_io_input_set; // @[Controllers.scala 76:50:@15875.4]
  wire  active_5_io_input_reset; // @[Controllers.scala 76:50:@15875.4]
  wire  active_5_io_input_asyn_reset; // @[Controllers.scala 76:50:@15875.4]
  wire  active_5_io_output; // @[Controllers.scala 76:50:@15875.4]
  wire  active_6_clock; // @[Controllers.scala 76:50:@15878.4]
  wire  active_6_reset; // @[Controllers.scala 76:50:@15878.4]
  wire  active_6_io_input_set; // @[Controllers.scala 76:50:@15878.4]
  wire  active_6_io_input_reset; // @[Controllers.scala 76:50:@15878.4]
  wire  active_6_io_input_asyn_reset; // @[Controllers.scala 76:50:@15878.4]
  wire  active_6_io_output; // @[Controllers.scala 76:50:@15878.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@15881.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@15881.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@15881.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@15881.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@15881.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@15881.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@15884.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@15884.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@15884.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@15884.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@15884.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@15884.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@15887.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@15887.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@15887.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@15887.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@15887.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@15887.4]
  wire  done_3_clock; // @[Controllers.scala 77:48:@15890.4]
  wire  done_3_reset; // @[Controllers.scala 77:48:@15890.4]
  wire  done_3_io_input_set; // @[Controllers.scala 77:48:@15890.4]
  wire  done_3_io_input_reset; // @[Controllers.scala 77:48:@15890.4]
  wire  done_3_io_input_asyn_reset; // @[Controllers.scala 77:48:@15890.4]
  wire  done_3_io_output; // @[Controllers.scala 77:48:@15890.4]
  wire  done_4_clock; // @[Controllers.scala 77:48:@15893.4]
  wire  done_4_reset; // @[Controllers.scala 77:48:@15893.4]
  wire  done_4_io_input_set; // @[Controllers.scala 77:48:@15893.4]
  wire  done_4_io_input_reset; // @[Controllers.scala 77:48:@15893.4]
  wire  done_4_io_input_asyn_reset; // @[Controllers.scala 77:48:@15893.4]
  wire  done_4_io_output; // @[Controllers.scala 77:48:@15893.4]
  wire  done_5_clock; // @[Controllers.scala 77:48:@15896.4]
  wire  done_5_reset; // @[Controllers.scala 77:48:@15896.4]
  wire  done_5_io_input_set; // @[Controllers.scala 77:48:@15896.4]
  wire  done_5_io_input_reset; // @[Controllers.scala 77:48:@15896.4]
  wire  done_5_io_input_asyn_reset; // @[Controllers.scala 77:48:@15896.4]
  wire  done_5_io_output; // @[Controllers.scala 77:48:@15896.4]
  wire  done_6_clock; // @[Controllers.scala 77:48:@15899.4]
  wire  done_6_reset; // @[Controllers.scala 77:48:@15899.4]
  wire  done_6_io_input_set; // @[Controllers.scala 77:48:@15899.4]
  wire  done_6_io_input_reset; // @[Controllers.scala 77:48:@15899.4]
  wire  done_6_io_input_asyn_reset; // @[Controllers.scala 77:48:@15899.4]
  wire  done_6_io_output; // @[Controllers.scala 77:48:@15899.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@15988.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@15988.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@15988.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@15988.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@15988.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@15988.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@15991.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@15991.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@15991.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@15991.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@15991.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@15991.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@15994.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@15994.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@15994.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@15994.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@15994.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@15994.4]
  wire  iterDone_3_clock; // @[Controllers.scala 90:52:@15997.4]
  wire  iterDone_3_reset; // @[Controllers.scala 90:52:@15997.4]
  wire  iterDone_3_io_input_set; // @[Controllers.scala 90:52:@15997.4]
  wire  iterDone_3_io_input_reset; // @[Controllers.scala 90:52:@15997.4]
  wire  iterDone_3_io_input_asyn_reset; // @[Controllers.scala 90:52:@15997.4]
  wire  iterDone_3_io_output; // @[Controllers.scala 90:52:@15997.4]
  wire  iterDone_4_clock; // @[Controllers.scala 90:52:@16000.4]
  wire  iterDone_4_reset; // @[Controllers.scala 90:52:@16000.4]
  wire  iterDone_4_io_input_set; // @[Controllers.scala 90:52:@16000.4]
  wire  iterDone_4_io_input_reset; // @[Controllers.scala 90:52:@16000.4]
  wire  iterDone_4_io_input_asyn_reset; // @[Controllers.scala 90:52:@16000.4]
  wire  iterDone_4_io_output; // @[Controllers.scala 90:52:@16000.4]
  wire  iterDone_5_clock; // @[Controllers.scala 90:52:@16003.4]
  wire  iterDone_5_reset; // @[Controllers.scala 90:52:@16003.4]
  wire  iterDone_5_io_input_set; // @[Controllers.scala 90:52:@16003.4]
  wire  iterDone_5_io_input_reset; // @[Controllers.scala 90:52:@16003.4]
  wire  iterDone_5_io_input_asyn_reset; // @[Controllers.scala 90:52:@16003.4]
  wire  iterDone_5_io_output; // @[Controllers.scala 90:52:@16003.4]
  wire  iterDone_6_clock; // @[Controllers.scala 90:52:@16006.4]
  wire  iterDone_6_reset; // @[Controllers.scala 90:52:@16006.4]
  wire  iterDone_6_io_input_set; // @[Controllers.scala 90:52:@16006.4]
  wire  iterDone_6_io_input_reset; // @[Controllers.scala 90:52:@16006.4]
  wire  iterDone_6_io_input_asyn_reset; // @[Controllers.scala 90:52:@16006.4]
  wire  iterDone_6_io_output; // @[Controllers.scala 90:52:@16006.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@16089.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@16089.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@16089.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@16089.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@16089.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@16102.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@16102.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@16102.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@16102.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@16102.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@16115.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@16115.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@16115.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@16115.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@16115.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@16128.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@16128.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@16128.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@16128.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@16128.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@16141.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@16141.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@16141.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@16141.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@16141.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@16154.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@16154.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@16154.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@16154.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@16154.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@16167.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@16167.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@16167.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@16167.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@16167.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@16198.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@16198.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@16198.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@16198.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@16198.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@16218.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@16218.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@16218.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@16218.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@16218.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@16242.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@16242.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@16242.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@16242.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@16242.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@16266.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@16266.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@16266.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@16266.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@16266.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@16290.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@16290.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@16290.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@16290.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@16290.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@16314.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@16314.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@16314.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@16314.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@16314.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@16338.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@16338.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@16338.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@16338.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@16338.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@16437.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@16437.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@16437.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@16437.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@16437.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@16454.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@16454.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@16454.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@16454.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@16454.4]
  wire  _T_77; // @[Controllers.scala 80:47:@15902.4]
  wire  _T_78; // @[Controllers.scala 80:47:@15903.4]
  wire  _T_79; // @[Controllers.scala 80:47:@15904.4]
  wire  _T_80; // @[Controllers.scala 80:47:@15905.4]
  wire  _T_81; // @[Controllers.scala 80:47:@15906.4]
  wire  allDone; // @[Controllers.scala 80:47:@15907.4]
  wire  _T_253; // @[Controllers.scala 102:95:@16088.4]
  wire  _T_247; // @[Controllers.scala 101:55:@16082.4]
  wire  _T_248; // @[Controllers.scala 101:55:@16083.4]
  wire  _T_249; // @[Controllers.scala 101:55:@16084.4]
  wire  _T_250; // @[Controllers.scala 101:55:@16085.4]
  wire  _T_251; // @[Controllers.scala 101:55:@16086.4]
  wire  _T_252; // @[Controllers.scala 101:55:@16087.4]
  wire  _T_257; // @[package.scala 96:25:@16094.4 package.scala 96:25:@16095.4]
  wire  _T_260; // @[Controllers.scala 102:142:@16097.4]
  wire  _T_261; // @[Controllers.scala 102:138:@16098.4]
  wire  _T_262; // @[Controllers.scala 102:123:@16099.4]
  wire  _T_263; // @[Controllers.scala 102:112:@16100.4]
  wire  _T_264; // @[Controllers.scala 102:95:@16101.4]
  wire  _T_268; // @[package.scala 96:25:@16107.4 package.scala 96:25:@16108.4]
  wire  _T_271; // @[Controllers.scala 102:142:@16110.4]
  wire  _T_272; // @[Controllers.scala 102:138:@16111.4]
  wire  _T_273; // @[Controllers.scala 102:123:@16112.4]
  wire  _T_274; // @[Controllers.scala 102:112:@16113.4]
  wire  _T_330; // @[Controllers.scala 102:164:@16179.4]
  wire  _T_275; // @[Controllers.scala 102:95:@16114.4]
  wire  _T_279; // @[package.scala 96:25:@16120.4 package.scala 96:25:@16121.4]
  wire  _T_282; // @[Controllers.scala 102:142:@16123.4]
  wire  _T_283; // @[Controllers.scala 102:138:@16124.4]
  wire  _T_284; // @[Controllers.scala 102:123:@16125.4]
  wire  _T_285; // @[Controllers.scala 102:112:@16126.4]
  wire  _T_331; // @[Controllers.scala 102:164:@16180.4]
  wire  _T_286; // @[Controllers.scala 102:95:@16127.4]
  wire  _T_290; // @[package.scala 96:25:@16133.4 package.scala 96:25:@16134.4]
  wire  _T_293; // @[Controllers.scala 102:142:@16136.4]
  wire  _T_294; // @[Controllers.scala 102:138:@16137.4]
  wire  _T_295; // @[Controllers.scala 102:123:@16138.4]
  wire  _T_296; // @[Controllers.scala 102:112:@16139.4]
  wire  _T_332; // @[Controllers.scala 102:164:@16181.4]
  wire  _T_297; // @[Controllers.scala 102:95:@16140.4]
  wire  _T_301; // @[package.scala 96:25:@16146.4 package.scala 96:25:@16147.4]
  wire  _T_304; // @[Controllers.scala 102:142:@16149.4]
  wire  _T_305; // @[Controllers.scala 102:138:@16150.4]
  wire  _T_306; // @[Controllers.scala 102:123:@16151.4]
  wire  _T_307; // @[Controllers.scala 102:112:@16152.4]
  wire  _T_333; // @[Controllers.scala 102:164:@16182.4]
  wire  _T_308; // @[Controllers.scala 102:95:@16153.4]
  wire  _T_312; // @[package.scala 96:25:@16159.4 package.scala 96:25:@16160.4]
  wire  _T_315; // @[Controllers.scala 102:142:@16162.4]
  wire  _T_316; // @[Controllers.scala 102:138:@16163.4]
  wire  _T_317; // @[Controllers.scala 102:123:@16164.4]
  wire  _T_318; // @[Controllers.scala 102:112:@16165.4]
  wire  _T_334; // @[Controllers.scala 102:164:@16183.4]
  wire  _T_319; // @[Controllers.scala 102:95:@16166.4]
  wire  _T_323; // @[package.scala 96:25:@16172.4 package.scala 96:25:@16173.4]
  wire  _T_326; // @[Controllers.scala 102:142:@16175.4]
  wire  _T_327; // @[Controllers.scala 102:138:@16176.4]
  wire  _T_328; // @[Controllers.scala 102:123:@16177.4]
  wire  _T_329; // @[Controllers.scala 102:112:@16178.4]
  wire  synchronize; // @[Controllers.scala 102:164:@16184.4]
  wire  _T_337; // @[Controllers.scala 105:33:@16186.4]
  wire  _T_339; // @[Controllers.scala 105:54:@16187.4]
  wire  _T_340; // @[Controllers.scala 105:52:@16188.4]
  wire  _T_346; // @[Controllers.scala 107:51:@16195.4]
  wire  _T_349; // @[Controllers.scala 107:64:@16197.4]
  wire  _T_353; // @[package.scala 96:25:@16203.4 package.scala 96:25:@16204.4]
  wire  _T_357; // @[Controllers.scala 107:89:@16206.4]
  wire  _T_358; // @[Controllers.scala 107:86:@16207.4]
  wire  _T_359; // @[Controllers.scala 107:108:@16208.4]
  wire  _T_374; // @[Controllers.scala 114:49:@16226.4]
  wire  _T_377; // @[Controllers.scala 115:57:@16230.4]
  wire  _T_393; // @[Controllers.scala 114:49:@16250.4]
  wire  _T_396; // @[Controllers.scala 115:57:@16254.4]
  wire  _T_412; // @[Controllers.scala 114:49:@16274.4]
  wire  _T_415; // @[Controllers.scala 115:57:@16278.4]
  wire  _T_431; // @[Controllers.scala 114:49:@16298.4]
  wire  _T_434; // @[Controllers.scala 115:57:@16302.4]
  wire  _T_450; // @[Controllers.scala 114:49:@16322.4]
  wire  _T_453; // @[Controllers.scala 115:57:@16326.4]
  wire  _T_469; // @[Controllers.scala 114:49:@16346.4]
  wire  _T_472; // @[Controllers.scala 115:57:@16350.4]
  wire  _T_488; // @[Controllers.scala 213:68:@16375.4]
  wire  _T_489; // @[Controllers.scala 213:92:@16376.4]
  wire  _T_490; // @[Controllers.scala 213:90:@16377.4]
  wire  _T_491; // @[Controllers.scala 213:115:@16378.4]
  wire  _T_492; // @[Controllers.scala 213:132:@16379.4]
  wire  _T_493; // @[Controllers.scala 213:130:@16380.4]
  wire  _T_494; // @[Controllers.scala 213:156:@16381.4]
  wire  _T_496; // @[Controllers.scala 213:68:@16384.4]
  wire  _T_497; // @[Controllers.scala 213:92:@16385.4]
  wire  _T_498; // @[Controllers.scala 213:90:@16386.4]
  wire  _T_499; // @[Controllers.scala 213:115:@16387.4]
  wire  _T_504; // @[Controllers.scala 213:68:@16392.4]
  wire  _T_505; // @[Controllers.scala 213:92:@16393.4]
  wire  _T_506; // @[Controllers.scala 213:90:@16394.4]
  wire  _T_507; // @[Controllers.scala 213:115:@16395.4]
  wire  _T_512; // @[Controllers.scala 213:68:@16400.4]
  wire  _T_513; // @[Controllers.scala 213:92:@16401.4]
  wire  _T_514; // @[Controllers.scala 213:90:@16402.4]
  wire  _T_520; // @[Controllers.scala 213:68:@16408.4]
  wire  _T_521; // @[Controllers.scala 213:92:@16409.4]
  wire  _T_522; // @[Controllers.scala 213:90:@16410.4]
  wire  _T_523; // @[Controllers.scala 213:115:@16411.4]
  wire  _T_528; // @[Controllers.scala 213:68:@16416.4]
  wire  _T_529; // @[Controllers.scala 213:92:@16417.4]
  wire  _T_530; // @[Controllers.scala 213:90:@16418.4]
  wire  _T_531; // @[Controllers.scala 213:115:@16419.4]
  wire  _T_536; // @[Controllers.scala 213:68:@16424.4]
  wire  _T_537; // @[Controllers.scala 213:92:@16425.4]
  wire  _T_538; // @[Controllers.scala 213:90:@16426.4]
  wire  _T_545; // @[package.scala 100:49:@16432.4]
  reg  _T_548; // @[package.scala 48:56:@16433.4]
  reg [31:0] _RAND_0;
  wire  _T_549; // @[package.scala 100:41:@16435.4]
  reg  _T_562; // @[package.scala 48:56:@16451.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@15860.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@15863.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@15866.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF active_3 ( // @[Controllers.scala 76:50:@15869.4]
    .clock(active_3_clock),
    .reset(active_3_reset),
    .io_input_set(active_3_io_input_set),
    .io_input_reset(active_3_io_input_reset),
    .io_input_asyn_reset(active_3_io_input_asyn_reset),
    .io_output(active_3_io_output)
  );
  SRFF active_4 ( // @[Controllers.scala 76:50:@15872.4]
    .clock(active_4_clock),
    .reset(active_4_reset),
    .io_input_set(active_4_io_input_set),
    .io_input_reset(active_4_io_input_reset),
    .io_input_asyn_reset(active_4_io_input_asyn_reset),
    .io_output(active_4_io_output)
  );
  SRFF active_5 ( // @[Controllers.scala 76:50:@15875.4]
    .clock(active_5_clock),
    .reset(active_5_reset),
    .io_input_set(active_5_io_input_set),
    .io_input_reset(active_5_io_input_reset),
    .io_input_asyn_reset(active_5_io_input_asyn_reset),
    .io_output(active_5_io_output)
  );
  SRFF active_6 ( // @[Controllers.scala 76:50:@15878.4]
    .clock(active_6_clock),
    .reset(active_6_reset),
    .io_input_set(active_6_io_input_set),
    .io_input_reset(active_6_io_input_reset),
    .io_input_asyn_reset(active_6_io_input_asyn_reset),
    .io_output(active_6_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@15881.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@15884.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@15887.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF done_3 ( // @[Controllers.scala 77:48:@15890.4]
    .clock(done_3_clock),
    .reset(done_3_reset),
    .io_input_set(done_3_io_input_set),
    .io_input_reset(done_3_io_input_reset),
    .io_input_asyn_reset(done_3_io_input_asyn_reset),
    .io_output(done_3_io_output)
  );
  SRFF done_4 ( // @[Controllers.scala 77:48:@15893.4]
    .clock(done_4_clock),
    .reset(done_4_reset),
    .io_input_set(done_4_io_input_set),
    .io_input_reset(done_4_io_input_reset),
    .io_input_asyn_reset(done_4_io_input_asyn_reset),
    .io_output(done_4_io_output)
  );
  SRFF done_5 ( // @[Controllers.scala 77:48:@15896.4]
    .clock(done_5_clock),
    .reset(done_5_reset),
    .io_input_set(done_5_io_input_set),
    .io_input_reset(done_5_io_input_reset),
    .io_input_asyn_reset(done_5_io_input_asyn_reset),
    .io_output(done_5_io_output)
  );
  SRFF done_6 ( // @[Controllers.scala 77:48:@15899.4]
    .clock(done_6_clock),
    .reset(done_6_reset),
    .io_input_set(done_6_io_input_set),
    .io_input_reset(done_6_io_input_reset),
    .io_input_asyn_reset(done_6_io_input_asyn_reset),
    .io_output(done_6_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@15988.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@15991.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@15994.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  SRFF iterDone_3 ( // @[Controllers.scala 90:52:@15997.4]
    .clock(iterDone_3_clock),
    .reset(iterDone_3_reset),
    .io_input_set(iterDone_3_io_input_set),
    .io_input_reset(iterDone_3_io_input_reset),
    .io_input_asyn_reset(iterDone_3_io_input_asyn_reset),
    .io_output(iterDone_3_io_output)
  );
  SRFF iterDone_4 ( // @[Controllers.scala 90:52:@16000.4]
    .clock(iterDone_4_clock),
    .reset(iterDone_4_reset),
    .io_input_set(iterDone_4_io_input_set),
    .io_input_reset(iterDone_4_io_input_reset),
    .io_input_asyn_reset(iterDone_4_io_input_asyn_reset),
    .io_output(iterDone_4_io_output)
  );
  SRFF iterDone_5 ( // @[Controllers.scala 90:52:@16003.4]
    .clock(iterDone_5_clock),
    .reset(iterDone_5_reset),
    .io_input_set(iterDone_5_io_input_set),
    .io_input_reset(iterDone_5_io_input_reset),
    .io_input_asyn_reset(iterDone_5_io_input_asyn_reset),
    .io_output(iterDone_5_io_output)
  );
  SRFF iterDone_6 ( // @[Controllers.scala 90:52:@16006.4]
    .clock(iterDone_6_clock),
    .reset(iterDone_6_reset),
    .io_input_set(iterDone_6_io_input_set),
    .io_input_reset(iterDone_6_io_input_reset),
    .io_input_asyn_reset(iterDone_6_io_input_asyn_reset),
    .io_output(iterDone_6_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@16089.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@16102.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@16115.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@16128.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@16141.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@16154.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@16167.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@16198.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@16218.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@16242.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@16266.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 ( // @[package.scala 93:22:@16290.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper RetimeWrapper_12 ( // @[package.scala 93:22:@16314.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 ( // @[package.scala 93:22:@16338.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@16437.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@16454.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@15902.4]
  assign _T_78 = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@15903.4]
  assign _T_79 = _T_78 & done_3_io_output; // @[Controllers.scala 80:47:@15904.4]
  assign _T_80 = _T_79 & done_4_io_output; // @[Controllers.scala 80:47:@15905.4]
  assign _T_81 = _T_80 & done_5_io_output; // @[Controllers.scala 80:47:@15906.4]
  assign allDone = _T_81 & done_6_io_output; // @[Controllers.scala 80:47:@15907.4]
  assign _T_253 = active_0_io_output == iterDone_0_io_output; // @[Controllers.scala 102:95:@16088.4]
  assign _T_247 = iterDone_0_io_output | iterDone_1_io_output; // @[Controllers.scala 101:55:@16082.4]
  assign _T_248 = _T_247 | iterDone_2_io_output; // @[Controllers.scala 101:55:@16083.4]
  assign _T_249 = _T_248 | iterDone_3_io_output; // @[Controllers.scala 101:55:@16084.4]
  assign _T_250 = _T_249 | iterDone_4_io_output; // @[Controllers.scala 101:55:@16085.4]
  assign _T_251 = _T_250 | iterDone_5_io_output; // @[Controllers.scala 101:55:@16086.4]
  assign _T_252 = _T_251 | iterDone_6_io_output; // @[Controllers.scala 101:55:@16087.4]
  assign _T_257 = RetimeWrapper_io_out; // @[package.scala 96:25:@16094.4 package.scala 96:25:@16095.4]
  assign _T_260 = ~ _T_257; // @[Controllers.scala 102:142:@16097.4]
  assign _T_261 = active_0_io_output == _T_260; // @[Controllers.scala 102:138:@16098.4]
  assign _T_262 = _T_252 & _T_261; // @[Controllers.scala 102:123:@16099.4]
  assign _T_263 = _T_253 | _T_262; // @[Controllers.scala 102:112:@16100.4]
  assign _T_264 = active_1_io_output == iterDone_1_io_output; // @[Controllers.scala 102:95:@16101.4]
  assign _T_268 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@16107.4 package.scala 96:25:@16108.4]
  assign _T_271 = ~ _T_268; // @[Controllers.scala 102:142:@16110.4]
  assign _T_272 = active_1_io_output == _T_271; // @[Controllers.scala 102:138:@16111.4]
  assign _T_273 = _T_252 & _T_272; // @[Controllers.scala 102:123:@16112.4]
  assign _T_274 = _T_264 | _T_273; // @[Controllers.scala 102:112:@16113.4]
  assign _T_330 = _T_263 & _T_274; // @[Controllers.scala 102:164:@16179.4]
  assign _T_275 = active_2_io_output == iterDone_2_io_output; // @[Controllers.scala 102:95:@16114.4]
  assign _T_279 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@16120.4 package.scala 96:25:@16121.4]
  assign _T_282 = ~ _T_279; // @[Controllers.scala 102:142:@16123.4]
  assign _T_283 = active_2_io_output == _T_282; // @[Controllers.scala 102:138:@16124.4]
  assign _T_284 = _T_252 & _T_283; // @[Controllers.scala 102:123:@16125.4]
  assign _T_285 = _T_275 | _T_284; // @[Controllers.scala 102:112:@16126.4]
  assign _T_331 = _T_330 & _T_285; // @[Controllers.scala 102:164:@16180.4]
  assign _T_286 = active_3_io_output == iterDone_3_io_output; // @[Controllers.scala 102:95:@16127.4]
  assign _T_290 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@16133.4 package.scala 96:25:@16134.4]
  assign _T_293 = ~ _T_290; // @[Controllers.scala 102:142:@16136.4]
  assign _T_294 = active_3_io_output == _T_293; // @[Controllers.scala 102:138:@16137.4]
  assign _T_295 = _T_252 & _T_294; // @[Controllers.scala 102:123:@16138.4]
  assign _T_296 = _T_286 | _T_295; // @[Controllers.scala 102:112:@16139.4]
  assign _T_332 = _T_331 & _T_296; // @[Controllers.scala 102:164:@16181.4]
  assign _T_297 = active_4_io_output == iterDone_4_io_output; // @[Controllers.scala 102:95:@16140.4]
  assign _T_301 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@16146.4 package.scala 96:25:@16147.4]
  assign _T_304 = ~ _T_301; // @[Controllers.scala 102:142:@16149.4]
  assign _T_305 = active_4_io_output == _T_304; // @[Controllers.scala 102:138:@16150.4]
  assign _T_306 = _T_252 & _T_305; // @[Controllers.scala 102:123:@16151.4]
  assign _T_307 = _T_297 | _T_306; // @[Controllers.scala 102:112:@16152.4]
  assign _T_333 = _T_332 & _T_307; // @[Controllers.scala 102:164:@16182.4]
  assign _T_308 = active_5_io_output == iterDone_5_io_output; // @[Controllers.scala 102:95:@16153.4]
  assign _T_312 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@16159.4 package.scala 96:25:@16160.4]
  assign _T_315 = ~ _T_312; // @[Controllers.scala 102:142:@16162.4]
  assign _T_316 = active_5_io_output == _T_315; // @[Controllers.scala 102:138:@16163.4]
  assign _T_317 = _T_252 & _T_316; // @[Controllers.scala 102:123:@16164.4]
  assign _T_318 = _T_308 | _T_317; // @[Controllers.scala 102:112:@16165.4]
  assign _T_334 = _T_333 & _T_318; // @[Controllers.scala 102:164:@16183.4]
  assign _T_319 = active_6_io_output == iterDone_6_io_output; // @[Controllers.scala 102:95:@16166.4]
  assign _T_323 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@16172.4 package.scala 96:25:@16173.4]
  assign _T_326 = ~ _T_323; // @[Controllers.scala 102:142:@16175.4]
  assign _T_327 = active_6_io_output == _T_326; // @[Controllers.scala 102:138:@16176.4]
  assign _T_328 = _T_252 & _T_327; // @[Controllers.scala 102:123:@16177.4]
  assign _T_329 = _T_319 | _T_328; // @[Controllers.scala 102:112:@16178.4]
  assign synchronize = _T_334 & _T_329; // @[Controllers.scala 102:164:@16184.4]
  assign _T_337 = done_0_io_output == 1'h0; // @[Controllers.scala 105:33:@16186.4]
  assign _T_339 = io_ctrDone == 1'h0; // @[Controllers.scala 105:54:@16187.4]
  assign _T_340 = _T_337 & _T_339; // @[Controllers.scala 105:52:@16188.4]
  assign _T_346 = synchronize == 1'h0; // @[Controllers.scala 107:51:@16195.4]
  assign _T_349 = _T_346 & _T_337; // @[Controllers.scala 107:64:@16197.4]
  assign _T_353 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@16203.4 package.scala 96:25:@16204.4]
  assign _T_357 = _T_353 == 1'h0; // @[Controllers.scala 107:89:@16206.4]
  assign _T_358 = _T_349 & _T_357; // @[Controllers.scala 107:86:@16207.4]
  assign _T_359 = _T_358 & io_enable; // @[Controllers.scala 107:108:@16208.4]
  assign _T_374 = synchronize & active_0_io_output; // @[Controllers.scala 114:49:@16226.4]
  assign _T_377 = done_0_io_output & synchronize; // @[Controllers.scala 115:57:@16230.4]
  assign _T_393 = synchronize & active_1_io_output; // @[Controllers.scala 114:49:@16250.4]
  assign _T_396 = done_1_io_output & synchronize; // @[Controllers.scala 115:57:@16254.4]
  assign _T_412 = synchronize & active_2_io_output; // @[Controllers.scala 114:49:@16274.4]
  assign _T_415 = done_2_io_output & synchronize; // @[Controllers.scala 115:57:@16278.4]
  assign _T_431 = synchronize & active_3_io_output; // @[Controllers.scala 114:49:@16298.4]
  assign _T_434 = done_3_io_output & synchronize; // @[Controllers.scala 115:57:@16302.4]
  assign _T_450 = synchronize & active_4_io_output; // @[Controllers.scala 114:49:@16322.4]
  assign _T_453 = done_4_io_output & synchronize; // @[Controllers.scala 115:57:@16326.4]
  assign _T_469 = synchronize & active_5_io_output; // @[Controllers.scala 114:49:@16346.4]
  assign _T_472 = done_5_io_output & synchronize; // @[Controllers.scala 115:57:@16350.4]
  assign _T_488 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@16375.4]
  assign _T_489 = ~ iterDone_0_io_output; // @[Controllers.scala 213:92:@16376.4]
  assign _T_490 = _T_488 & _T_489; // @[Controllers.scala 213:90:@16377.4]
  assign _T_491 = _T_490 & io_maskIn_0; // @[Controllers.scala 213:115:@16378.4]
  assign _T_492 = ~ allDone; // @[Controllers.scala 213:132:@16379.4]
  assign _T_493 = _T_491 & _T_492; // @[Controllers.scala 213:130:@16380.4]
  assign _T_494 = ~ io_ctrDone; // @[Controllers.scala 213:156:@16381.4]
  assign _T_496 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@16384.4]
  assign _T_497 = ~ iterDone_1_io_output; // @[Controllers.scala 213:92:@16385.4]
  assign _T_498 = _T_496 & _T_497; // @[Controllers.scala 213:90:@16386.4]
  assign _T_499 = _T_498 & io_maskIn_1; // @[Controllers.scala 213:115:@16387.4]
  assign _T_504 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@16392.4]
  assign _T_505 = ~ iterDone_2_io_output; // @[Controllers.scala 213:92:@16393.4]
  assign _T_506 = _T_504 & _T_505; // @[Controllers.scala 213:90:@16394.4]
  assign _T_507 = _T_506 & io_maskIn_2; // @[Controllers.scala 213:115:@16395.4]
  assign _T_512 = io_enable & active_3_io_output; // @[Controllers.scala 213:68:@16400.4]
  assign _T_513 = ~ iterDone_3_io_output; // @[Controllers.scala 213:92:@16401.4]
  assign _T_514 = _T_512 & _T_513; // @[Controllers.scala 213:90:@16402.4]
  assign _T_520 = io_enable & active_4_io_output; // @[Controllers.scala 213:68:@16408.4]
  assign _T_521 = ~ iterDone_4_io_output; // @[Controllers.scala 213:92:@16409.4]
  assign _T_522 = _T_520 & _T_521; // @[Controllers.scala 213:90:@16410.4]
  assign _T_523 = _T_522 & io_maskIn_4; // @[Controllers.scala 213:115:@16411.4]
  assign _T_528 = io_enable & active_5_io_output; // @[Controllers.scala 213:68:@16416.4]
  assign _T_529 = ~ iterDone_5_io_output; // @[Controllers.scala 213:92:@16417.4]
  assign _T_530 = _T_528 & _T_529; // @[Controllers.scala 213:90:@16418.4]
  assign _T_531 = _T_530 & io_maskIn_5; // @[Controllers.scala 213:115:@16419.4]
  assign _T_536 = io_enable & active_6_io_output; // @[Controllers.scala 213:68:@16424.4]
  assign _T_537 = ~ iterDone_6_io_output; // @[Controllers.scala 213:92:@16425.4]
  assign _T_538 = _T_536 & _T_537; // @[Controllers.scala 213:90:@16426.4]
  assign _T_545 = allDone == 1'h0; // @[package.scala 100:49:@16432.4]
  assign _T_549 = allDone & _T_548; // @[package.scala 100:41:@16435.4]
  assign io_done = RetimeWrapper_15_io_out; // @[Controllers.scala 245:13:@16461.4]
  assign io_ctrInc = iterDone_0_io_output & synchronize; // @[Controllers.scala 98:17:@16081.4]
  assign io_ctrRst = RetimeWrapper_14_io_out; // @[Controllers.scala 215:13:@16444.4]
  assign io_enableOut_0 = _T_493 & _T_494; // @[Controllers.scala 213:55:@16383.4]
  assign io_enableOut_1 = _T_499 & _T_492; // @[Controllers.scala 213:55:@16391.4]
  assign io_enableOut_2 = _T_507 & _T_492; // @[Controllers.scala 213:55:@16399.4]
  assign io_enableOut_3 = _T_514 & _T_492; // @[Controllers.scala 213:55:@16407.4]
  assign io_enableOut_4 = _T_523 & _T_492; // @[Controllers.scala 213:55:@16415.4]
  assign io_enableOut_5 = _T_531 & _T_492; // @[Controllers.scala 213:55:@16423.4]
  assign io_enableOut_6 = _T_538 & _T_492; // @[Controllers.scala 213:55:@16431.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@16362.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@16364.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@16366.4]
  assign io_childAck_3 = iterDone_3_io_output; // @[Controllers.scala 212:58:@16368.4]
  assign io_childAck_4 = iterDone_4_io_output; // @[Controllers.scala 212:58:@16370.4]
  assign io_childAck_5 = iterDone_5_io_output; // @[Controllers.scala 212:58:@16372.4]
  assign io_childAck_6 = iterDone_6_io_output; // @[Controllers.scala 212:58:@16374.4]
  assign active_0_clock = clock; // @[:@15861.4]
  assign active_0_reset = reset; // @[:@15862.4]
  assign active_0_io_input_set = _T_340 & io_enable; // @[Controllers.scala 105:30:@16191.4]
  assign active_0_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 106:32:@16194.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@15910.4]
  assign active_1_clock = clock; // @[:@15864.4]
  assign active_1_reset = reset; // @[:@15865.4]
  assign active_1_io_input_set = _T_374 & io_enable; // @[Controllers.scala 114:32:@16229.4]
  assign active_1_io_input_reset = _T_377 | io_parentAck; // @[Controllers.scala 115:34:@16233.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@15911.4]
  assign active_2_clock = clock; // @[:@15867.4]
  assign active_2_reset = reset; // @[:@15868.4]
  assign active_2_io_input_set = _T_393 & io_enable; // @[Controllers.scala 114:32:@16253.4]
  assign active_2_io_input_reset = _T_396 | io_parentAck; // @[Controllers.scala 115:34:@16257.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@15912.4]
  assign active_3_clock = clock; // @[:@15870.4]
  assign active_3_reset = reset; // @[:@15871.4]
  assign active_3_io_input_set = _T_412 & io_enable; // @[Controllers.scala 114:32:@16277.4]
  assign active_3_io_input_reset = _T_415 | io_parentAck; // @[Controllers.scala 115:34:@16281.4]
  assign active_3_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@15913.4]
  assign active_4_clock = clock; // @[:@15873.4]
  assign active_4_reset = reset; // @[:@15874.4]
  assign active_4_io_input_set = _T_431 & io_enable; // @[Controllers.scala 114:32:@16301.4]
  assign active_4_io_input_reset = _T_434 | io_parentAck; // @[Controllers.scala 115:34:@16305.4]
  assign active_4_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@15914.4]
  assign active_5_clock = clock; // @[:@15876.4]
  assign active_5_reset = reset; // @[:@15877.4]
  assign active_5_io_input_set = _T_450 & io_enable; // @[Controllers.scala 114:32:@16325.4]
  assign active_5_io_input_reset = _T_453 | io_parentAck; // @[Controllers.scala 115:34:@16329.4]
  assign active_5_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@15915.4]
  assign active_6_clock = clock; // @[:@15879.4]
  assign active_6_reset = reset; // @[:@15880.4]
  assign active_6_io_input_set = _T_469 & io_enable; // @[Controllers.scala 114:32:@16349.4]
  assign active_6_io_input_reset = _T_472 | io_parentAck; // @[Controllers.scala 115:34:@16353.4]
  assign active_6_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@15916.4]
  assign done_0_clock = clock; // @[:@15882.4]
  assign done_0_reset = reset; // @[:@15883.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 108:28:@16216.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@15932.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@15917.4]
  assign done_1_clock = clock; // @[:@15885.4]
  assign done_1_reset = reset; // @[:@15886.4]
  assign done_1_io_input_set = done_0_io_output & synchronize; // @[Controllers.scala 117:30:@16240.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@15941.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@15918.4]
  assign done_2_clock = clock; // @[:@15888.4]
  assign done_2_reset = reset; // @[:@15889.4]
  assign done_2_io_input_set = done_1_io_output & synchronize; // @[Controllers.scala 117:30:@16264.4]
  assign done_2_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@15950.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@15919.4]
  assign done_3_clock = clock; // @[:@15891.4]
  assign done_3_reset = reset; // @[:@15892.4]
  assign done_3_io_input_set = done_2_io_output & synchronize; // @[Controllers.scala 117:30:@16288.4]
  assign done_3_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@15959.4]
  assign done_3_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@15920.4]
  assign done_4_clock = clock; // @[:@15894.4]
  assign done_4_reset = reset; // @[:@15895.4]
  assign done_4_io_input_set = done_3_io_output & synchronize; // @[Controllers.scala 117:30:@16312.4]
  assign done_4_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@15968.4]
  assign done_4_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@15921.4]
  assign done_5_clock = clock; // @[:@15897.4]
  assign done_5_reset = reset; // @[:@15898.4]
  assign done_5_io_input_set = done_4_io_output & synchronize; // @[Controllers.scala 117:30:@16336.4]
  assign done_5_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@15977.4]
  assign done_5_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@15922.4]
  assign done_6_clock = clock; // @[:@15900.4]
  assign done_6_reset = reset; // @[:@15901.4]
  assign done_6_io_input_set = done_5_io_output & synchronize; // @[Controllers.scala 117:30:@16360.4]
  assign done_6_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@15986.4]
  assign done_6_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@15923.4]
  assign iterDone_0_clock = clock; // @[:@15989.4]
  assign iterDone_0_reset = reset; // @[:@15990.4]
  assign iterDone_0_io_input_set = io_doneIn_0 | _T_359; // @[Controllers.scala 107:32:@16212.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@16024.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@16009.4]
  assign iterDone_1_clock = clock; // @[:@15992.4]
  assign iterDone_1_reset = reset; // @[:@15993.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 116:34:@16235.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@16033.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@16010.4]
  assign iterDone_2_clock = clock; // @[:@15995.4]
  assign iterDone_2_reset = reset; // @[:@15996.4]
  assign iterDone_2_io_input_set = io_doneIn_2; // @[Controllers.scala 116:34:@16259.4]
  assign iterDone_2_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@16042.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@16011.4]
  assign iterDone_3_clock = clock; // @[:@15998.4]
  assign iterDone_3_reset = reset; // @[:@15999.4]
  assign iterDone_3_io_input_set = io_doneIn_3; // @[Controllers.scala 116:34:@16283.4]
  assign iterDone_3_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@16051.4]
  assign iterDone_3_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@16012.4]
  assign iterDone_4_clock = clock; // @[:@16001.4]
  assign iterDone_4_reset = reset; // @[:@16002.4]
  assign iterDone_4_io_input_set = io_doneIn_4; // @[Controllers.scala 116:34:@16307.4]
  assign iterDone_4_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@16060.4]
  assign iterDone_4_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@16013.4]
  assign iterDone_5_clock = clock; // @[:@16004.4]
  assign iterDone_5_reset = reset; // @[:@16005.4]
  assign iterDone_5_io_input_set = io_doneIn_5; // @[Controllers.scala 116:34:@16331.4]
  assign iterDone_5_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@16069.4]
  assign iterDone_5_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@16014.4]
  assign iterDone_6_clock = clock; // @[:@16007.4]
  assign iterDone_6_reset = reset; // @[:@16008.4]
  assign iterDone_6_io_input_set = io_doneIn_6; // @[Controllers.scala 116:34:@16355.4]
  assign iterDone_6_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@16078.4]
  assign iterDone_6_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@16015.4]
  assign RetimeWrapper_clock = clock; // @[:@16090.4]
  assign RetimeWrapper_reset = reset; // @[:@16091.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@16093.4]
  assign RetimeWrapper_io_in = io_maskIn_0; // @[package.scala 94:16:@16092.4]
  assign RetimeWrapper_1_clock = clock; // @[:@16103.4]
  assign RetimeWrapper_1_reset = reset; // @[:@16104.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@16106.4]
  assign RetimeWrapper_1_io_in = io_maskIn_1; // @[package.scala 94:16:@16105.4]
  assign RetimeWrapper_2_clock = clock; // @[:@16116.4]
  assign RetimeWrapper_2_reset = reset; // @[:@16117.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@16119.4]
  assign RetimeWrapper_2_io_in = io_maskIn_2; // @[package.scala 94:16:@16118.4]
  assign RetimeWrapper_3_clock = clock; // @[:@16129.4]
  assign RetimeWrapper_3_reset = reset; // @[:@16130.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@16132.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@16131.4]
  assign RetimeWrapper_4_clock = clock; // @[:@16142.4]
  assign RetimeWrapper_4_reset = reset; // @[:@16143.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@16145.4]
  assign RetimeWrapper_4_io_in = io_maskIn_4; // @[package.scala 94:16:@16144.4]
  assign RetimeWrapper_5_clock = clock; // @[:@16155.4]
  assign RetimeWrapper_5_reset = reset; // @[:@16156.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@16158.4]
  assign RetimeWrapper_5_io_in = io_maskIn_5; // @[package.scala 94:16:@16157.4]
  assign RetimeWrapper_6_clock = clock; // @[:@16168.4]
  assign RetimeWrapper_6_reset = reset; // @[:@16169.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@16171.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@16170.4]
  assign RetimeWrapper_7_clock = clock; // @[:@16199.4]
  assign RetimeWrapper_7_reset = reset; // @[:@16200.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@16202.4]
  assign RetimeWrapper_7_io_in = io_maskIn_0; // @[package.scala 94:16:@16201.4]
  assign RetimeWrapper_8_clock = clock; // @[:@16219.4]
  assign RetimeWrapper_8_reset = reset; // @[:@16220.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@16222.4]
  assign RetimeWrapper_8_io_in = synchronize & iterDone_0_io_output; // @[package.scala 94:16:@16221.4]
  assign RetimeWrapper_9_clock = clock; // @[:@16243.4]
  assign RetimeWrapper_9_reset = reset; // @[:@16244.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@16246.4]
  assign RetimeWrapper_9_io_in = synchronize & iterDone_1_io_output; // @[package.scala 94:16:@16245.4]
  assign RetimeWrapper_10_clock = clock; // @[:@16267.4]
  assign RetimeWrapper_10_reset = reset; // @[:@16268.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@16270.4]
  assign RetimeWrapper_10_io_in = synchronize & iterDone_2_io_output; // @[package.scala 94:16:@16269.4]
  assign RetimeWrapper_11_clock = clock; // @[:@16291.4]
  assign RetimeWrapper_11_reset = reset; // @[:@16292.4]
  assign RetimeWrapper_11_io_flow = 1'h1; // @[package.scala 95:18:@16294.4]
  assign RetimeWrapper_11_io_in = synchronize & iterDone_3_io_output; // @[package.scala 94:16:@16293.4]
  assign RetimeWrapper_12_clock = clock; // @[:@16315.4]
  assign RetimeWrapper_12_reset = reset; // @[:@16316.4]
  assign RetimeWrapper_12_io_flow = 1'h1; // @[package.scala 95:18:@16318.4]
  assign RetimeWrapper_12_io_in = synchronize & iterDone_4_io_output; // @[package.scala 94:16:@16317.4]
  assign RetimeWrapper_13_clock = clock; // @[:@16339.4]
  assign RetimeWrapper_13_reset = reset; // @[:@16340.4]
  assign RetimeWrapper_13_io_flow = 1'h1; // @[package.scala 95:18:@16342.4]
  assign RetimeWrapper_13_io_in = synchronize & iterDone_5_io_output; // @[package.scala 94:16:@16341.4]
  assign RetimeWrapper_14_clock = clock; // @[:@16438.4]
  assign RetimeWrapper_14_reset = reset; // @[:@16439.4]
  assign RetimeWrapper_14_io_flow = 1'h1; // @[package.scala 95:18:@16441.4]
  assign RetimeWrapper_14_io_in = _T_549 | io_parentAck; // @[package.scala 94:16:@16440.4]
  assign RetimeWrapper_15_clock = clock; // @[:@16455.4]
  assign RetimeWrapper_15_reset = reset; // @[:@16456.4]
  assign RetimeWrapper_15_io_flow = io_enable; // @[package.scala 95:18:@16458.4]
  assign RetimeWrapper_15_io_in = allDone & _T_562; // @[package.scala 94:16:@16457.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_548 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_562 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_548 <= 1'h0;
    end else begin
      _T_548 <= _T_545;
    end
    if (reset) begin
      _T_562 <= 1'h0;
    end else begin
      _T_562 <= _T_545;
    end
  end
endmodule
module RetimeWrapper_179( // @[:@17795.2]
  input         clock, // @[:@17796.4]
  input         reset, // @[:@17797.4]
  input         io_flow, // @[:@17798.4]
  input  [31:0] io_in, // @[:@17798.4]
  output [31:0] io_out // @[:@17798.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17800.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17800.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17800.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17800.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17800.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17800.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@17800.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17813.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17812.4]
  assign sr_init = 32'h6; // @[RetimeShiftRegister.scala 19:16:@17811.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17810.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17809.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17807.4]
endmodule
module NBufCtr_9( // @[:@17815.2]
  input         clock, // @[:@17816.4]
  input         reset, // @[:@17817.4]
  input         io_input_countUp, // @[:@17818.4]
  input         io_input_enable, // @[:@17818.4]
  output [31:0] io_output_count // @[:@17818.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@17855.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@17855.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@17855.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@17855.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@17855.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@17860.4 package.scala 96:25:@17861.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@17821.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@17822.4]
  wire  _T_21; // @[Counter.scala 49:55:@17823.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@17824.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@17825.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@17826.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@17827.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@17828.4]
  wire  _T_33; // @[Counter.scala 51:52:@17832.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@17833.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@17834.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@17835.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@17836.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@17837.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@17838.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@17839.4]
  wire  _T_45; // @[Counter.scala 52:70:@17840.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@17842.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@17843.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@17844.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@17845.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@17846.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@17847.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@17850.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@17851.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@17853.4]
  RetimeWrapper_179 RetimeWrapper ( // @[package.scala 93:22:@17855.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@17860.4 package.scala 96:25:@17861.4]
  assign _T_18 = {{1'd0}, _T_66}; // @[Counter.scala 49:32:@17821.4]
  assign _T_19 = _T_18[31:0]; // @[Counter.scala 49:32:@17822.4]
  assign _T_21 = _T_19 >= 32'h7; // @[Counter.scala 49:55:@17823.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@17824.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh7); // @[Counter.scala 49:91:@17825.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh7); // @[Counter.scala 49:91:@17826.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@17827.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@17828.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@17832.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@17833.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@17834.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@17835.4]
  assign _T_39 = _T_33 ? 32'h6 : _T_38; // @[Counter.scala 51:47:@17836.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@17837.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@17838.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@17839.4]
  assign _T_45 = _T_43 >= 32'h7; // @[Counter.scala 52:70:@17840.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@17842.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@17843.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@17844.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@17845.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@17846.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@17847.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@17850.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@17851.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@17853.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@17863.4]
  assign RetimeWrapper_clock = clock; // @[:@17856.4]
  assign RetimeWrapper_reset = reset; // @[:@17857.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@17859.4]
  assign RetimeWrapper_io_in = reset ? 32'h6 : _T_62; // @[package.scala 94:16:@17858.4]
endmodule
module NBufCtr_11( // @[:@17979.2]
  input         clock, // @[:@17980.4]
  input         reset, // @[:@17981.4]
  input         io_input_countUp, // @[:@17982.4]
  input         io_input_enable, // @[:@17982.4]
  output [31:0] io_output_count // @[:@17982.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@18019.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@18019.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@18019.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@18019.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@18019.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@18024.4 package.scala 96:25:@18025.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@17985.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@17986.4]
  wire  _T_21; // @[Counter.scala 49:55:@17987.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@17988.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@17989.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@17990.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@17991.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@17992.4]
  wire  _T_33; // @[Counter.scala 51:52:@17996.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@17997.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@17998.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@17999.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@18000.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@18001.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@18010.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@18011.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@18014.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@18015.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@18017.4]
  RetimeWrapper_179 RetimeWrapper ( // @[package.scala 93:22:@18019.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@18024.4 package.scala 96:25:@18025.4]
  assign _T_18 = _T_66 + 32'h1; // @[Counter.scala 49:32:@17985.4]
  assign _T_19 = _T_66 + 32'h1; // @[Counter.scala 49:32:@17986.4]
  assign _T_21 = _T_19 >= 32'h7; // @[Counter.scala 49:55:@17987.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@17988.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 49:91:@17989.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 49:91:@17990.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@17991.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@17992.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@17996.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@17997.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@17998.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@17999.4]
  assign _T_39 = _T_33 ? 32'h6 : _T_38; // @[Counter.scala 51:47:@18000.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@18001.4]
  assign _T_53 = {{1'd0}, _T_27}; // @[Counter.scala 52:107:@18010.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@18011.4]
  assign _T_58 = _T_21 ? _T_54 : _T_19; // @[Counter.scala 52:45:@18014.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@18015.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@18017.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@18027.4]
  assign RetimeWrapper_clock = clock; // @[:@18020.4]
  assign RetimeWrapper_reset = reset; // @[:@18021.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@18023.4]
  assign RetimeWrapper_io_in = reset ? 32'h6 : _T_62; // @[package.scala 94:16:@18022.4]
endmodule
module NBufCtr_12( // @[:@18061.2]
  input         clock, // @[:@18062.4]
  input         reset, // @[:@18063.4]
  input         io_input_countUp, // @[:@18064.4]
  input         io_input_enable, // @[:@18064.4]
  output [31:0] io_output_count // @[:@18064.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@18101.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@18101.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@18101.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@18101.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@18101.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@18106.4 package.scala 96:25:@18107.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@18067.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@18068.4]
  wire  _T_21; // @[Counter.scala 49:55:@18069.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@18070.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@18071.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@18072.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@18073.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@18074.4]
  wire  _T_33; // @[Counter.scala 51:52:@18078.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@18079.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@18080.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@18081.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@18082.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@18083.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@18084.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@18085.4]
  wire  _T_45; // @[Counter.scala 52:70:@18086.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@18088.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@18089.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@18090.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@18091.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@18092.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@18093.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@18096.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@18097.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@18099.4]
  RetimeWrapper_179 RetimeWrapper ( // @[package.scala 93:22:@18101.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@18106.4 package.scala 96:25:@18107.4]
  assign _T_18 = _T_66 + 32'h2; // @[Counter.scala 49:32:@18067.4]
  assign _T_19 = _T_66 + 32'h2; // @[Counter.scala 49:32:@18068.4]
  assign _T_21 = _T_19 >= 32'h7; // @[Counter.scala 49:55:@18069.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@18070.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 49:91:@18071.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 49:91:@18072.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@18073.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@18074.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@18078.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@18079.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@18080.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@18081.4]
  assign _T_39 = _T_33 ? 32'h6 : _T_38; // @[Counter.scala 51:47:@18082.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@18083.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@18084.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@18085.4]
  assign _T_45 = _T_43 >= 32'h7; // @[Counter.scala 52:70:@18086.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@18088.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@18089.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@18090.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@18091.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@18092.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@18093.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@18096.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@18097.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@18099.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@18109.4]
  assign RetimeWrapper_clock = clock; // @[:@18102.4]
  assign RetimeWrapper_reset = reset; // @[:@18103.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@18105.4]
  assign RetimeWrapper_io_in = reset ? 32'h6 : _T_62; // @[package.scala 94:16:@18104.4]
endmodule
module NBufCtr_13( // @[:@18143.2]
  input         clock, // @[:@18144.4]
  input         reset, // @[:@18145.4]
  input         io_input_countUp, // @[:@18146.4]
  input         io_input_enable, // @[:@18146.4]
  output [31:0] io_output_count // @[:@18146.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@18183.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@18183.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@18183.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@18183.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@18183.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@18188.4 package.scala 96:25:@18189.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@18149.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@18150.4]
  wire  _T_21; // @[Counter.scala 49:55:@18151.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@18152.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@18153.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@18154.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@18155.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@18156.4]
  wire  _T_33; // @[Counter.scala 51:52:@18160.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@18161.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@18162.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@18163.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@18164.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@18165.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@18166.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@18167.4]
  wire  _T_45; // @[Counter.scala 52:70:@18168.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@18170.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@18171.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@18172.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@18173.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@18174.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@18175.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@18178.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@18179.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@18181.4]
  RetimeWrapper_179 RetimeWrapper ( // @[package.scala 93:22:@18183.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@18188.4 package.scala 96:25:@18189.4]
  assign _T_18 = _T_66 + 32'h3; // @[Counter.scala 49:32:@18149.4]
  assign _T_19 = _T_66 + 32'h3; // @[Counter.scala 49:32:@18150.4]
  assign _T_21 = _T_19 >= 32'h7; // @[Counter.scala 49:55:@18151.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@18152.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh4); // @[Counter.scala 49:91:@18153.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh4); // @[Counter.scala 49:91:@18154.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@18155.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@18156.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@18160.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@18161.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@18162.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@18163.4]
  assign _T_39 = _T_33 ? 32'h6 : _T_38; // @[Counter.scala 51:47:@18164.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@18165.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@18166.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@18167.4]
  assign _T_45 = _T_43 >= 32'h7; // @[Counter.scala 52:70:@18168.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@18170.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@18171.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@18172.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@18173.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@18174.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@18175.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@18178.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@18179.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@18181.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@18191.4]
  assign RetimeWrapper_clock = clock; // @[:@18184.4]
  assign RetimeWrapper_reset = reset; // @[:@18185.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@18187.4]
  assign RetimeWrapper_io_in = reset ? 32'h6 : _T_62; // @[package.scala 94:16:@18186.4]
endmodule
module NBufCtr_14( // @[:@18225.2]
  input         clock, // @[:@18226.4]
  input         reset, // @[:@18227.4]
  input         io_input_countUp, // @[:@18228.4]
  input         io_input_enable, // @[:@18228.4]
  output [31:0] io_output_count // @[:@18228.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@18265.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@18265.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@18265.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@18265.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@18265.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@18270.4 package.scala 96:25:@18271.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@18231.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@18232.4]
  wire  _T_21; // @[Counter.scala 49:55:@18233.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@18234.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@18235.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@18236.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@18237.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@18238.4]
  wire  _T_33; // @[Counter.scala 51:52:@18242.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@18243.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@18244.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@18245.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@18246.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@18247.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@18248.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@18249.4]
  wire  _T_45; // @[Counter.scala 52:70:@18250.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@18252.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@18253.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@18254.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@18255.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@18256.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@18257.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@18260.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@18261.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@18263.4]
  RetimeWrapper_179 RetimeWrapper ( // @[package.scala 93:22:@18265.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@18270.4 package.scala 96:25:@18271.4]
  assign _T_18 = _T_66 + 32'h4; // @[Counter.scala 49:32:@18231.4]
  assign _T_19 = _T_66 + 32'h4; // @[Counter.scala 49:32:@18232.4]
  assign _T_21 = _T_19 >= 32'h7; // @[Counter.scala 49:55:@18233.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@18234.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh3); // @[Counter.scala 49:91:@18235.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh3); // @[Counter.scala 49:91:@18236.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@18237.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@18238.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@18242.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@18243.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@18244.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@18245.4]
  assign _T_39 = _T_33 ? 32'h6 : _T_38; // @[Counter.scala 51:47:@18246.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@18247.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@18248.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@18249.4]
  assign _T_45 = _T_43 >= 32'h7; // @[Counter.scala 52:70:@18250.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@18252.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@18253.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@18254.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@18255.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@18256.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@18257.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@18260.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@18261.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@18263.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@18273.4]
  assign RetimeWrapper_clock = clock; // @[:@18266.4]
  assign RetimeWrapper_reset = reset; // @[:@18267.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@18269.4]
  assign RetimeWrapper_io_in = reset ? 32'h6 : _T_62; // @[package.scala 94:16:@18268.4]
endmodule
module NBufCtr_15( // @[:@18307.2]
  input         clock, // @[:@18308.4]
  input         reset, // @[:@18309.4]
  input         io_input_countUp, // @[:@18310.4]
  input         io_input_enable, // @[:@18310.4]
  output [31:0] io_output_count // @[:@18310.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@18347.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@18347.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@18347.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@18347.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@18347.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@18352.4 package.scala 96:25:@18353.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@18313.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@18314.4]
  wire  _T_21; // @[Counter.scala 49:55:@18315.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@18316.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@18317.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@18318.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@18319.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@18320.4]
  wire  _T_33; // @[Counter.scala 51:52:@18324.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@18325.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@18326.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@18327.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@18328.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@18329.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@18330.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@18331.4]
  wire  _T_45; // @[Counter.scala 52:70:@18332.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@18334.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@18335.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@18336.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@18337.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@18338.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@18339.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@18342.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@18343.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@18345.4]
  RetimeWrapper_179 RetimeWrapper ( // @[package.scala 93:22:@18347.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@18352.4 package.scala 96:25:@18353.4]
  assign _T_18 = _T_66 + 32'h5; // @[Counter.scala 49:32:@18313.4]
  assign _T_19 = _T_66 + 32'h5; // @[Counter.scala 49:32:@18314.4]
  assign _T_21 = _T_19 >= 32'h7; // @[Counter.scala 49:55:@18315.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@18316.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh2); // @[Counter.scala 49:91:@18317.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh2); // @[Counter.scala 49:91:@18318.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@18319.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@18320.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@18324.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@18325.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@18326.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@18327.4]
  assign _T_39 = _T_33 ? 32'h6 : _T_38; // @[Counter.scala 51:47:@18328.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@18329.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@18330.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@18331.4]
  assign _T_45 = _T_43 >= 32'h7; // @[Counter.scala 52:70:@18332.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@18334.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@18335.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@18336.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@18337.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@18338.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@18339.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@18342.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@18343.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@18345.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@18355.4]
  assign RetimeWrapper_clock = clock; // @[:@18348.4]
  assign RetimeWrapper_reset = reset; // @[:@18349.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@18351.4]
  assign RetimeWrapper_io_in = reset ? 32'h6 : _T_62; // @[package.scala 94:16:@18350.4]
endmodule
module NBufCtr_16( // @[:@18389.2]
  input         clock, // @[:@18390.4]
  input         reset, // @[:@18391.4]
  input         io_input_countUp, // @[:@18392.4]
  input         io_input_enable, // @[:@18392.4]
  output [31:0] io_output_count // @[:@18392.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@18429.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@18429.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@18429.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@18429.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@18429.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@18434.4 package.scala 96:25:@18435.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@18395.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@18396.4]
  wire  _T_21; // @[Counter.scala 49:55:@18397.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@18398.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@18399.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@18400.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@18401.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@18402.4]
  wire  _T_33; // @[Counter.scala 51:52:@18406.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@18407.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@18408.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@18409.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@18410.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@18411.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@18412.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@18413.4]
  wire  _T_45; // @[Counter.scala 52:70:@18414.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@18416.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@18417.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@18418.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@18419.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@18420.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@18421.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@18424.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@18425.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@18427.4]
  RetimeWrapper_179 RetimeWrapper ( // @[package.scala 93:22:@18429.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@18434.4 package.scala 96:25:@18435.4]
  assign _T_18 = _T_66 + 32'h6; // @[Counter.scala 49:32:@18395.4]
  assign _T_19 = _T_66 + 32'h6; // @[Counter.scala 49:32:@18396.4]
  assign _T_21 = _T_19 >= 32'h7; // @[Counter.scala 49:55:@18397.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@18398.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 49:91:@18399.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 49:91:@18400.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@18401.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@18402.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@18406.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@18407.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@18408.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@18409.4]
  assign _T_39 = _T_33 ? 32'h6 : _T_38; // @[Counter.scala 51:47:@18410.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@18411.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@18412.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@18413.4]
  assign _T_45 = _T_43 >= 32'h7; // @[Counter.scala 52:70:@18414.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@18416.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@18417.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@18418.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@18419.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@18420.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@18421.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@18424.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@18425.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@18427.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@18437.4]
  assign RetimeWrapper_clock = clock; // @[:@18430.4]
  assign RetimeWrapper_reset = reset; // @[:@18431.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@18433.4]
  assign RetimeWrapper_io_in = reset ? 32'h6 : _T_62; // @[package.scala 94:16:@18432.4]
endmodule
module NBufController_3( // @[:@18439.2]
  input        clock, // @[:@18440.4]
  input        reset, // @[:@18441.4]
  input        io_sEn_0, // @[:@18442.4]
  input        io_sEn_1, // @[:@18442.4]
  input        io_sEn_2, // @[:@18442.4]
  input        io_sEn_3, // @[:@18442.4]
  input        io_sEn_4, // @[:@18442.4]
  input        io_sEn_5, // @[:@18442.4]
  input        io_sEn_6, // @[:@18442.4]
  input        io_sDone_0, // @[:@18442.4]
  input        io_sDone_1, // @[:@18442.4]
  input        io_sDone_2, // @[:@18442.4]
  input        io_sDone_3, // @[:@18442.4]
  input        io_sDone_4, // @[:@18442.4]
  input        io_sDone_5, // @[:@18442.4]
  input        io_sDone_6, // @[:@18442.4]
  output [3:0] io_statesInW_0, // @[:@18442.4]
  output [3:0] io_statesInR_1, // @[:@18442.4]
  output [3:0] io_statesInR_2, // @[:@18442.4]
  output [3:0] io_statesInR_3, // @[:@18442.4]
  output [3:0] io_statesInR_4, // @[:@18442.4]
  output [3:0] io_statesInR_5, // @[:@18442.4]
  output [3:0] io_statesInR_6 // @[:@18442.4]
);
  wire  sEn_latch_0_clock; // @[NBuffers.scala 21:52:@18444.4]
  wire  sEn_latch_0_reset; // @[NBuffers.scala 21:52:@18444.4]
  wire  sEn_latch_0_io_input_set; // @[NBuffers.scala 21:52:@18444.4]
  wire  sEn_latch_0_io_input_reset; // @[NBuffers.scala 21:52:@18444.4]
  wire  sEn_latch_0_io_input_asyn_reset; // @[NBuffers.scala 21:52:@18444.4]
  wire  sEn_latch_0_io_output; // @[NBuffers.scala 21:52:@18444.4]
  wire  sEn_latch_1_clock; // @[NBuffers.scala 21:52:@18447.4]
  wire  sEn_latch_1_reset; // @[NBuffers.scala 21:52:@18447.4]
  wire  sEn_latch_1_io_input_set; // @[NBuffers.scala 21:52:@18447.4]
  wire  sEn_latch_1_io_input_reset; // @[NBuffers.scala 21:52:@18447.4]
  wire  sEn_latch_1_io_input_asyn_reset; // @[NBuffers.scala 21:52:@18447.4]
  wire  sEn_latch_1_io_output; // @[NBuffers.scala 21:52:@18447.4]
  wire  sEn_latch_2_clock; // @[NBuffers.scala 21:52:@18450.4]
  wire  sEn_latch_2_reset; // @[NBuffers.scala 21:52:@18450.4]
  wire  sEn_latch_2_io_input_set; // @[NBuffers.scala 21:52:@18450.4]
  wire  sEn_latch_2_io_input_reset; // @[NBuffers.scala 21:52:@18450.4]
  wire  sEn_latch_2_io_input_asyn_reset; // @[NBuffers.scala 21:52:@18450.4]
  wire  sEn_latch_2_io_output; // @[NBuffers.scala 21:52:@18450.4]
  wire  sEn_latch_3_clock; // @[NBuffers.scala 21:52:@18453.4]
  wire  sEn_latch_3_reset; // @[NBuffers.scala 21:52:@18453.4]
  wire  sEn_latch_3_io_input_set; // @[NBuffers.scala 21:52:@18453.4]
  wire  sEn_latch_3_io_input_reset; // @[NBuffers.scala 21:52:@18453.4]
  wire  sEn_latch_3_io_input_asyn_reset; // @[NBuffers.scala 21:52:@18453.4]
  wire  sEn_latch_3_io_output; // @[NBuffers.scala 21:52:@18453.4]
  wire  sEn_latch_4_clock; // @[NBuffers.scala 21:52:@18456.4]
  wire  sEn_latch_4_reset; // @[NBuffers.scala 21:52:@18456.4]
  wire  sEn_latch_4_io_input_set; // @[NBuffers.scala 21:52:@18456.4]
  wire  sEn_latch_4_io_input_reset; // @[NBuffers.scala 21:52:@18456.4]
  wire  sEn_latch_4_io_input_asyn_reset; // @[NBuffers.scala 21:52:@18456.4]
  wire  sEn_latch_4_io_output; // @[NBuffers.scala 21:52:@18456.4]
  wire  sEn_latch_5_clock; // @[NBuffers.scala 21:52:@18459.4]
  wire  sEn_latch_5_reset; // @[NBuffers.scala 21:52:@18459.4]
  wire  sEn_latch_5_io_input_set; // @[NBuffers.scala 21:52:@18459.4]
  wire  sEn_latch_5_io_input_reset; // @[NBuffers.scala 21:52:@18459.4]
  wire  sEn_latch_5_io_input_asyn_reset; // @[NBuffers.scala 21:52:@18459.4]
  wire  sEn_latch_5_io_output; // @[NBuffers.scala 21:52:@18459.4]
  wire  sEn_latch_6_clock; // @[NBuffers.scala 21:52:@18462.4]
  wire  sEn_latch_6_reset; // @[NBuffers.scala 21:52:@18462.4]
  wire  sEn_latch_6_io_input_set; // @[NBuffers.scala 21:52:@18462.4]
  wire  sEn_latch_6_io_input_reset; // @[NBuffers.scala 21:52:@18462.4]
  wire  sEn_latch_6_io_input_asyn_reset; // @[NBuffers.scala 21:52:@18462.4]
  wire  sEn_latch_6_io_output; // @[NBuffers.scala 21:52:@18462.4]
  wire  sDone_latch_0_clock; // @[NBuffers.scala 22:54:@18465.4]
  wire  sDone_latch_0_reset; // @[NBuffers.scala 22:54:@18465.4]
  wire  sDone_latch_0_io_input_set; // @[NBuffers.scala 22:54:@18465.4]
  wire  sDone_latch_0_io_input_reset; // @[NBuffers.scala 22:54:@18465.4]
  wire  sDone_latch_0_io_input_asyn_reset; // @[NBuffers.scala 22:54:@18465.4]
  wire  sDone_latch_0_io_output; // @[NBuffers.scala 22:54:@18465.4]
  wire  sDone_latch_1_clock; // @[NBuffers.scala 22:54:@18468.4]
  wire  sDone_latch_1_reset; // @[NBuffers.scala 22:54:@18468.4]
  wire  sDone_latch_1_io_input_set; // @[NBuffers.scala 22:54:@18468.4]
  wire  sDone_latch_1_io_input_reset; // @[NBuffers.scala 22:54:@18468.4]
  wire  sDone_latch_1_io_input_asyn_reset; // @[NBuffers.scala 22:54:@18468.4]
  wire  sDone_latch_1_io_output; // @[NBuffers.scala 22:54:@18468.4]
  wire  sDone_latch_2_clock; // @[NBuffers.scala 22:54:@18471.4]
  wire  sDone_latch_2_reset; // @[NBuffers.scala 22:54:@18471.4]
  wire  sDone_latch_2_io_input_set; // @[NBuffers.scala 22:54:@18471.4]
  wire  sDone_latch_2_io_input_reset; // @[NBuffers.scala 22:54:@18471.4]
  wire  sDone_latch_2_io_input_asyn_reset; // @[NBuffers.scala 22:54:@18471.4]
  wire  sDone_latch_2_io_output; // @[NBuffers.scala 22:54:@18471.4]
  wire  sDone_latch_3_clock; // @[NBuffers.scala 22:54:@18474.4]
  wire  sDone_latch_3_reset; // @[NBuffers.scala 22:54:@18474.4]
  wire  sDone_latch_3_io_input_set; // @[NBuffers.scala 22:54:@18474.4]
  wire  sDone_latch_3_io_input_reset; // @[NBuffers.scala 22:54:@18474.4]
  wire  sDone_latch_3_io_input_asyn_reset; // @[NBuffers.scala 22:54:@18474.4]
  wire  sDone_latch_3_io_output; // @[NBuffers.scala 22:54:@18474.4]
  wire  sDone_latch_4_clock; // @[NBuffers.scala 22:54:@18477.4]
  wire  sDone_latch_4_reset; // @[NBuffers.scala 22:54:@18477.4]
  wire  sDone_latch_4_io_input_set; // @[NBuffers.scala 22:54:@18477.4]
  wire  sDone_latch_4_io_input_reset; // @[NBuffers.scala 22:54:@18477.4]
  wire  sDone_latch_4_io_input_asyn_reset; // @[NBuffers.scala 22:54:@18477.4]
  wire  sDone_latch_4_io_output; // @[NBuffers.scala 22:54:@18477.4]
  wire  sDone_latch_5_clock; // @[NBuffers.scala 22:54:@18480.4]
  wire  sDone_latch_5_reset; // @[NBuffers.scala 22:54:@18480.4]
  wire  sDone_latch_5_io_input_set; // @[NBuffers.scala 22:54:@18480.4]
  wire  sDone_latch_5_io_input_reset; // @[NBuffers.scala 22:54:@18480.4]
  wire  sDone_latch_5_io_input_asyn_reset; // @[NBuffers.scala 22:54:@18480.4]
  wire  sDone_latch_5_io_output; // @[NBuffers.scala 22:54:@18480.4]
  wire  sDone_latch_6_clock; // @[NBuffers.scala 22:54:@18483.4]
  wire  sDone_latch_6_reset; // @[NBuffers.scala 22:54:@18483.4]
  wire  sDone_latch_6_io_input_set; // @[NBuffers.scala 22:54:@18483.4]
  wire  sDone_latch_6_io_input_reset; // @[NBuffers.scala 22:54:@18483.4]
  wire  sDone_latch_6_io_input_asyn_reset; // @[NBuffers.scala 22:54:@18483.4]
  wire  sDone_latch_6_io_output; // @[NBuffers.scala 22:54:@18483.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@18490.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@18490.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@18490.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@18490.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@18490.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@18498.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@18498.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@18498.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@18498.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@18498.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@18507.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@18507.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@18507.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@18507.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@18507.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@18515.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@18515.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@18515.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@18515.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@18515.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@18526.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@18526.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@18526.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@18526.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@18526.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@18534.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@18534.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@18534.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@18534.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@18534.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@18543.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@18543.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@18543.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@18543.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@18543.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@18551.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@18551.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@18551.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@18551.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@18551.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@18562.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@18562.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@18562.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@18562.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@18562.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@18570.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@18570.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@18570.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@18570.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@18570.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@18579.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@18579.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@18579.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@18579.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@18579.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@18587.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@18587.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@18587.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@18587.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@18587.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@18598.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@18598.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@18598.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@18598.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@18598.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@18606.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@18606.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@18606.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@18606.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@18606.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@18615.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@18615.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@18615.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@18615.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@18615.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@18623.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@18623.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@18623.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@18623.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@18623.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@18634.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@18634.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@18634.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@18634.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@18634.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@18642.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@18642.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@18642.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@18642.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@18642.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@18651.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@18651.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@18651.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@18651.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@18651.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@18659.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@18659.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@18659.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@18659.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@18659.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@18670.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@18670.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@18670.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@18670.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@18670.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@18678.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@18678.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@18678.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@18678.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@18678.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@18687.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@18687.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@18687.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@18687.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@18687.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@18695.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@18695.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@18695.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@18695.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@18695.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@18706.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@18706.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@18706.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@18706.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@18706.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@18714.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@18714.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@18714.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@18714.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@18714.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@18723.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@18723.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@18723.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@18723.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@18723.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@18731.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@18731.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@18731.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@18731.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@18731.4]
  wire  NBufCtr_clock; // @[NBuffers.scala 40:19:@18772.4]
  wire  NBufCtr_reset; // @[NBuffers.scala 40:19:@18772.4]
  wire  NBufCtr_io_input_countUp; // @[NBuffers.scala 40:19:@18772.4]
  wire  NBufCtr_io_input_enable; // @[NBuffers.scala 40:19:@18772.4]
  wire [31:0] NBufCtr_io_output_count; // @[NBuffers.scala 40:19:@18772.4]
  wire  statesInR_0_clock; // @[NBuffers.scala 50:19:@18783.4]
  wire  statesInR_0_reset; // @[NBuffers.scala 50:19:@18783.4]
  wire  statesInR_0_io_input_countUp; // @[NBuffers.scala 50:19:@18783.4]
  wire  statesInR_0_io_input_enable; // @[NBuffers.scala 50:19:@18783.4]
  wire [31:0] statesInR_0_io_output_count; // @[NBuffers.scala 50:19:@18783.4]
  wire  statesInR_1_clock; // @[NBuffers.scala 50:19:@18794.4]
  wire  statesInR_1_reset; // @[NBuffers.scala 50:19:@18794.4]
  wire  statesInR_1_io_input_countUp; // @[NBuffers.scala 50:19:@18794.4]
  wire  statesInR_1_io_input_enable; // @[NBuffers.scala 50:19:@18794.4]
  wire [31:0] statesInR_1_io_output_count; // @[NBuffers.scala 50:19:@18794.4]
  wire  statesInR_2_clock; // @[NBuffers.scala 50:19:@18805.4]
  wire  statesInR_2_reset; // @[NBuffers.scala 50:19:@18805.4]
  wire  statesInR_2_io_input_countUp; // @[NBuffers.scala 50:19:@18805.4]
  wire  statesInR_2_io_input_enable; // @[NBuffers.scala 50:19:@18805.4]
  wire [31:0] statesInR_2_io_output_count; // @[NBuffers.scala 50:19:@18805.4]
  wire  statesInR_3_clock; // @[NBuffers.scala 50:19:@18816.4]
  wire  statesInR_3_reset; // @[NBuffers.scala 50:19:@18816.4]
  wire  statesInR_3_io_input_countUp; // @[NBuffers.scala 50:19:@18816.4]
  wire  statesInR_3_io_input_enable; // @[NBuffers.scala 50:19:@18816.4]
  wire [31:0] statesInR_3_io_output_count; // @[NBuffers.scala 50:19:@18816.4]
  wire  statesInR_4_clock; // @[NBuffers.scala 50:19:@18827.4]
  wire  statesInR_4_reset; // @[NBuffers.scala 50:19:@18827.4]
  wire  statesInR_4_io_input_countUp; // @[NBuffers.scala 50:19:@18827.4]
  wire  statesInR_4_io_input_enable; // @[NBuffers.scala 50:19:@18827.4]
  wire [31:0] statesInR_4_io_output_count; // @[NBuffers.scala 50:19:@18827.4]
  wire  statesInR_5_clock; // @[NBuffers.scala 50:19:@18838.4]
  wire  statesInR_5_reset; // @[NBuffers.scala 50:19:@18838.4]
  wire  statesInR_5_io_input_countUp; // @[NBuffers.scala 50:19:@18838.4]
  wire  statesInR_5_io_input_enable; // @[NBuffers.scala 50:19:@18838.4]
  wire [31:0] statesInR_5_io_output_count; // @[NBuffers.scala 50:19:@18838.4]
  wire  statesInR_6_clock; // @[NBuffers.scala 50:19:@18849.4]
  wire  statesInR_6_reset; // @[NBuffers.scala 50:19:@18849.4]
  wire  statesInR_6_io_input_countUp; // @[NBuffers.scala 50:19:@18849.4]
  wire  statesInR_6_io_input_enable; // @[NBuffers.scala 50:19:@18849.4]
  wire [31:0] statesInR_6_io_output_count; // @[NBuffers.scala 50:19:@18849.4]
  wire  _T_33; // @[NBuffers.scala 26:46:@18487.4]
  wire  _T_48; // @[NBuffers.scala 26:46:@18523.4]
  wire  _T_63; // @[NBuffers.scala 26:46:@18559.4]
  wire  _T_78; // @[NBuffers.scala 26:46:@18595.4]
  wire  _T_93; // @[NBuffers.scala 26:46:@18631.4]
  wire  _T_108; // @[NBuffers.scala 26:46:@18667.4]
  wire  _T_123; // @[NBuffers.scala 26:46:@18703.4]
  wire  _T_137; // @[NBuffers.scala 33:64:@18739.4]
  wire  _T_138; // @[NBuffers.scala 33:64:@18740.4]
  wire  _T_139; // @[NBuffers.scala 33:64:@18741.4]
  wire  _T_140; // @[NBuffers.scala 33:64:@18742.4]
  wire  _T_141; // @[NBuffers.scala 33:64:@18743.4]
  wire  anyEnabled; // @[NBuffers.scala 33:64:@18744.4]
  wire  _T_142; // @[NBuffers.scala 34:124:@18745.4]
  wire  _T_143; // @[NBuffers.scala 34:104:@18746.4]
  wire  _T_144; // @[NBuffers.scala 34:124:@18747.4]
  wire  _T_145; // @[NBuffers.scala 34:104:@18748.4]
  wire  _T_146; // @[NBuffers.scala 34:124:@18749.4]
  wire  _T_147; // @[NBuffers.scala 34:104:@18750.4]
  wire  _T_148; // @[NBuffers.scala 34:124:@18751.4]
  wire  _T_149; // @[NBuffers.scala 34:104:@18752.4]
  wire  _T_150; // @[NBuffers.scala 34:124:@18753.4]
  wire  _T_151; // @[NBuffers.scala 34:104:@18754.4]
  wire  _T_152; // @[NBuffers.scala 34:124:@18755.4]
  wire  _T_153; // @[NBuffers.scala 34:104:@18756.4]
  wire  _T_154; // @[NBuffers.scala 34:124:@18757.4]
  wire  _T_155; // @[NBuffers.scala 34:104:@18758.4]
  wire  _T_156; // @[NBuffers.scala 34:150:@18759.4]
  wire  _T_157; // @[NBuffers.scala 34:150:@18760.4]
  wire  _T_158; // @[NBuffers.scala 34:150:@18761.4]
  wire  _T_159; // @[NBuffers.scala 34:150:@18762.4]
  wire  _T_160; // @[NBuffers.scala 34:150:@18763.4]
  wire  _T_161; // @[NBuffers.scala 34:150:@18764.4]
  wire  _T_162; // @[NBuffers.scala 34:154:@18765.4]
  wire  _T_164; // @[package.scala 100:49:@18766.4]
  reg  _T_167; // @[package.scala 48:56:@18767.4]
  reg [31:0] _RAND_0;
  SRFF sEn_latch_0 ( // @[NBuffers.scala 21:52:@18444.4]
    .clock(sEn_latch_0_clock),
    .reset(sEn_latch_0_reset),
    .io_input_set(sEn_latch_0_io_input_set),
    .io_input_reset(sEn_latch_0_io_input_reset),
    .io_input_asyn_reset(sEn_latch_0_io_input_asyn_reset),
    .io_output(sEn_latch_0_io_output)
  );
  SRFF sEn_latch_1 ( // @[NBuffers.scala 21:52:@18447.4]
    .clock(sEn_latch_1_clock),
    .reset(sEn_latch_1_reset),
    .io_input_set(sEn_latch_1_io_input_set),
    .io_input_reset(sEn_latch_1_io_input_reset),
    .io_input_asyn_reset(sEn_latch_1_io_input_asyn_reset),
    .io_output(sEn_latch_1_io_output)
  );
  SRFF sEn_latch_2 ( // @[NBuffers.scala 21:52:@18450.4]
    .clock(sEn_latch_2_clock),
    .reset(sEn_latch_2_reset),
    .io_input_set(sEn_latch_2_io_input_set),
    .io_input_reset(sEn_latch_2_io_input_reset),
    .io_input_asyn_reset(sEn_latch_2_io_input_asyn_reset),
    .io_output(sEn_latch_2_io_output)
  );
  SRFF sEn_latch_3 ( // @[NBuffers.scala 21:52:@18453.4]
    .clock(sEn_latch_3_clock),
    .reset(sEn_latch_3_reset),
    .io_input_set(sEn_latch_3_io_input_set),
    .io_input_reset(sEn_latch_3_io_input_reset),
    .io_input_asyn_reset(sEn_latch_3_io_input_asyn_reset),
    .io_output(sEn_latch_3_io_output)
  );
  SRFF sEn_latch_4 ( // @[NBuffers.scala 21:52:@18456.4]
    .clock(sEn_latch_4_clock),
    .reset(sEn_latch_4_reset),
    .io_input_set(sEn_latch_4_io_input_set),
    .io_input_reset(sEn_latch_4_io_input_reset),
    .io_input_asyn_reset(sEn_latch_4_io_input_asyn_reset),
    .io_output(sEn_latch_4_io_output)
  );
  SRFF sEn_latch_5 ( // @[NBuffers.scala 21:52:@18459.4]
    .clock(sEn_latch_5_clock),
    .reset(sEn_latch_5_reset),
    .io_input_set(sEn_latch_5_io_input_set),
    .io_input_reset(sEn_latch_5_io_input_reset),
    .io_input_asyn_reset(sEn_latch_5_io_input_asyn_reset),
    .io_output(sEn_latch_5_io_output)
  );
  SRFF sEn_latch_6 ( // @[NBuffers.scala 21:52:@18462.4]
    .clock(sEn_latch_6_clock),
    .reset(sEn_latch_6_reset),
    .io_input_set(sEn_latch_6_io_input_set),
    .io_input_reset(sEn_latch_6_io_input_reset),
    .io_input_asyn_reset(sEn_latch_6_io_input_asyn_reset),
    .io_output(sEn_latch_6_io_output)
  );
  SRFF sDone_latch_0 ( // @[NBuffers.scala 22:54:@18465.4]
    .clock(sDone_latch_0_clock),
    .reset(sDone_latch_0_reset),
    .io_input_set(sDone_latch_0_io_input_set),
    .io_input_reset(sDone_latch_0_io_input_reset),
    .io_input_asyn_reset(sDone_latch_0_io_input_asyn_reset),
    .io_output(sDone_latch_0_io_output)
  );
  SRFF sDone_latch_1 ( // @[NBuffers.scala 22:54:@18468.4]
    .clock(sDone_latch_1_clock),
    .reset(sDone_latch_1_reset),
    .io_input_set(sDone_latch_1_io_input_set),
    .io_input_reset(sDone_latch_1_io_input_reset),
    .io_input_asyn_reset(sDone_latch_1_io_input_asyn_reset),
    .io_output(sDone_latch_1_io_output)
  );
  SRFF sDone_latch_2 ( // @[NBuffers.scala 22:54:@18471.4]
    .clock(sDone_latch_2_clock),
    .reset(sDone_latch_2_reset),
    .io_input_set(sDone_latch_2_io_input_set),
    .io_input_reset(sDone_latch_2_io_input_reset),
    .io_input_asyn_reset(sDone_latch_2_io_input_asyn_reset),
    .io_output(sDone_latch_2_io_output)
  );
  SRFF sDone_latch_3 ( // @[NBuffers.scala 22:54:@18474.4]
    .clock(sDone_latch_3_clock),
    .reset(sDone_latch_3_reset),
    .io_input_set(sDone_latch_3_io_input_set),
    .io_input_reset(sDone_latch_3_io_input_reset),
    .io_input_asyn_reset(sDone_latch_3_io_input_asyn_reset),
    .io_output(sDone_latch_3_io_output)
  );
  SRFF sDone_latch_4 ( // @[NBuffers.scala 22:54:@18477.4]
    .clock(sDone_latch_4_clock),
    .reset(sDone_latch_4_reset),
    .io_input_set(sDone_latch_4_io_input_set),
    .io_input_reset(sDone_latch_4_io_input_reset),
    .io_input_asyn_reset(sDone_latch_4_io_input_asyn_reset),
    .io_output(sDone_latch_4_io_output)
  );
  SRFF sDone_latch_5 ( // @[NBuffers.scala 22:54:@18480.4]
    .clock(sDone_latch_5_clock),
    .reset(sDone_latch_5_reset),
    .io_input_set(sDone_latch_5_io_input_set),
    .io_input_reset(sDone_latch_5_io_input_reset),
    .io_input_asyn_reset(sDone_latch_5_io_input_asyn_reset),
    .io_output(sDone_latch_5_io_output)
  );
  SRFF sDone_latch_6 ( // @[NBuffers.scala 22:54:@18483.4]
    .clock(sDone_latch_6_clock),
    .reset(sDone_latch_6_reset),
    .io_input_set(sDone_latch_6_io_input_set),
    .io_input_reset(sDone_latch_6_io_input_reset),
    .io_input_asyn_reset(sDone_latch_6_io_input_asyn_reset),
    .io_output(sDone_latch_6_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@18490.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@18498.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@18507.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@18515.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@18526.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@18534.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@18543.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@18551.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@18562.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@18570.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@18579.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 ( // @[package.scala 93:22:@18587.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper RetimeWrapper_12 ( // @[package.scala 93:22:@18598.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 ( // @[package.scala 93:22:@18606.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@18615.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@18623.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 ( // @[package.scala 93:22:@18634.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper RetimeWrapper_17 ( // @[package.scala 93:22:@18642.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 ( // @[package.scala 93:22:@18651.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper RetimeWrapper_19 ( // @[package.scala 93:22:@18659.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper RetimeWrapper_20 ( // @[package.scala 93:22:@18670.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper RetimeWrapper_21 ( // @[package.scala 93:22:@18678.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper RetimeWrapper_22 ( // @[package.scala 93:22:@18687.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper RetimeWrapper_23 ( // @[package.scala 93:22:@18695.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper RetimeWrapper_24 ( // @[package.scala 93:22:@18706.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@18714.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper RetimeWrapper_26 ( // @[package.scala 93:22:@18723.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper RetimeWrapper_27 ( // @[package.scala 93:22:@18731.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  NBufCtr_9 NBufCtr ( // @[NBuffers.scala 40:19:@18772.4]
    .clock(NBufCtr_clock),
    .reset(NBufCtr_reset),
    .io_input_countUp(NBufCtr_io_input_countUp),
    .io_input_enable(NBufCtr_io_input_enable),
    .io_output_count(NBufCtr_io_output_count)
  );
  NBufCtr_9 statesInR_0 ( // @[NBuffers.scala 50:19:@18783.4]
    .clock(statesInR_0_clock),
    .reset(statesInR_0_reset),
    .io_input_countUp(statesInR_0_io_input_countUp),
    .io_input_enable(statesInR_0_io_input_enable),
    .io_output_count(statesInR_0_io_output_count)
  );
  NBufCtr_11 statesInR_1 ( // @[NBuffers.scala 50:19:@18794.4]
    .clock(statesInR_1_clock),
    .reset(statesInR_1_reset),
    .io_input_countUp(statesInR_1_io_input_countUp),
    .io_input_enable(statesInR_1_io_input_enable),
    .io_output_count(statesInR_1_io_output_count)
  );
  NBufCtr_12 statesInR_2 ( // @[NBuffers.scala 50:19:@18805.4]
    .clock(statesInR_2_clock),
    .reset(statesInR_2_reset),
    .io_input_countUp(statesInR_2_io_input_countUp),
    .io_input_enable(statesInR_2_io_input_enable),
    .io_output_count(statesInR_2_io_output_count)
  );
  NBufCtr_13 statesInR_3 ( // @[NBuffers.scala 50:19:@18816.4]
    .clock(statesInR_3_clock),
    .reset(statesInR_3_reset),
    .io_input_countUp(statesInR_3_io_input_countUp),
    .io_input_enable(statesInR_3_io_input_enable),
    .io_output_count(statesInR_3_io_output_count)
  );
  NBufCtr_14 statesInR_4 ( // @[NBuffers.scala 50:19:@18827.4]
    .clock(statesInR_4_clock),
    .reset(statesInR_4_reset),
    .io_input_countUp(statesInR_4_io_input_countUp),
    .io_input_enable(statesInR_4_io_input_enable),
    .io_output_count(statesInR_4_io_output_count)
  );
  NBufCtr_15 statesInR_5 ( // @[NBuffers.scala 50:19:@18838.4]
    .clock(statesInR_5_clock),
    .reset(statesInR_5_reset),
    .io_input_countUp(statesInR_5_io_input_countUp),
    .io_input_enable(statesInR_5_io_input_enable),
    .io_output_count(statesInR_5_io_output_count)
  );
  NBufCtr_16 statesInR_6 ( // @[NBuffers.scala 50:19:@18849.4]
    .clock(statesInR_6_clock),
    .reset(statesInR_6_reset),
    .io_input_countUp(statesInR_6_io_input_countUp),
    .io_input_enable(statesInR_6_io_input_enable),
    .io_output_count(statesInR_6_io_output_count)
  );
  assign _T_33 = io_sDone_0 == 1'h0; // @[NBuffers.scala 26:46:@18487.4]
  assign _T_48 = io_sDone_1 == 1'h0; // @[NBuffers.scala 26:46:@18523.4]
  assign _T_63 = io_sDone_2 == 1'h0; // @[NBuffers.scala 26:46:@18559.4]
  assign _T_78 = io_sDone_3 == 1'h0; // @[NBuffers.scala 26:46:@18595.4]
  assign _T_93 = io_sDone_4 == 1'h0; // @[NBuffers.scala 26:46:@18631.4]
  assign _T_108 = io_sDone_5 == 1'h0; // @[NBuffers.scala 26:46:@18667.4]
  assign _T_123 = io_sDone_6 == 1'h0; // @[NBuffers.scala 26:46:@18703.4]
  assign _T_137 = sEn_latch_0_io_output | sEn_latch_1_io_output; // @[NBuffers.scala 33:64:@18739.4]
  assign _T_138 = _T_137 | sEn_latch_2_io_output; // @[NBuffers.scala 33:64:@18740.4]
  assign _T_139 = _T_138 | sEn_latch_3_io_output; // @[NBuffers.scala 33:64:@18741.4]
  assign _T_140 = _T_139 | sEn_latch_4_io_output; // @[NBuffers.scala 33:64:@18742.4]
  assign _T_141 = _T_140 | sEn_latch_5_io_output; // @[NBuffers.scala 33:64:@18743.4]
  assign anyEnabled = _T_141 | sEn_latch_6_io_output; // @[NBuffers.scala 33:64:@18744.4]
  assign _T_142 = sDone_latch_0_io_output | io_sDone_0; // @[NBuffers.scala 34:124:@18745.4]
  assign _T_143 = sEn_latch_0_io_output == _T_142; // @[NBuffers.scala 34:104:@18746.4]
  assign _T_144 = sDone_latch_1_io_output | io_sDone_1; // @[NBuffers.scala 34:124:@18747.4]
  assign _T_145 = sEn_latch_1_io_output == _T_144; // @[NBuffers.scala 34:104:@18748.4]
  assign _T_146 = sDone_latch_2_io_output | io_sDone_2; // @[NBuffers.scala 34:124:@18749.4]
  assign _T_147 = sEn_latch_2_io_output == _T_146; // @[NBuffers.scala 34:104:@18750.4]
  assign _T_148 = sDone_latch_3_io_output | io_sDone_3; // @[NBuffers.scala 34:124:@18751.4]
  assign _T_149 = sEn_latch_3_io_output == _T_148; // @[NBuffers.scala 34:104:@18752.4]
  assign _T_150 = sDone_latch_4_io_output | io_sDone_4; // @[NBuffers.scala 34:124:@18753.4]
  assign _T_151 = sEn_latch_4_io_output == _T_150; // @[NBuffers.scala 34:104:@18754.4]
  assign _T_152 = sDone_latch_5_io_output | io_sDone_5; // @[NBuffers.scala 34:124:@18755.4]
  assign _T_153 = sEn_latch_5_io_output == _T_152; // @[NBuffers.scala 34:104:@18756.4]
  assign _T_154 = sDone_latch_6_io_output | io_sDone_6; // @[NBuffers.scala 34:124:@18757.4]
  assign _T_155 = sEn_latch_6_io_output == _T_154; // @[NBuffers.scala 34:104:@18758.4]
  assign _T_156 = _T_143 & _T_145; // @[NBuffers.scala 34:150:@18759.4]
  assign _T_157 = _T_156 & _T_147; // @[NBuffers.scala 34:150:@18760.4]
  assign _T_158 = _T_157 & _T_149; // @[NBuffers.scala 34:150:@18761.4]
  assign _T_159 = _T_158 & _T_151; // @[NBuffers.scala 34:150:@18762.4]
  assign _T_160 = _T_159 & _T_153; // @[NBuffers.scala 34:150:@18763.4]
  assign _T_161 = _T_160 & _T_155; // @[NBuffers.scala 34:150:@18764.4]
  assign _T_162 = _T_161 & anyEnabled; // @[NBuffers.scala 34:154:@18765.4]
  assign _T_164 = _T_162 == 1'h0; // @[package.scala 100:49:@18766.4]
  assign io_statesInW_0 = NBufCtr_io_output_count[3:0]; // @[NBuffers.scala 44:21:@18782.4]
  assign io_statesInR_1 = statesInR_1_io_output_count[3:0]; // @[NBuffers.scala 54:21:@18804.4]
  assign io_statesInR_2 = statesInR_2_io_output_count[3:0]; // @[NBuffers.scala 54:21:@18815.4]
  assign io_statesInR_3 = statesInR_3_io_output_count[3:0]; // @[NBuffers.scala 54:21:@18826.4]
  assign io_statesInR_4 = statesInR_4_io_output_count[3:0]; // @[NBuffers.scala 54:21:@18837.4]
  assign io_statesInR_5 = statesInR_5_io_output_count[3:0]; // @[NBuffers.scala 54:21:@18848.4]
  assign io_statesInR_6 = statesInR_6_io_output_count[3:0]; // @[NBuffers.scala 54:21:@18859.4]
  assign sEn_latch_0_clock = clock; // @[:@18445.4]
  assign sEn_latch_0_reset = reset; // @[:@18446.4]
  assign sEn_latch_0_io_input_set = io_sEn_0 & _T_33; // @[NBuffers.scala 26:31:@18489.4]
  assign sEn_latch_0_io_input_reset = RetimeWrapper_io_out; // @[NBuffers.scala 27:33:@18497.4]
  assign sEn_latch_0_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[NBuffers.scala 28:38:@18505.4]
  assign sEn_latch_1_clock = clock; // @[:@18448.4]
  assign sEn_latch_1_reset = reset; // @[:@18449.4]
  assign sEn_latch_1_io_input_set = io_sEn_1 & _T_48; // @[NBuffers.scala 26:31:@18525.4]
  assign sEn_latch_1_io_input_reset = RetimeWrapper_4_io_out; // @[NBuffers.scala 27:33:@18533.4]
  assign sEn_latch_1_io_input_asyn_reset = RetimeWrapper_5_io_out; // @[NBuffers.scala 28:38:@18541.4]
  assign sEn_latch_2_clock = clock; // @[:@18451.4]
  assign sEn_latch_2_reset = reset; // @[:@18452.4]
  assign sEn_latch_2_io_input_set = io_sEn_2 & _T_63; // @[NBuffers.scala 26:31:@18561.4]
  assign sEn_latch_2_io_input_reset = RetimeWrapper_8_io_out; // @[NBuffers.scala 27:33:@18569.4]
  assign sEn_latch_2_io_input_asyn_reset = RetimeWrapper_9_io_out; // @[NBuffers.scala 28:38:@18577.4]
  assign sEn_latch_3_clock = clock; // @[:@18454.4]
  assign sEn_latch_3_reset = reset; // @[:@18455.4]
  assign sEn_latch_3_io_input_set = io_sEn_3 & _T_78; // @[NBuffers.scala 26:31:@18597.4]
  assign sEn_latch_3_io_input_reset = RetimeWrapper_12_io_out; // @[NBuffers.scala 27:33:@18605.4]
  assign sEn_latch_3_io_input_asyn_reset = RetimeWrapper_13_io_out; // @[NBuffers.scala 28:38:@18613.4]
  assign sEn_latch_4_clock = clock; // @[:@18457.4]
  assign sEn_latch_4_reset = reset; // @[:@18458.4]
  assign sEn_latch_4_io_input_set = io_sEn_4 & _T_93; // @[NBuffers.scala 26:31:@18633.4]
  assign sEn_latch_4_io_input_reset = RetimeWrapper_16_io_out; // @[NBuffers.scala 27:33:@18641.4]
  assign sEn_latch_4_io_input_asyn_reset = RetimeWrapper_17_io_out; // @[NBuffers.scala 28:38:@18649.4]
  assign sEn_latch_5_clock = clock; // @[:@18460.4]
  assign sEn_latch_5_reset = reset; // @[:@18461.4]
  assign sEn_latch_5_io_input_set = io_sEn_5 & _T_108; // @[NBuffers.scala 26:31:@18669.4]
  assign sEn_latch_5_io_input_reset = RetimeWrapper_20_io_out; // @[NBuffers.scala 27:33:@18677.4]
  assign sEn_latch_5_io_input_asyn_reset = RetimeWrapper_21_io_out; // @[NBuffers.scala 28:38:@18685.4]
  assign sEn_latch_6_clock = clock; // @[:@18463.4]
  assign sEn_latch_6_reset = reset; // @[:@18464.4]
  assign sEn_latch_6_io_input_set = io_sEn_6 & _T_123; // @[NBuffers.scala 26:31:@18705.4]
  assign sEn_latch_6_io_input_reset = RetimeWrapper_24_io_out; // @[NBuffers.scala 27:33:@18713.4]
  assign sEn_latch_6_io_input_asyn_reset = RetimeWrapper_25_io_out; // @[NBuffers.scala 28:38:@18721.4]
  assign sDone_latch_0_clock = clock; // @[:@18466.4]
  assign sDone_latch_0_reset = reset; // @[:@18467.4]
  assign sDone_latch_0_io_input_set = io_sDone_0; // @[NBuffers.scala 29:33:@18506.4]
  assign sDone_latch_0_io_input_reset = RetimeWrapper_2_io_out; // @[NBuffers.scala 30:35:@18514.4]
  assign sDone_latch_0_io_input_asyn_reset = RetimeWrapper_3_io_out; // @[NBuffers.scala 31:40:@18522.4]
  assign sDone_latch_1_clock = clock; // @[:@18469.4]
  assign sDone_latch_1_reset = reset; // @[:@18470.4]
  assign sDone_latch_1_io_input_set = io_sDone_1; // @[NBuffers.scala 29:33:@18542.4]
  assign sDone_latch_1_io_input_reset = RetimeWrapper_6_io_out; // @[NBuffers.scala 30:35:@18550.4]
  assign sDone_latch_1_io_input_asyn_reset = RetimeWrapper_7_io_out; // @[NBuffers.scala 31:40:@18558.4]
  assign sDone_latch_2_clock = clock; // @[:@18472.4]
  assign sDone_latch_2_reset = reset; // @[:@18473.4]
  assign sDone_latch_2_io_input_set = io_sDone_2; // @[NBuffers.scala 29:33:@18578.4]
  assign sDone_latch_2_io_input_reset = RetimeWrapper_10_io_out; // @[NBuffers.scala 30:35:@18586.4]
  assign sDone_latch_2_io_input_asyn_reset = RetimeWrapper_11_io_out; // @[NBuffers.scala 31:40:@18594.4]
  assign sDone_latch_3_clock = clock; // @[:@18475.4]
  assign sDone_latch_3_reset = reset; // @[:@18476.4]
  assign sDone_latch_3_io_input_set = io_sDone_3; // @[NBuffers.scala 29:33:@18614.4]
  assign sDone_latch_3_io_input_reset = RetimeWrapper_14_io_out; // @[NBuffers.scala 30:35:@18622.4]
  assign sDone_latch_3_io_input_asyn_reset = RetimeWrapper_15_io_out; // @[NBuffers.scala 31:40:@18630.4]
  assign sDone_latch_4_clock = clock; // @[:@18478.4]
  assign sDone_latch_4_reset = reset; // @[:@18479.4]
  assign sDone_latch_4_io_input_set = io_sDone_4; // @[NBuffers.scala 29:33:@18650.4]
  assign sDone_latch_4_io_input_reset = RetimeWrapper_18_io_out; // @[NBuffers.scala 30:35:@18658.4]
  assign sDone_latch_4_io_input_asyn_reset = RetimeWrapper_19_io_out; // @[NBuffers.scala 31:40:@18666.4]
  assign sDone_latch_5_clock = clock; // @[:@18481.4]
  assign sDone_latch_5_reset = reset; // @[:@18482.4]
  assign sDone_latch_5_io_input_set = io_sDone_5; // @[NBuffers.scala 29:33:@18686.4]
  assign sDone_latch_5_io_input_reset = RetimeWrapper_22_io_out; // @[NBuffers.scala 30:35:@18694.4]
  assign sDone_latch_5_io_input_asyn_reset = RetimeWrapper_23_io_out; // @[NBuffers.scala 31:40:@18702.4]
  assign sDone_latch_6_clock = clock; // @[:@18484.4]
  assign sDone_latch_6_reset = reset; // @[:@18485.4]
  assign sDone_latch_6_io_input_set = io_sDone_6; // @[NBuffers.scala 29:33:@18722.4]
  assign sDone_latch_6_io_input_reset = RetimeWrapper_26_io_out; // @[NBuffers.scala 30:35:@18730.4]
  assign sDone_latch_6_io_input_asyn_reset = RetimeWrapper_27_io_out; // @[NBuffers.scala 31:40:@18738.4]
  assign RetimeWrapper_clock = clock; // @[:@18491.4]
  assign RetimeWrapper_reset = reset; // @[:@18492.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@18494.4]
  assign RetimeWrapper_io_in = _T_162 & _T_167; // @[package.scala 94:16:@18493.4]
  assign RetimeWrapper_1_clock = clock; // @[:@18499.4]
  assign RetimeWrapper_1_reset = reset; // @[:@18500.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@18502.4]
  assign RetimeWrapper_1_io_in = reset; // @[package.scala 94:16:@18501.4]
  assign RetimeWrapper_2_clock = clock; // @[:@18508.4]
  assign RetimeWrapper_2_reset = reset; // @[:@18509.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@18511.4]
  assign RetimeWrapper_2_io_in = _T_162 & _T_167; // @[package.scala 94:16:@18510.4]
  assign RetimeWrapper_3_clock = clock; // @[:@18516.4]
  assign RetimeWrapper_3_reset = reset; // @[:@18517.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@18519.4]
  assign RetimeWrapper_3_io_in = reset; // @[package.scala 94:16:@18518.4]
  assign RetimeWrapper_4_clock = clock; // @[:@18527.4]
  assign RetimeWrapper_4_reset = reset; // @[:@18528.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@18530.4]
  assign RetimeWrapper_4_io_in = _T_162 & _T_167; // @[package.scala 94:16:@18529.4]
  assign RetimeWrapper_5_clock = clock; // @[:@18535.4]
  assign RetimeWrapper_5_reset = reset; // @[:@18536.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@18538.4]
  assign RetimeWrapper_5_io_in = reset; // @[package.scala 94:16:@18537.4]
  assign RetimeWrapper_6_clock = clock; // @[:@18544.4]
  assign RetimeWrapper_6_reset = reset; // @[:@18545.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@18547.4]
  assign RetimeWrapper_6_io_in = _T_162 & _T_167; // @[package.scala 94:16:@18546.4]
  assign RetimeWrapper_7_clock = clock; // @[:@18552.4]
  assign RetimeWrapper_7_reset = reset; // @[:@18553.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@18555.4]
  assign RetimeWrapper_7_io_in = reset; // @[package.scala 94:16:@18554.4]
  assign RetimeWrapper_8_clock = clock; // @[:@18563.4]
  assign RetimeWrapper_8_reset = reset; // @[:@18564.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@18566.4]
  assign RetimeWrapper_8_io_in = _T_162 & _T_167; // @[package.scala 94:16:@18565.4]
  assign RetimeWrapper_9_clock = clock; // @[:@18571.4]
  assign RetimeWrapper_9_reset = reset; // @[:@18572.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@18574.4]
  assign RetimeWrapper_9_io_in = reset; // @[package.scala 94:16:@18573.4]
  assign RetimeWrapper_10_clock = clock; // @[:@18580.4]
  assign RetimeWrapper_10_reset = reset; // @[:@18581.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@18583.4]
  assign RetimeWrapper_10_io_in = _T_162 & _T_167; // @[package.scala 94:16:@18582.4]
  assign RetimeWrapper_11_clock = clock; // @[:@18588.4]
  assign RetimeWrapper_11_reset = reset; // @[:@18589.4]
  assign RetimeWrapper_11_io_flow = 1'h1; // @[package.scala 95:18:@18591.4]
  assign RetimeWrapper_11_io_in = reset; // @[package.scala 94:16:@18590.4]
  assign RetimeWrapper_12_clock = clock; // @[:@18599.4]
  assign RetimeWrapper_12_reset = reset; // @[:@18600.4]
  assign RetimeWrapper_12_io_flow = 1'h1; // @[package.scala 95:18:@18602.4]
  assign RetimeWrapper_12_io_in = _T_162 & _T_167; // @[package.scala 94:16:@18601.4]
  assign RetimeWrapper_13_clock = clock; // @[:@18607.4]
  assign RetimeWrapper_13_reset = reset; // @[:@18608.4]
  assign RetimeWrapper_13_io_flow = 1'h1; // @[package.scala 95:18:@18610.4]
  assign RetimeWrapper_13_io_in = reset; // @[package.scala 94:16:@18609.4]
  assign RetimeWrapper_14_clock = clock; // @[:@18616.4]
  assign RetimeWrapper_14_reset = reset; // @[:@18617.4]
  assign RetimeWrapper_14_io_flow = 1'h1; // @[package.scala 95:18:@18619.4]
  assign RetimeWrapper_14_io_in = _T_162 & _T_167; // @[package.scala 94:16:@18618.4]
  assign RetimeWrapper_15_clock = clock; // @[:@18624.4]
  assign RetimeWrapper_15_reset = reset; // @[:@18625.4]
  assign RetimeWrapper_15_io_flow = 1'h1; // @[package.scala 95:18:@18627.4]
  assign RetimeWrapper_15_io_in = reset; // @[package.scala 94:16:@18626.4]
  assign RetimeWrapper_16_clock = clock; // @[:@18635.4]
  assign RetimeWrapper_16_reset = reset; // @[:@18636.4]
  assign RetimeWrapper_16_io_flow = 1'h1; // @[package.scala 95:18:@18638.4]
  assign RetimeWrapper_16_io_in = _T_162 & _T_167; // @[package.scala 94:16:@18637.4]
  assign RetimeWrapper_17_clock = clock; // @[:@18643.4]
  assign RetimeWrapper_17_reset = reset; // @[:@18644.4]
  assign RetimeWrapper_17_io_flow = 1'h1; // @[package.scala 95:18:@18646.4]
  assign RetimeWrapper_17_io_in = reset; // @[package.scala 94:16:@18645.4]
  assign RetimeWrapper_18_clock = clock; // @[:@18652.4]
  assign RetimeWrapper_18_reset = reset; // @[:@18653.4]
  assign RetimeWrapper_18_io_flow = 1'h1; // @[package.scala 95:18:@18655.4]
  assign RetimeWrapper_18_io_in = _T_162 & _T_167; // @[package.scala 94:16:@18654.4]
  assign RetimeWrapper_19_clock = clock; // @[:@18660.4]
  assign RetimeWrapper_19_reset = reset; // @[:@18661.4]
  assign RetimeWrapper_19_io_flow = 1'h1; // @[package.scala 95:18:@18663.4]
  assign RetimeWrapper_19_io_in = reset; // @[package.scala 94:16:@18662.4]
  assign RetimeWrapper_20_clock = clock; // @[:@18671.4]
  assign RetimeWrapper_20_reset = reset; // @[:@18672.4]
  assign RetimeWrapper_20_io_flow = 1'h1; // @[package.scala 95:18:@18674.4]
  assign RetimeWrapper_20_io_in = _T_162 & _T_167; // @[package.scala 94:16:@18673.4]
  assign RetimeWrapper_21_clock = clock; // @[:@18679.4]
  assign RetimeWrapper_21_reset = reset; // @[:@18680.4]
  assign RetimeWrapper_21_io_flow = 1'h1; // @[package.scala 95:18:@18682.4]
  assign RetimeWrapper_21_io_in = reset; // @[package.scala 94:16:@18681.4]
  assign RetimeWrapper_22_clock = clock; // @[:@18688.4]
  assign RetimeWrapper_22_reset = reset; // @[:@18689.4]
  assign RetimeWrapper_22_io_flow = 1'h1; // @[package.scala 95:18:@18691.4]
  assign RetimeWrapper_22_io_in = _T_162 & _T_167; // @[package.scala 94:16:@18690.4]
  assign RetimeWrapper_23_clock = clock; // @[:@18696.4]
  assign RetimeWrapper_23_reset = reset; // @[:@18697.4]
  assign RetimeWrapper_23_io_flow = 1'h1; // @[package.scala 95:18:@18699.4]
  assign RetimeWrapper_23_io_in = reset; // @[package.scala 94:16:@18698.4]
  assign RetimeWrapper_24_clock = clock; // @[:@18707.4]
  assign RetimeWrapper_24_reset = reset; // @[:@18708.4]
  assign RetimeWrapper_24_io_flow = 1'h1; // @[package.scala 95:18:@18710.4]
  assign RetimeWrapper_24_io_in = _T_162 & _T_167; // @[package.scala 94:16:@18709.4]
  assign RetimeWrapper_25_clock = clock; // @[:@18715.4]
  assign RetimeWrapper_25_reset = reset; // @[:@18716.4]
  assign RetimeWrapper_25_io_flow = 1'h1; // @[package.scala 95:18:@18718.4]
  assign RetimeWrapper_25_io_in = reset; // @[package.scala 94:16:@18717.4]
  assign RetimeWrapper_26_clock = clock; // @[:@18724.4]
  assign RetimeWrapper_26_reset = reset; // @[:@18725.4]
  assign RetimeWrapper_26_io_flow = 1'h1; // @[package.scala 95:18:@18727.4]
  assign RetimeWrapper_26_io_in = _T_162 & _T_167; // @[package.scala 94:16:@18726.4]
  assign RetimeWrapper_27_clock = clock; // @[:@18732.4]
  assign RetimeWrapper_27_reset = reset; // @[:@18733.4]
  assign RetimeWrapper_27_io_flow = 1'h1; // @[package.scala 95:18:@18735.4]
  assign RetimeWrapper_27_io_in = reset; // @[package.scala 94:16:@18734.4]
  assign NBufCtr_clock = clock; // @[:@18773.4]
  assign NBufCtr_reset = reset; // @[:@18774.4]
  assign NBufCtr_io_input_countUp = 1'h0; // @[NBuffers.scala 43:24:@18781.4]
  assign NBufCtr_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 42:23:@18780.4]
  assign statesInR_0_clock = clock; // @[:@18784.4]
  assign statesInR_0_reset = reset; // @[:@18785.4]
  assign statesInR_0_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@18792.4]
  assign statesInR_0_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@18791.4]
  assign statesInR_1_clock = clock; // @[:@18795.4]
  assign statesInR_1_reset = reset; // @[:@18796.4]
  assign statesInR_1_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@18803.4]
  assign statesInR_1_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@18802.4]
  assign statesInR_2_clock = clock; // @[:@18806.4]
  assign statesInR_2_reset = reset; // @[:@18807.4]
  assign statesInR_2_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@18814.4]
  assign statesInR_2_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@18813.4]
  assign statesInR_3_clock = clock; // @[:@18817.4]
  assign statesInR_3_reset = reset; // @[:@18818.4]
  assign statesInR_3_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@18825.4]
  assign statesInR_3_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@18824.4]
  assign statesInR_4_clock = clock; // @[:@18828.4]
  assign statesInR_4_reset = reset; // @[:@18829.4]
  assign statesInR_4_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@18836.4]
  assign statesInR_4_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@18835.4]
  assign statesInR_5_clock = clock; // @[:@18839.4]
  assign statesInR_5_reset = reset; // @[:@18840.4]
  assign statesInR_5_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@18847.4]
  assign statesInR_5_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@18846.4]
  assign statesInR_6_clock = clock; // @[:@18850.4]
  assign statesInR_6_reset = reset; // @[:@18851.4]
  assign statesInR_6_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@18858.4]
  assign statesInR_6_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@18857.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_167 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_167 <= 1'h0;
    end else begin
      _T_167 <= _T_164;
    end
  end
endmodule
module FF_13( // @[:@18861.2]
  input         clock, // @[:@18862.4]
  input         reset, // @[:@18863.4]
  output [31:0] io_rPort_5_output_0, // @[:@18864.4]
  output [31:0] io_rPort_4_output_0, // @[:@18864.4]
  output [31:0] io_rPort_3_output_0, // @[:@18864.4]
  output [31:0] io_rPort_2_output_0, // @[:@18864.4]
  output [31:0] io_rPort_1_output_0, // @[:@18864.4]
  output [31:0] io_rPort_0_output_0, // @[:@18864.4]
  input  [31:0] io_wPort_0_data_0, // @[:@18864.4]
  input         io_wPort_0_reset, // @[:@18864.4]
  input         io_wPort_0_en_0 // @[:@18864.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@18904.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_198; // @[MemPrimitives.scala 325:32:@18906.4]
  wire [31:0] _T_199; // @[MemPrimitives.scala 325:12:@18907.4]
  assign _T_198 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@18906.4]
  assign _T_199 = io_wPort_0_reset ? 32'h0 : _T_198; // @[MemPrimitives.scala 325:12:@18907.4]
  assign io_rPort_5_output_0 = ff; // @[MemPrimitives.scala 326:34:@18914.4]
  assign io_rPort_4_output_0 = ff; // @[MemPrimitives.scala 326:34:@18913.4]
  assign io_rPort_3_output_0 = ff; // @[MemPrimitives.scala 326:34:@18912.4]
  assign io_rPort_2_output_0 = ff; // @[MemPrimitives.scala 326:34:@18911.4]
  assign io_rPort_1_output_0 = ff; // @[MemPrimitives.scala 326:34:@18910.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@18909.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module NBuf_2( // @[:@19246.2]
  input         clock, // @[:@19247.4]
  input         reset, // @[:@19248.4]
  output [31:0] io_rPort_5_output_0, // @[:@19249.4]
  output [31:0] io_rPort_4_output_0, // @[:@19249.4]
  output [31:0] io_rPort_3_output_0, // @[:@19249.4]
  output [31:0] io_rPort_2_output_0, // @[:@19249.4]
  output [31:0] io_rPort_1_output_0, // @[:@19249.4]
  output [31:0] io_rPort_0_output_0, // @[:@19249.4]
  input  [31:0] io_wPort_0_data_0, // @[:@19249.4]
  input         io_wPort_0_reset, // @[:@19249.4]
  input         io_wPort_0_en_0, // @[:@19249.4]
  input         io_sEn_0, // @[:@19249.4]
  input         io_sEn_1, // @[:@19249.4]
  input         io_sEn_2, // @[:@19249.4]
  input         io_sEn_3, // @[:@19249.4]
  input         io_sEn_4, // @[:@19249.4]
  input         io_sEn_5, // @[:@19249.4]
  input         io_sEn_6, // @[:@19249.4]
  input         io_sDone_0, // @[:@19249.4]
  input         io_sDone_1, // @[:@19249.4]
  input         io_sDone_2, // @[:@19249.4]
  input         io_sDone_3, // @[:@19249.4]
  input         io_sDone_4, // @[:@19249.4]
  input         io_sDone_5, // @[:@19249.4]
  input         io_sDone_6 // @[:@19249.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@19257.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@19257.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@19257.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@19257.4]
  wire  ctrl_io_sEn_2; // @[NBuffers.scala 83:20:@19257.4]
  wire  ctrl_io_sEn_3; // @[NBuffers.scala 83:20:@19257.4]
  wire  ctrl_io_sEn_4; // @[NBuffers.scala 83:20:@19257.4]
  wire  ctrl_io_sEn_5; // @[NBuffers.scala 83:20:@19257.4]
  wire  ctrl_io_sEn_6; // @[NBuffers.scala 83:20:@19257.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@19257.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@19257.4]
  wire  ctrl_io_sDone_2; // @[NBuffers.scala 83:20:@19257.4]
  wire  ctrl_io_sDone_3; // @[NBuffers.scala 83:20:@19257.4]
  wire  ctrl_io_sDone_4; // @[NBuffers.scala 83:20:@19257.4]
  wire  ctrl_io_sDone_5; // @[NBuffers.scala 83:20:@19257.4]
  wire  ctrl_io_sDone_6; // @[NBuffers.scala 83:20:@19257.4]
  wire [3:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@19257.4]
  wire [3:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@19257.4]
  wire [3:0] ctrl_io_statesInR_2; // @[NBuffers.scala 83:20:@19257.4]
  wire [3:0] ctrl_io_statesInR_3; // @[NBuffers.scala 83:20:@19257.4]
  wire [3:0] ctrl_io_statesInR_4; // @[NBuffers.scala 83:20:@19257.4]
  wire [3:0] ctrl_io_statesInR_5; // @[NBuffers.scala 83:20:@19257.4]
  wire [3:0] ctrl_io_statesInR_6; // @[NBuffers.scala 83:20:@19257.4]
  wire  FF_clock; // @[NBuffers.scala 146:23:@19274.4]
  wire  FF_reset; // @[NBuffers.scala 146:23:@19274.4]
  wire [31:0] FF_io_rPort_5_output_0; // @[NBuffers.scala 146:23:@19274.4]
  wire [31:0] FF_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@19274.4]
  wire [31:0] FF_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@19274.4]
  wire [31:0] FF_io_rPort_2_output_0; // @[NBuffers.scala 146:23:@19274.4]
  wire [31:0] FF_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@19274.4]
  wire [31:0] FF_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@19274.4]
  wire [31:0] FF_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@19274.4]
  wire  FF_io_wPort_0_reset; // @[NBuffers.scala 146:23:@19274.4]
  wire  FF_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@19274.4]
  wire  FF_1_clock; // @[NBuffers.scala 146:23:@19315.4]
  wire  FF_1_reset; // @[NBuffers.scala 146:23:@19315.4]
  wire [31:0] FF_1_io_rPort_5_output_0; // @[NBuffers.scala 146:23:@19315.4]
  wire [31:0] FF_1_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@19315.4]
  wire [31:0] FF_1_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@19315.4]
  wire [31:0] FF_1_io_rPort_2_output_0; // @[NBuffers.scala 146:23:@19315.4]
  wire [31:0] FF_1_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@19315.4]
  wire [31:0] FF_1_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@19315.4]
  wire [31:0] FF_1_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@19315.4]
  wire  FF_1_io_wPort_0_reset; // @[NBuffers.scala 146:23:@19315.4]
  wire  FF_1_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@19315.4]
  wire  FF_2_clock; // @[NBuffers.scala 146:23:@19356.4]
  wire  FF_2_reset; // @[NBuffers.scala 146:23:@19356.4]
  wire [31:0] FF_2_io_rPort_5_output_0; // @[NBuffers.scala 146:23:@19356.4]
  wire [31:0] FF_2_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@19356.4]
  wire [31:0] FF_2_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@19356.4]
  wire [31:0] FF_2_io_rPort_2_output_0; // @[NBuffers.scala 146:23:@19356.4]
  wire [31:0] FF_2_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@19356.4]
  wire [31:0] FF_2_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@19356.4]
  wire [31:0] FF_2_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@19356.4]
  wire  FF_2_io_wPort_0_reset; // @[NBuffers.scala 146:23:@19356.4]
  wire  FF_2_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@19356.4]
  wire  FF_3_clock; // @[NBuffers.scala 146:23:@19397.4]
  wire  FF_3_reset; // @[NBuffers.scala 146:23:@19397.4]
  wire [31:0] FF_3_io_rPort_5_output_0; // @[NBuffers.scala 146:23:@19397.4]
  wire [31:0] FF_3_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@19397.4]
  wire [31:0] FF_3_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@19397.4]
  wire [31:0] FF_3_io_rPort_2_output_0; // @[NBuffers.scala 146:23:@19397.4]
  wire [31:0] FF_3_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@19397.4]
  wire [31:0] FF_3_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@19397.4]
  wire [31:0] FF_3_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@19397.4]
  wire  FF_3_io_wPort_0_reset; // @[NBuffers.scala 146:23:@19397.4]
  wire  FF_3_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@19397.4]
  wire  FF_4_clock; // @[NBuffers.scala 146:23:@19438.4]
  wire  FF_4_reset; // @[NBuffers.scala 146:23:@19438.4]
  wire [31:0] FF_4_io_rPort_5_output_0; // @[NBuffers.scala 146:23:@19438.4]
  wire [31:0] FF_4_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@19438.4]
  wire [31:0] FF_4_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@19438.4]
  wire [31:0] FF_4_io_rPort_2_output_0; // @[NBuffers.scala 146:23:@19438.4]
  wire [31:0] FF_4_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@19438.4]
  wire [31:0] FF_4_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@19438.4]
  wire [31:0] FF_4_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@19438.4]
  wire  FF_4_io_wPort_0_reset; // @[NBuffers.scala 146:23:@19438.4]
  wire  FF_4_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@19438.4]
  wire  FF_5_clock; // @[NBuffers.scala 146:23:@19479.4]
  wire  FF_5_reset; // @[NBuffers.scala 146:23:@19479.4]
  wire [31:0] FF_5_io_rPort_5_output_0; // @[NBuffers.scala 146:23:@19479.4]
  wire [31:0] FF_5_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@19479.4]
  wire [31:0] FF_5_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@19479.4]
  wire [31:0] FF_5_io_rPort_2_output_0; // @[NBuffers.scala 146:23:@19479.4]
  wire [31:0] FF_5_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@19479.4]
  wire [31:0] FF_5_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@19479.4]
  wire [31:0] FF_5_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@19479.4]
  wire  FF_5_io_wPort_0_reset; // @[NBuffers.scala 146:23:@19479.4]
  wire  FF_5_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@19479.4]
  wire  FF_6_clock; // @[NBuffers.scala 146:23:@19520.4]
  wire  FF_6_reset; // @[NBuffers.scala 146:23:@19520.4]
  wire [31:0] FF_6_io_rPort_5_output_0; // @[NBuffers.scala 146:23:@19520.4]
  wire [31:0] FF_6_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@19520.4]
  wire [31:0] FF_6_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@19520.4]
  wire [31:0] FF_6_io_rPort_2_output_0; // @[NBuffers.scala 146:23:@19520.4]
  wire [31:0] FF_6_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@19520.4]
  wire [31:0] FF_6_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@19520.4]
  wire [31:0] FF_6_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@19520.4]
  wire  FF_6_io_wPort_0_reset; // @[NBuffers.scala 146:23:@19520.4]
  wire  FF_6_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@19520.4]
  wire  _T_236; // @[NBuffers.scala 153:105:@19568.4]
  wire  _T_240; // @[NBuffers.scala 157:92:@19578.4]
  wire  _T_243; // @[NBuffers.scala 157:92:@19584.4]
  wire  _T_246; // @[NBuffers.scala 157:92:@19590.4]
  wire  _T_249; // @[NBuffers.scala 157:92:@19596.4]
  wire  _T_252; // @[NBuffers.scala 157:92:@19602.4]
  wire  _T_255; // @[NBuffers.scala 157:92:@19608.4]
  wire  _T_258; // @[NBuffers.scala 153:105:@19614.4]
  wire  _T_262; // @[NBuffers.scala 157:92:@19624.4]
  wire  _T_265; // @[NBuffers.scala 157:92:@19630.4]
  wire  _T_268; // @[NBuffers.scala 157:92:@19636.4]
  wire  _T_271; // @[NBuffers.scala 157:92:@19642.4]
  wire  _T_274; // @[NBuffers.scala 157:92:@19648.4]
  wire  _T_277; // @[NBuffers.scala 157:92:@19654.4]
  wire  _T_280; // @[NBuffers.scala 153:105:@19660.4]
  wire  _T_284; // @[NBuffers.scala 157:92:@19670.4]
  wire  _T_287; // @[NBuffers.scala 157:92:@19676.4]
  wire  _T_290; // @[NBuffers.scala 157:92:@19682.4]
  wire  _T_293; // @[NBuffers.scala 157:92:@19688.4]
  wire  _T_296; // @[NBuffers.scala 157:92:@19694.4]
  wire  _T_299; // @[NBuffers.scala 157:92:@19700.4]
  wire  _T_302; // @[NBuffers.scala 153:105:@19706.4]
  wire  _T_306; // @[NBuffers.scala 157:92:@19716.4]
  wire  _T_309; // @[NBuffers.scala 157:92:@19722.4]
  wire  _T_312; // @[NBuffers.scala 157:92:@19728.4]
  wire  _T_315; // @[NBuffers.scala 157:92:@19734.4]
  wire  _T_318; // @[NBuffers.scala 157:92:@19740.4]
  wire  _T_321; // @[NBuffers.scala 157:92:@19746.4]
  wire  _T_324; // @[NBuffers.scala 153:105:@19752.4]
  wire  _T_328; // @[NBuffers.scala 157:92:@19762.4]
  wire  _T_331; // @[NBuffers.scala 157:92:@19768.4]
  wire  _T_334; // @[NBuffers.scala 157:92:@19774.4]
  wire  _T_337; // @[NBuffers.scala 157:92:@19780.4]
  wire  _T_340; // @[NBuffers.scala 157:92:@19786.4]
  wire  _T_343; // @[NBuffers.scala 157:92:@19792.4]
  wire  _T_346; // @[NBuffers.scala 153:105:@19798.4]
  wire  _T_350; // @[NBuffers.scala 157:92:@19808.4]
  wire  _T_353; // @[NBuffers.scala 157:92:@19814.4]
  wire  _T_356; // @[NBuffers.scala 157:92:@19820.4]
  wire  _T_359; // @[NBuffers.scala 157:92:@19826.4]
  wire  _T_362; // @[NBuffers.scala 157:92:@19832.4]
  wire  _T_365; // @[NBuffers.scala 157:92:@19838.4]
  wire  _T_368; // @[NBuffers.scala 153:105:@19844.4]
  wire  _T_372; // @[NBuffers.scala 157:92:@19854.4]
  wire  _T_375; // @[NBuffers.scala 157:92:@19860.4]
  wire  _T_378; // @[NBuffers.scala 157:92:@19866.4]
  wire  _T_381; // @[NBuffers.scala 157:92:@19872.4]
  wire  _T_384; // @[NBuffers.scala 157:92:@19878.4]
  wire  _T_387; // @[NBuffers.scala 157:92:@19884.4]
  wire [31:0] _T_405; // @[Mux.scala 19:72:@19897.4]
  wire [31:0] _T_407; // @[Mux.scala 19:72:@19898.4]
  wire [31:0] _T_409; // @[Mux.scala 19:72:@19899.4]
  wire [31:0] _T_411; // @[Mux.scala 19:72:@19900.4]
  wire [31:0] _T_413; // @[Mux.scala 19:72:@19901.4]
  wire [31:0] _T_415; // @[Mux.scala 19:72:@19902.4]
  wire [31:0] _T_417; // @[Mux.scala 19:72:@19903.4]
  wire [31:0] _T_418; // @[Mux.scala 19:72:@19904.4]
  wire [31:0] _T_419; // @[Mux.scala 19:72:@19905.4]
  wire [31:0] _T_420; // @[Mux.scala 19:72:@19906.4]
  wire [31:0] _T_421; // @[Mux.scala 19:72:@19907.4]
  wire [31:0] _T_422; // @[Mux.scala 19:72:@19908.4]
  wire [31:0] _T_442; // @[Mux.scala 19:72:@19920.4]
  wire [31:0] _T_444; // @[Mux.scala 19:72:@19921.4]
  wire [31:0] _T_446; // @[Mux.scala 19:72:@19922.4]
  wire [31:0] _T_448; // @[Mux.scala 19:72:@19923.4]
  wire [31:0] _T_450; // @[Mux.scala 19:72:@19924.4]
  wire [31:0] _T_452; // @[Mux.scala 19:72:@19925.4]
  wire [31:0] _T_454; // @[Mux.scala 19:72:@19926.4]
  wire [31:0] _T_455; // @[Mux.scala 19:72:@19927.4]
  wire [31:0] _T_456; // @[Mux.scala 19:72:@19928.4]
  wire [31:0] _T_457; // @[Mux.scala 19:72:@19929.4]
  wire [31:0] _T_458; // @[Mux.scala 19:72:@19930.4]
  wire [31:0] _T_459; // @[Mux.scala 19:72:@19931.4]
  wire [31:0] _T_479; // @[Mux.scala 19:72:@19943.4]
  wire [31:0] _T_481; // @[Mux.scala 19:72:@19944.4]
  wire [31:0] _T_483; // @[Mux.scala 19:72:@19945.4]
  wire [31:0] _T_485; // @[Mux.scala 19:72:@19946.4]
  wire [31:0] _T_487; // @[Mux.scala 19:72:@19947.4]
  wire [31:0] _T_489; // @[Mux.scala 19:72:@19948.4]
  wire [31:0] _T_491; // @[Mux.scala 19:72:@19949.4]
  wire [31:0] _T_492; // @[Mux.scala 19:72:@19950.4]
  wire [31:0] _T_493; // @[Mux.scala 19:72:@19951.4]
  wire [31:0] _T_494; // @[Mux.scala 19:72:@19952.4]
  wire [31:0] _T_495; // @[Mux.scala 19:72:@19953.4]
  wire [31:0] _T_496; // @[Mux.scala 19:72:@19954.4]
  wire [31:0] _T_516; // @[Mux.scala 19:72:@19966.4]
  wire [31:0] _T_518; // @[Mux.scala 19:72:@19967.4]
  wire [31:0] _T_520; // @[Mux.scala 19:72:@19968.4]
  wire [31:0] _T_522; // @[Mux.scala 19:72:@19969.4]
  wire [31:0] _T_524; // @[Mux.scala 19:72:@19970.4]
  wire [31:0] _T_526; // @[Mux.scala 19:72:@19971.4]
  wire [31:0] _T_528; // @[Mux.scala 19:72:@19972.4]
  wire [31:0] _T_529; // @[Mux.scala 19:72:@19973.4]
  wire [31:0] _T_530; // @[Mux.scala 19:72:@19974.4]
  wire [31:0] _T_531; // @[Mux.scala 19:72:@19975.4]
  wire [31:0] _T_532; // @[Mux.scala 19:72:@19976.4]
  wire [31:0] _T_533; // @[Mux.scala 19:72:@19977.4]
  wire [31:0] _T_553; // @[Mux.scala 19:72:@19989.4]
  wire [31:0] _T_555; // @[Mux.scala 19:72:@19990.4]
  wire [31:0] _T_557; // @[Mux.scala 19:72:@19991.4]
  wire [31:0] _T_559; // @[Mux.scala 19:72:@19992.4]
  wire [31:0] _T_561; // @[Mux.scala 19:72:@19993.4]
  wire [31:0] _T_563; // @[Mux.scala 19:72:@19994.4]
  wire [31:0] _T_565; // @[Mux.scala 19:72:@19995.4]
  wire [31:0] _T_566; // @[Mux.scala 19:72:@19996.4]
  wire [31:0] _T_567; // @[Mux.scala 19:72:@19997.4]
  wire [31:0] _T_568; // @[Mux.scala 19:72:@19998.4]
  wire [31:0] _T_569; // @[Mux.scala 19:72:@19999.4]
  wire [31:0] _T_570; // @[Mux.scala 19:72:@20000.4]
  wire [31:0] _T_590; // @[Mux.scala 19:72:@20012.4]
  wire [31:0] _T_592; // @[Mux.scala 19:72:@20013.4]
  wire [31:0] _T_594; // @[Mux.scala 19:72:@20014.4]
  wire [31:0] _T_596; // @[Mux.scala 19:72:@20015.4]
  wire [31:0] _T_598; // @[Mux.scala 19:72:@20016.4]
  wire [31:0] _T_600; // @[Mux.scala 19:72:@20017.4]
  wire [31:0] _T_602; // @[Mux.scala 19:72:@20018.4]
  wire [31:0] _T_603; // @[Mux.scala 19:72:@20019.4]
  wire [31:0] _T_604; // @[Mux.scala 19:72:@20020.4]
  wire [31:0] _T_605; // @[Mux.scala 19:72:@20021.4]
  wire [31:0] _T_606; // @[Mux.scala 19:72:@20022.4]
  wire [31:0] _T_607; // @[Mux.scala 19:72:@20023.4]
  NBufController_3 ctrl ( // @[NBuffers.scala 83:20:@19257.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sEn_2(ctrl_io_sEn_2),
    .io_sEn_3(ctrl_io_sEn_3),
    .io_sEn_4(ctrl_io_sEn_4),
    .io_sEn_5(ctrl_io_sEn_5),
    .io_sEn_6(ctrl_io_sEn_6),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_sDone_2(ctrl_io_sDone_2),
    .io_sDone_3(ctrl_io_sDone_3),
    .io_sDone_4(ctrl_io_sDone_4),
    .io_sDone_5(ctrl_io_sDone_5),
    .io_sDone_6(ctrl_io_sDone_6),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1),
    .io_statesInR_2(ctrl_io_statesInR_2),
    .io_statesInR_3(ctrl_io_statesInR_3),
    .io_statesInR_4(ctrl_io_statesInR_4),
    .io_statesInR_5(ctrl_io_statesInR_5),
    .io_statesInR_6(ctrl_io_statesInR_6)
  );
  FF_13 FF ( // @[NBuffers.scala 146:23:@19274.4]
    .clock(FF_clock),
    .reset(FF_reset),
    .io_rPort_5_output_0(FF_io_rPort_5_output_0),
    .io_rPort_4_output_0(FF_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_io_rPort_3_output_0),
    .io_rPort_2_output_0(FF_io_rPort_2_output_0),
    .io_rPort_1_output_0(FF_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_io_wPort_0_en_0)
  );
  FF_13 FF_1 ( // @[NBuffers.scala 146:23:@19315.4]
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_rPort_5_output_0(FF_1_io_rPort_5_output_0),
    .io_rPort_4_output_0(FF_1_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_1_io_rPort_3_output_0),
    .io_rPort_2_output_0(FF_1_io_rPort_2_output_0),
    .io_rPort_1_output_0(FF_1_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_1_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_1_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_1_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_1_io_wPort_0_en_0)
  );
  FF_13 FF_2 ( // @[NBuffers.scala 146:23:@19356.4]
    .clock(FF_2_clock),
    .reset(FF_2_reset),
    .io_rPort_5_output_0(FF_2_io_rPort_5_output_0),
    .io_rPort_4_output_0(FF_2_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_2_io_rPort_3_output_0),
    .io_rPort_2_output_0(FF_2_io_rPort_2_output_0),
    .io_rPort_1_output_0(FF_2_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_2_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_2_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_2_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_2_io_wPort_0_en_0)
  );
  FF_13 FF_3 ( // @[NBuffers.scala 146:23:@19397.4]
    .clock(FF_3_clock),
    .reset(FF_3_reset),
    .io_rPort_5_output_0(FF_3_io_rPort_5_output_0),
    .io_rPort_4_output_0(FF_3_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_3_io_rPort_3_output_0),
    .io_rPort_2_output_0(FF_3_io_rPort_2_output_0),
    .io_rPort_1_output_0(FF_3_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_3_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_3_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_3_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_3_io_wPort_0_en_0)
  );
  FF_13 FF_4 ( // @[NBuffers.scala 146:23:@19438.4]
    .clock(FF_4_clock),
    .reset(FF_4_reset),
    .io_rPort_5_output_0(FF_4_io_rPort_5_output_0),
    .io_rPort_4_output_0(FF_4_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_4_io_rPort_3_output_0),
    .io_rPort_2_output_0(FF_4_io_rPort_2_output_0),
    .io_rPort_1_output_0(FF_4_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_4_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_4_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_4_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_4_io_wPort_0_en_0)
  );
  FF_13 FF_5 ( // @[NBuffers.scala 146:23:@19479.4]
    .clock(FF_5_clock),
    .reset(FF_5_reset),
    .io_rPort_5_output_0(FF_5_io_rPort_5_output_0),
    .io_rPort_4_output_0(FF_5_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_5_io_rPort_3_output_0),
    .io_rPort_2_output_0(FF_5_io_rPort_2_output_0),
    .io_rPort_1_output_0(FF_5_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_5_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_5_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_5_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_5_io_wPort_0_en_0)
  );
  FF_13 FF_6 ( // @[NBuffers.scala 146:23:@19520.4]
    .clock(FF_6_clock),
    .reset(FF_6_reset),
    .io_rPort_5_output_0(FF_6_io_rPort_5_output_0),
    .io_rPort_4_output_0(FF_6_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_6_io_rPort_3_output_0),
    .io_rPort_2_output_0(FF_6_io_rPort_2_output_0),
    .io_rPort_1_output_0(FF_6_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_6_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_6_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_6_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_6_io_wPort_0_en_0)
  );
  assign _T_236 = ctrl_io_statesInW_0 == 4'h0; // @[NBuffers.scala 153:105:@19568.4]
  assign _T_240 = ctrl_io_statesInR_1 == 4'h0; // @[NBuffers.scala 157:92:@19578.4]
  assign _T_243 = ctrl_io_statesInR_2 == 4'h0; // @[NBuffers.scala 157:92:@19584.4]
  assign _T_246 = ctrl_io_statesInR_3 == 4'h0; // @[NBuffers.scala 157:92:@19590.4]
  assign _T_249 = ctrl_io_statesInR_4 == 4'h0; // @[NBuffers.scala 157:92:@19596.4]
  assign _T_252 = ctrl_io_statesInR_5 == 4'h0; // @[NBuffers.scala 157:92:@19602.4]
  assign _T_255 = ctrl_io_statesInR_6 == 4'h0; // @[NBuffers.scala 157:92:@19608.4]
  assign _T_258 = ctrl_io_statesInW_0 == 4'h1; // @[NBuffers.scala 153:105:@19614.4]
  assign _T_262 = ctrl_io_statesInR_1 == 4'h1; // @[NBuffers.scala 157:92:@19624.4]
  assign _T_265 = ctrl_io_statesInR_2 == 4'h1; // @[NBuffers.scala 157:92:@19630.4]
  assign _T_268 = ctrl_io_statesInR_3 == 4'h1; // @[NBuffers.scala 157:92:@19636.4]
  assign _T_271 = ctrl_io_statesInR_4 == 4'h1; // @[NBuffers.scala 157:92:@19642.4]
  assign _T_274 = ctrl_io_statesInR_5 == 4'h1; // @[NBuffers.scala 157:92:@19648.4]
  assign _T_277 = ctrl_io_statesInR_6 == 4'h1; // @[NBuffers.scala 157:92:@19654.4]
  assign _T_280 = ctrl_io_statesInW_0 == 4'h2; // @[NBuffers.scala 153:105:@19660.4]
  assign _T_284 = ctrl_io_statesInR_1 == 4'h2; // @[NBuffers.scala 157:92:@19670.4]
  assign _T_287 = ctrl_io_statesInR_2 == 4'h2; // @[NBuffers.scala 157:92:@19676.4]
  assign _T_290 = ctrl_io_statesInR_3 == 4'h2; // @[NBuffers.scala 157:92:@19682.4]
  assign _T_293 = ctrl_io_statesInR_4 == 4'h2; // @[NBuffers.scala 157:92:@19688.4]
  assign _T_296 = ctrl_io_statesInR_5 == 4'h2; // @[NBuffers.scala 157:92:@19694.4]
  assign _T_299 = ctrl_io_statesInR_6 == 4'h2; // @[NBuffers.scala 157:92:@19700.4]
  assign _T_302 = ctrl_io_statesInW_0 == 4'h3; // @[NBuffers.scala 153:105:@19706.4]
  assign _T_306 = ctrl_io_statesInR_1 == 4'h3; // @[NBuffers.scala 157:92:@19716.4]
  assign _T_309 = ctrl_io_statesInR_2 == 4'h3; // @[NBuffers.scala 157:92:@19722.4]
  assign _T_312 = ctrl_io_statesInR_3 == 4'h3; // @[NBuffers.scala 157:92:@19728.4]
  assign _T_315 = ctrl_io_statesInR_4 == 4'h3; // @[NBuffers.scala 157:92:@19734.4]
  assign _T_318 = ctrl_io_statesInR_5 == 4'h3; // @[NBuffers.scala 157:92:@19740.4]
  assign _T_321 = ctrl_io_statesInR_6 == 4'h3; // @[NBuffers.scala 157:92:@19746.4]
  assign _T_324 = ctrl_io_statesInW_0 == 4'h4; // @[NBuffers.scala 153:105:@19752.4]
  assign _T_328 = ctrl_io_statesInR_1 == 4'h4; // @[NBuffers.scala 157:92:@19762.4]
  assign _T_331 = ctrl_io_statesInR_2 == 4'h4; // @[NBuffers.scala 157:92:@19768.4]
  assign _T_334 = ctrl_io_statesInR_3 == 4'h4; // @[NBuffers.scala 157:92:@19774.4]
  assign _T_337 = ctrl_io_statesInR_4 == 4'h4; // @[NBuffers.scala 157:92:@19780.4]
  assign _T_340 = ctrl_io_statesInR_5 == 4'h4; // @[NBuffers.scala 157:92:@19786.4]
  assign _T_343 = ctrl_io_statesInR_6 == 4'h4; // @[NBuffers.scala 157:92:@19792.4]
  assign _T_346 = ctrl_io_statesInW_0 == 4'h5; // @[NBuffers.scala 153:105:@19798.4]
  assign _T_350 = ctrl_io_statesInR_1 == 4'h5; // @[NBuffers.scala 157:92:@19808.4]
  assign _T_353 = ctrl_io_statesInR_2 == 4'h5; // @[NBuffers.scala 157:92:@19814.4]
  assign _T_356 = ctrl_io_statesInR_3 == 4'h5; // @[NBuffers.scala 157:92:@19820.4]
  assign _T_359 = ctrl_io_statesInR_4 == 4'h5; // @[NBuffers.scala 157:92:@19826.4]
  assign _T_362 = ctrl_io_statesInR_5 == 4'h5; // @[NBuffers.scala 157:92:@19832.4]
  assign _T_365 = ctrl_io_statesInR_6 == 4'h5; // @[NBuffers.scala 157:92:@19838.4]
  assign _T_368 = ctrl_io_statesInW_0 == 4'h6; // @[NBuffers.scala 153:105:@19844.4]
  assign _T_372 = ctrl_io_statesInR_1 == 4'h6; // @[NBuffers.scala 157:92:@19854.4]
  assign _T_375 = ctrl_io_statesInR_2 == 4'h6; // @[NBuffers.scala 157:92:@19860.4]
  assign _T_378 = ctrl_io_statesInR_3 == 4'h6; // @[NBuffers.scala 157:92:@19866.4]
  assign _T_381 = ctrl_io_statesInR_4 == 4'h6; // @[NBuffers.scala 157:92:@19872.4]
  assign _T_384 = ctrl_io_statesInR_5 == 4'h6; // @[NBuffers.scala 157:92:@19878.4]
  assign _T_387 = ctrl_io_statesInR_6 == 4'h6; // @[NBuffers.scala 157:92:@19884.4]
  assign _T_405 = _T_240 ? FF_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@19897.4]
  assign _T_407 = _T_262 ? FF_1_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@19898.4]
  assign _T_409 = _T_284 ? FF_2_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@19899.4]
  assign _T_411 = _T_306 ? FF_3_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@19900.4]
  assign _T_413 = _T_328 ? FF_4_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@19901.4]
  assign _T_415 = _T_350 ? FF_5_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@19902.4]
  assign _T_417 = _T_372 ? FF_6_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@19903.4]
  assign _T_418 = _T_405 | _T_407; // @[Mux.scala 19:72:@19904.4]
  assign _T_419 = _T_418 | _T_409; // @[Mux.scala 19:72:@19905.4]
  assign _T_420 = _T_419 | _T_411; // @[Mux.scala 19:72:@19906.4]
  assign _T_421 = _T_420 | _T_413; // @[Mux.scala 19:72:@19907.4]
  assign _T_422 = _T_421 | _T_415; // @[Mux.scala 19:72:@19908.4]
  assign _T_442 = _T_243 ? FF_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@19920.4]
  assign _T_444 = _T_265 ? FF_1_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@19921.4]
  assign _T_446 = _T_287 ? FF_2_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@19922.4]
  assign _T_448 = _T_309 ? FF_3_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@19923.4]
  assign _T_450 = _T_331 ? FF_4_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@19924.4]
  assign _T_452 = _T_353 ? FF_5_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@19925.4]
  assign _T_454 = _T_375 ? FF_6_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@19926.4]
  assign _T_455 = _T_442 | _T_444; // @[Mux.scala 19:72:@19927.4]
  assign _T_456 = _T_455 | _T_446; // @[Mux.scala 19:72:@19928.4]
  assign _T_457 = _T_456 | _T_448; // @[Mux.scala 19:72:@19929.4]
  assign _T_458 = _T_457 | _T_450; // @[Mux.scala 19:72:@19930.4]
  assign _T_459 = _T_458 | _T_452; // @[Mux.scala 19:72:@19931.4]
  assign _T_479 = _T_246 ? FF_io_rPort_2_output_0 : 32'h0; // @[Mux.scala 19:72:@19943.4]
  assign _T_481 = _T_268 ? FF_1_io_rPort_2_output_0 : 32'h0; // @[Mux.scala 19:72:@19944.4]
  assign _T_483 = _T_290 ? FF_2_io_rPort_2_output_0 : 32'h0; // @[Mux.scala 19:72:@19945.4]
  assign _T_485 = _T_312 ? FF_3_io_rPort_2_output_0 : 32'h0; // @[Mux.scala 19:72:@19946.4]
  assign _T_487 = _T_334 ? FF_4_io_rPort_2_output_0 : 32'h0; // @[Mux.scala 19:72:@19947.4]
  assign _T_489 = _T_356 ? FF_5_io_rPort_2_output_0 : 32'h0; // @[Mux.scala 19:72:@19948.4]
  assign _T_491 = _T_378 ? FF_6_io_rPort_2_output_0 : 32'h0; // @[Mux.scala 19:72:@19949.4]
  assign _T_492 = _T_479 | _T_481; // @[Mux.scala 19:72:@19950.4]
  assign _T_493 = _T_492 | _T_483; // @[Mux.scala 19:72:@19951.4]
  assign _T_494 = _T_493 | _T_485; // @[Mux.scala 19:72:@19952.4]
  assign _T_495 = _T_494 | _T_487; // @[Mux.scala 19:72:@19953.4]
  assign _T_496 = _T_495 | _T_489; // @[Mux.scala 19:72:@19954.4]
  assign _T_516 = _T_249 ? FF_io_rPort_3_output_0 : 32'h0; // @[Mux.scala 19:72:@19966.4]
  assign _T_518 = _T_271 ? FF_1_io_rPort_3_output_0 : 32'h0; // @[Mux.scala 19:72:@19967.4]
  assign _T_520 = _T_293 ? FF_2_io_rPort_3_output_0 : 32'h0; // @[Mux.scala 19:72:@19968.4]
  assign _T_522 = _T_315 ? FF_3_io_rPort_3_output_0 : 32'h0; // @[Mux.scala 19:72:@19969.4]
  assign _T_524 = _T_337 ? FF_4_io_rPort_3_output_0 : 32'h0; // @[Mux.scala 19:72:@19970.4]
  assign _T_526 = _T_359 ? FF_5_io_rPort_3_output_0 : 32'h0; // @[Mux.scala 19:72:@19971.4]
  assign _T_528 = _T_381 ? FF_6_io_rPort_3_output_0 : 32'h0; // @[Mux.scala 19:72:@19972.4]
  assign _T_529 = _T_516 | _T_518; // @[Mux.scala 19:72:@19973.4]
  assign _T_530 = _T_529 | _T_520; // @[Mux.scala 19:72:@19974.4]
  assign _T_531 = _T_530 | _T_522; // @[Mux.scala 19:72:@19975.4]
  assign _T_532 = _T_531 | _T_524; // @[Mux.scala 19:72:@19976.4]
  assign _T_533 = _T_532 | _T_526; // @[Mux.scala 19:72:@19977.4]
  assign _T_553 = _T_252 ? FF_io_rPort_4_output_0 : 32'h0; // @[Mux.scala 19:72:@19989.4]
  assign _T_555 = _T_274 ? FF_1_io_rPort_4_output_0 : 32'h0; // @[Mux.scala 19:72:@19990.4]
  assign _T_557 = _T_296 ? FF_2_io_rPort_4_output_0 : 32'h0; // @[Mux.scala 19:72:@19991.4]
  assign _T_559 = _T_318 ? FF_3_io_rPort_4_output_0 : 32'h0; // @[Mux.scala 19:72:@19992.4]
  assign _T_561 = _T_340 ? FF_4_io_rPort_4_output_0 : 32'h0; // @[Mux.scala 19:72:@19993.4]
  assign _T_563 = _T_362 ? FF_5_io_rPort_4_output_0 : 32'h0; // @[Mux.scala 19:72:@19994.4]
  assign _T_565 = _T_384 ? FF_6_io_rPort_4_output_0 : 32'h0; // @[Mux.scala 19:72:@19995.4]
  assign _T_566 = _T_553 | _T_555; // @[Mux.scala 19:72:@19996.4]
  assign _T_567 = _T_566 | _T_557; // @[Mux.scala 19:72:@19997.4]
  assign _T_568 = _T_567 | _T_559; // @[Mux.scala 19:72:@19998.4]
  assign _T_569 = _T_568 | _T_561; // @[Mux.scala 19:72:@19999.4]
  assign _T_570 = _T_569 | _T_563; // @[Mux.scala 19:72:@20000.4]
  assign _T_590 = _T_255 ? FF_io_rPort_5_output_0 : 32'h0; // @[Mux.scala 19:72:@20012.4]
  assign _T_592 = _T_277 ? FF_1_io_rPort_5_output_0 : 32'h0; // @[Mux.scala 19:72:@20013.4]
  assign _T_594 = _T_299 ? FF_2_io_rPort_5_output_0 : 32'h0; // @[Mux.scala 19:72:@20014.4]
  assign _T_596 = _T_321 ? FF_3_io_rPort_5_output_0 : 32'h0; // @[Mux.scala 19:72:@20015.4]
  assign _T_598 = _T_343 ? FF_4_io_rPort_5_output_0 : 32'h0; // @[Mux.scala 19:72:@20016.4]
  assign _T_600 = _T_365 ? FF_5_io_rPort_5_output_0 : 32'h0; // @[Mux.scala 19:72:@20017.4]
  assign _T_602 = _T_387 ? FF_6_io_rPort_5_output_0 : 32'h0; // @[Mux.scala 19:72:@20018.4]
  assign _T_603 = _T_590 | _T_592; // @[Mux.scala 19:72:@20019.4]
  assign _T_604 = _T_603 | _T_594; // @[Mux.scala 19:72:@20020.4]
  assign _T_605 = _T_604 | _T_596; // @[Mux.scala 19:72:@20021.4]
  assign _T_606 = _T_605 | _T_598; // @[Mux.scala 19:72:@20022.4]
  assign _T_607 = _T_606 | _T_600; // @[Mux.scala 19:72:@20023.4]
  assign io_rPort_5_output_0 = _T_607 | _T_602; // @[NBuffers.scala 163:66:@20027.4]
  assign io_rPort_4_output_0 = _T_570 | _T_565; // @[NBuffers.scala 163:66:@20004.4]
  assign io_rPort_3_output_0 = _T_533 | _T_528; // @[NBuffers.scala 163:66:@19981.4]
  assign io_rPort_2_output_0 = _T_496 | _T_491; // @[NBuffers.scala 163:66:@19958.4]
  assign io_rPort_1_output_0 = _T_459 | _T_454; // @[NBuffers.scala 163:66:@19935.4]
  assign io_rPort_0_output_0 = _T_422 | _T_417; // @[NBuffers.scala 163:66:@19912.4]
  assign ctrl_clock = clock; // @[:@19258.4]
  assign ctrl_reset = reset; // @[:@19259.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@19260.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@19262.4]
  assign ctrl_io_sEn_2 = io_sEn_2; // @[NBuffers.scala 85:20:@19264.4]
  assign ctrl_io_sEn_3 = io_sEn_3; // @[NBuffers.scala 85:20:@19266.4]
  assign ctrl_io_sEn_4 = io_sEn_4; // @[NBuffers.scala 85:20:@19268.4]
  assign ctrl_io_sEn_5 = io_sEn_5; // @[NBuffers.scala 85:20:@19270.4]
  assign ctrl_io_sEn_6 = io_sEn_6; // @[NBuffers.scala 85:20:@19272.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@19261.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@19263.4]
  assign ctrl_io_sDone_2 = io_sDone_2; // @[NBuffers.scala 86:22:@19265.4]
  assign ctrl_io_sDone_3 = io_sDone_3; // @[NBuffers.scala 86:22:@19267.4]
  assign ctrl_io_sDone_4 = io_sDone_4; // @[NBuffers.scala 86:22:@19269.4]
  assign ctrl_io_sDone_5 = io_sDone_5; // @[NBuffers.scala 86:22:@19271.4]
  assign ctrl_io_sDone_6 = io_sDone_6; // @[NBuffers.scala 86:22:@19273.4]
  assign FF_clock = clock; // @[:@19275.4]
  assign FF_reset = reset; // @[:@19276.4]
  assign FF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@19571.4]
  assign FF_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@19572.4]
  assign FF_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_236; // @[MemPrimitives.scala 37:29:@19577.4]
  assign FF_1_clock = clock; // @[:@19316.4]
  assign FF_1_reset = reset; // @[:@19317.4]
  assign FF_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@19617.4]
  assign FF_1_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@19618.4]
  assign FF_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_258; // @[MemPrimitives.scala 37:29:@19623.4]
  assign FF_2_clock = clock; // @[:@19357.4]
  assign FF_2_reset = reset; // @[:@19358.4]
  assign FF_2_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@19663.4]
  assign FF_2_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@19664.4]
  assign FF_2_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_280; // @[MemPrimitives.scala 37:29:@19669.4]
  assign FF_3_clock = clock; // @[:@19398.4]
  assign FF_3_reset = reset; // @[:@19399.4]
  assign FF_3_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@19709.4]
  assign FF_3_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@19710.4]
  assign FF_3_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_302; // @[MemPrimitives.scala 37:29:@19715.4]
  assign FF_4_clock = clock; // @[:@19439.4]
  assign FF_4_reset = reset; // @[:@19440.4]
  assign FF_4_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@19755.4]
  assign FF_4_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@19756.4]
  assign FF_4_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_324; // @[MemPrimitives.scala 37:29:@19761.4]
  assign FF_5_clock = clock; // @[:@19480.4]
  assign FF_5_reset = reset; // @[:@19481.4]
  assign FF_5_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@19801.4]
  assign FF_5_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@19802.4]
  assign FF_5_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_346; // @[MemPrimitives.scala 37:29:@19807.4]
  assign FF_6_clock = clock; // @[:@19521.4]
  assign FF_6_reset = reset; // @[:@19522.4]
  assign FF_6_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@19847.4]
  assign FF_6_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@19848.4]
  assign FF_6_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_368; // @[MemPrimitives.scala 37:29:@19853.4]
endmodule
module b550_chain( // @[:@20029.2]
  input         clock, // @[:@20030.4]
  input         reset, // @[:@20031.4]
  output [31:0] io_rPort_5_output_0, // @[:@20032.4]
  output [31:0] io_rPort_4_output_0, // @[:@20032.4]
  output [31:0] io_rPort_3_output_0, // @[:@20032.4]
  output [31:0] io_rPort_2_output_0, // @[:@20032.4]
  output [31:0] io_rPort_1_output_0, // @[:@20032.4]
  output [31:0] io_rPort_0_output_0, // @[:@20032.4]
  input  [31:0] io_wPort_0_data_0, // @[:@20032.4]
  input         io_wPort_0_reset, // @[:@20032.4]
  input         io_wPort_0_en_0, // @[:@20032.4]
  input         io_sEn_0, // @[:@20032.4]
  input         io_sEn_1, // @[:@20032.4]
  input         io_sEn_2, // @[:@20032.4]
  input         io_sEn_3, // @[:@20032.4]
  input         io_sEn_4, // @[:@20032.4]
  input         io_sEn_5, // @[:@20032.4]
  input         io_sEn_6, // @[:@20032.4]
  input         io_sDone_0, // @[:@20032.4]
  input         io_sDone_1, // @[:@20032.4]
  input         io_sDone_2, // @[:@20032.4]
  input         io_sDone_3, // @[:@20032.4]
  input         io_sDone_4, // @[:@20032.4]
  input         io_sDone_5, // @[:@20032.4]
  input         io_sDone_6 // @[:@20032.4]
);
  wire  nbufFF_clock; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_reset; // @[NBuffers.scala 298:22:@20040.4]
  wire [31:0] nbufFF_io_rPort_5_output_0; // @[NBuffers.scala 298:22:@20040.4]
  wire [31:0] nbufFF_io_rPort_4_output_0; // @[NBuffers.scala 298:22:@20040.4]
  wire [31:0] nbufFF_io_rPort_3_output_0; // @[NBuffers.scala 298:22:@20040.4]
  wire [31:0] nbufFF_io_rPort_2_output_0; // @[NBuffers.scala 298:22:@20040.4]
  wire [31:0] nbufFF_io_rPort_1_output_0; // @[NBuffers.scala 298:22:@20040.4]
  wire [31:0] nbufFF_io_rPort_0_output_0; // @[NBuffers.scala 298:22:@20040.4]
  wire [31:0] nbufFF_io_wPort_0_data_0; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_io_wPort_0_reset; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_io_wPort_0_en_0; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_io_sEn_0; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_io_sEn_1; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_io_sEn_2; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_io_sEn_3; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_io_sEn_4; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_io_sEn_5; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_io_sEn_6; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_io_sDone_0; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_io_sDone_1; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_io_sDone_2; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_io_sDone_3; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_io_sDone_4; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_io_sDone_5; // @[NBuffers.scala 298:22:@20040.4]
  wire  nbufFF_io_sDone_6; // @[NBuffers.scala 298:22:@20040.4]
  NBuf_2 nbufFF ( // @[NBuffers.scala 298:22:@20040.4]
    .clock(nbufFF_clock),
    .reset(nbufFF_reset),
    .io_rPort_5_output_0(nbufFF_io_rPort_5_output_0),
    .io_rPort_4_output_0(nbufFF_io_rPort_4_output_0),
    .io_rPort_3_output_0(nbufFF_io_rPort_3_output_0),
    .io_rPort_2_output_0(nbufFF_io_rPort_2_output_0),
    .io_rPort_1_output_0(nbufFF_io_rPort_1_output_0),
    .io_rPort_0_output_0(nbufFF_io_rPort_0_output_0),
    .io_wPort_0_data_0(nbufFF_io_wPort_0_data_0),
    .io_wPort_0_reset(nbufFF_io_wPort_0_reset),
    .io_wPort_0_en_0(nbufFF_io_wPort_0_en_0),
    .io_sEn_0(nbufFF_io_sEn_0),
    .io_sEn_1(nbufFF_io_sEn_1),
    .io_sEn_2(nbufFF_io_sEn_2),
    .io_sEn_3(nbufFF_io_sEn_3),
    .io_sEn_4(nbufFF_io_sEn_4),
    .io_sEn_5(nbufFF_io_sEn_5),
    .io_sEn_6(nbufFF_io_sEn_6),
    .io_sDone_0(nbufFF_io_sDone_0),
    .io_sDone_1(nbufFF_io_sDone_1),
    .io_sDone_2(nbufFF_io_sDone_2),
    .io_sDone_3(nbufFF_io_sDone_3),
    .io_sDone_4(nbufFF_io_sDone_4),
    .io_sDone_5(nbufFF_io_sDone_5),
    .io_sDone_6(nbufFF_io_sDone_6)
  );
  assign io_rPort_5_output_0 = nbufFF_io_rPort_5_output_0; // @[NBuffers.scala 299:6:@20097.4]
  assign io_rPort_4_output_0 = nbufFF_io_rPort_4_output_0; // @[NBuffers.scala 299:6:@20092.4]
  assign io_rPort_3_output_0 = nbufFF_io_rPort_3_output_0; // @[NBuffers.scala 299:6:@20087.4]
  assign io_rPort_2_output_0 = nbufFF_io_rPort_2_output_0; // @[NBuffers.scala 299:6:@20082.4]
  assign io_rPort_1_output_0 = nbufFF_io_rPort_1_output_0; // @[NBuffers.scala 299:6:@20077.4]
  assign io_rPort_0_output_0 = nbufFF_io_rPort_0_output_0; // @[NBuffers.scala 299:6:@20072.4]
  assign nbufFF_clock = clock; // @[:@20041.4]
  assign nbufFF_reset = reset; // @[:@20042.4]
  assign nbufFF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[NBuffers.scala 299:6:@20069.4]
  assign nbufFF_io_wPort_0_reset = io_wPort_0_reset; // @[NBuffers.scala 299:6:@20068.4]
  assign nbufFF_io_wPort_0_en_0 = io_wPort_0_en_0; // @[NBuffers.scala 299:6:@20065.4]
  assign nbufFF_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 299:6:@20050.4]
  assign nbufFF_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 299:6:@20051.4]
  assign nbufFF_io_sEn_2 = io_sEn_2; // @[NBuffers.scala 299:6:@20052.4]
  assign nbufFF_io_sEn_3 = io_sEn_3; // @[NBuffers.scala 299:6:@20053.4]
  assign nbufFF_io_sEn_4 = io_sEn_4; // @[NBuffers.scala 299:6:@20054.4]
  assign nbufFF_io_sEn_5 = io_sEn_5; // @[NBuffers.scala 299:6:@20055.4]
  assign nbufFF_io_sEn_6 = io_sEn_6; // @[NBuffers.scala 299:6:@20056.4]
  assign nbufFF_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 299:6:@20043.4]
  assign nbufFF_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 299:6:@20044.4]
  assign nbufFF_io_sDone_2 = io_sDone_2; // @[NBuffers.scala 299:6:@20045.4]
  assign nbufFF_io_sDone_3 = io_sDone_3; // @[NBuffers.scala 299:6:@20046.4]
  assign nbufFF_io_sDone_4 = io_sDone_4; // @[NBuffers.scala 299:6:@20047.4]
  assign nbufFF_io_sDone_5 = io_sDone_5; // @[NBuffers.scala 299:6:@20048.4]
  assign nbufFF_io_sDone_6 = io_sDone_6; // @[NBuffers.scala 299:6:@20049.4]
endmodule
module FF_20( // @[:@22537.2]
  input   clock, // @[:@22538.4]
  input   reset, // @[:@22539.4]
  output  io_rPort_4_output_0, // @[:@22540.4]
  output  io_rPort_3_output_0, // @[:@22540.4]
  output  io_rPort_1_output_0, // @[:@22540.4]
  output  io_rPort_0_output_0, // @[:@22540.4]
  input   io_wPort_0_data_0, // @[:@22540.4]
  input   io_wPort_0_reset, // @[:@22540.4]
  input   io_wPort_0_en_0 // @[:@22540.4]
);
  reg  ff; // @[MemPrimitives.scala 321:19:@22580.4]
  reg [31:0] _RAND_0;
  wire  _T_198; // @[MemPrimitives.scala 325:32:@22582.4]
  wire  _T_199; // @[MemPrimitives.scala 325:12:@22583.4]
  assign _T_198 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@22582.4]
  assign _T_199 = io_wPort_0_reset ? 1'h0 : _T_198; // @[MemPrimitives.scala 325:12:@22583.4]
  assign io_rPort_4_output_0 = ff; // @[MemPrimitives.scala 326:34:@22589.4]
  assign io_rPort_3_output_0 = ff; // @[MemPrimitives.scala 326:34:@22588.4]
  assign io_rPort_1_output_0 = ff; // @[MemPrimitives.scala 326:34:@22586.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@22585.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 1'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 1'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module NBuf_3( // @[:@22922.2]
  input   clock, // @[:@22923.4]
  input   reset, // @[:@22924.4]
  output  io_rPort_4_output_0, // @[:@22925.4]
  output  io_rPort_3_output_0, // @[:@22925.4]
  output  io_rPort_1_output_0, // @[:@22925.4]
  output  io_rPort_0_output_0, // @[:@22925.4]
  input   io_wPort_0_data_0, // @[:@22925.4]
  input   io_wPort_0_reset, // @[:@22925.4]
  input   io_wPort_0_en_0, // @[:@22925.4]
  input   io_sEn_0, // @[:@22925.4]
  input   io_sEn_1, // @[:@22925.4]
  input   io_sEn_2, // @[:@22925.4]
  input   io_sEn_3, // @[:@22925.4]
  input   io_sEn_4, // @[:@22925.4]
  input   io_sEn_5, // @[:@22925.4]
  input   io_sEn_6, // @[:@22925.4]
  input   io_sDone_0, // @[:@22925.4]
  input   io_sDone_1, // @[:@22925.4]
  input   io_sDone_2, // @[:@22925.4]
  input   io_sDone_3, // @[:@22925.4]
  input   io_sDone_4, // @[:@22925.4]
  input   io_sDone_5, // @[:@22925.4]
  input   io_sDone_6 // @[:@22925.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@22933.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@22933.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@22933.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@22933.4]
  wire  ctrl_io_sEn_2; // @[NBuffers.scala 83:20:@22933.4]
  wire  ctrl_io_sEn_3; // @[NBuffers.scala 83:20:@22933.4]
  wire  ctrl_io_sEn_4; // @[NBuffers.scala 83:20:@22933.4]
  wire  ctrl_io_sEn_5; // @[NBuffers.scala 83:20:@22933.4]
  wire  ctrl_io_sEn_6; // @[NBuffers.scala 83:20:@22933.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@22933.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@22933.4]
  wire  ctrl_io_sDone_2; // @[NBuffers.scala 83:20:@22933.4]
  wire  ctrl_io_sDone_3; // @[NBuffers.scala 83:20:@22933.4]
  wire  ctrl_io_sDone_4; // @[NBuffers.scala 83:20:@22933.4]
  wire  ctrl_io_sDone_5; // @[NBuffers.scala 83:20:@22933.4]
  wire  ctrl_io_sDone_6; // @[NBuffers.scala 83:20:@22933.4]
  wire [3:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@22933.4]
  wire [3:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@22933.4]
  wire [3:0] ctrl_io_statesInR_2; // @[NBuffers.scala 83:20:@22933.4]
  wire [3:0] ctrl_io_statesInR_3; // @[NBuffers.scala 83:20:@22933.4]
  wire [3:0] ctrl_io_statesInR_4; // @[NBuffers.scala 83:20:@22933.4]
  wire [3:0] ctrl_io_statesInR_5; // @[NBuffers.scala 83:20:@22933.4]
  wire [3:0] ctrl_io_statesInR_6; // @[NBuffers.scala 83:20:@22933.4]
  wire  FF_clock; // @[NBuffers.scala 146:23:@22950.4]
  wire  FF_reset; // @[NBuffers.scala 146:23:@22950.4]
  wire  FF_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@22950.4]
  wire  FF_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@22950.4]
  wire  FF_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@22950.4]
  wire  FF_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@22950.4]
  wire  FF_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@22950.4]
  wire  FF_io_wPort_0_reset; // @[NBuffers.scala 146:23:@22950.4]
  wire  FF_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@22950.4]
  wire  FF_1_clock; // @[NBuffers.scala 146:23:@22991.4]
  wire  FF_1_reset; // @[NBuffers.scala 146:23:@22991.4]
  wire  FF_1_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@22991.4]
  wire  FF_1_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@22991.4]
  wire  FF_1_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@22991.4]
  wire  FF_1_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@22991.4]
  wire  FF_1_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@22991.4]
  wire  FF_1_io_wPort_0_reset; // @[NBuffers.scala 146:23:@22991.4]
  wire  FF_1_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@22991.4]
  wire  FF_2_clock; // @[NBuffers.scala 146:23:@23032.4]
  wire  FF_2_reset; // @[NBuffers.scala 146:23:@23032.4]
  wire  FF_2_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@23032.4]
  wire  FF_2_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@23032.4]
  wire  FF_2_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@23032.4]
  wire  FF_2_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@23032.4]
  wire  FF_2_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@23032.4]
  wire  FF_2_io_wPort_0_reset; // @[NBuffers.scala 146:23:@23032.4]
  wire  FF_2_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@23032.4]
  wire  FF_3_clock; // @[NBuffers.scala 146:23:@23073.4]
  wire  FF_3_reset; // @[NBuffers.scala 146:23:@23073.4]
  wire  FF_3_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@23073.4]
  wire  FF_3_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@23073.4]
  wire  FF_3_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@23073.4]
  wire  FF_3_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@23073.4]
  wire  FF_3_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@23073.4]
  wire  FF_3_io_wPort_0_reset; // @[NBuffers.scala 146:23:@23073.4]
  wire  FF_3_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@23073.4]
  wire  FF_4_clock; // @[NBuffers.scala 146:23:@23114.4]
  wire  FF_4_reset; // @[NBuffers.scala 146:23:@23114.4]
  wire  FF_4_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@23114.4]
  wire  FF_4_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@23114.4]
  wire  FF_4_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@23114.4]
  wire  FF_4_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@23114.4]
  wire  FF_4_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@23114.4]
  wire  FF_4_io_wPort_0_reset; // @[NBuffers.scala 146:23:@23114.4]
  wire  FF_4_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@23114.4]
  wire  FF_5_clock; // @[NBuffers.scala 146:23:@23155.4]
  wire  FF_5_reset; // @[NBuffers.scala 146:23:@23155.4]
  wire  FF_5_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@23155.4]
  wire  FF_5_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@23155.4]
  wire  FF_5_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@23155.4]
  wire  FF_5_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@23155.4]
  wire  FF_5_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@23155.4]
  wire  FF_5_io_wPort_0_reset; // @[NBuffers.scala 146:23:@23155.4]
  wire  FF_5_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@23155.4]
  wire  FF_6_clock; // @[NBuffers.scala 146:23:@23196.4]
  wire  FF_6_reset; // @[NBuffers.scala 146:23:@23196.4]
  wire  FF_6_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@23196.4]
  wire  FF_6_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@23196.4]
  wire  FF_6_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@23196.4]
  wire  FF_6_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@23196.4]
  wire  FF_6_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@23196.4]
  wire  FF_6_io_wPort_0_reset; // @[NBuffers.scala 146:23:@23196.4]
  wire  FF_6_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@23196.4]
  wire  _T_236; // @[NBuffers.scala 153:105:@23244.4]
  wire  _T_240; // @[NBuffers.scala 157:92:@23254.4]
  wire  _T_243; // @[NBuffers.scala 157:92:@23260.4]
  wire  _T_249; // @[NBuffers.scala 157:92:@23272.4]
  wire  _T_252; // @[NBuffers.scala 157:92:@23278.4]
  wire  _T_258; // @[NBuffers.scala 153:105:@23290.4]
  wire  _T_262; // @[NBuffers.scala 157:92:@23300.4]
  wire  _T_265; // @[NBuffers.scala 157:92:@23306.4]
  wire  _T_271; // @[NBuffers.scala 157:92:@23318.4]
  wire  _T_274; // @[NBuffers.scala 157:92:@23324.4]
  wire  _T_280; // @[NBuffers.scala 153:105:@23336.4]
  wire  _T_284; // @[NBuffers.scala 157:92:@23346.4]
  wire  _T_287; // @[NBuffers.scala 157:92:@23352.4]
  wire  _T_293; // @[NBuffers.scala 157:92:@23364.4]
  wire  _T_296; // @[NBuffers.scala 157:92:@23370.4]
  wire  _T_302; // @[NBuffers.scala 153:105:@23382.4]
  wire  _T_306; // @[NBuffers.scala 157:92:@23392.4]
  wire  _T_309; // @[NBuffers.scala 157:92:@23398.4]
  wire  _T_315; // @[NBuffers.scala 157:92:@23410.4]
  wire  _T_318; // @[NBuffers.scala 157:92:@23416.4]
  wire  _T_324; // @[NBuffers.scala 153:105:@23428.4]
  wire  _T_328; // @[NBuffers.scala 157:92:@23438.4]
  wire  _T_331; // @[NBuffers.scala 157:92:@23444.4]
  wire  _T_337; // @[NBuffers.scala 157:92:@23456.4]
  wire  _T_340; // @[NBuffers.scala 157:92:@23462.4]
  wire  _T_346; // @[NBuffers.scala 153:105:@23474.4]
  wire  _T_350; // @[NBuffers.scala 157:92:@23484.4]
  wire  _T_353; // @[NBuffers.scala 157:92:@23490.4]
  wire  _T_359; // @[NBuffers.scala 157:92:@23502.4]
  wire  _T_362; // @[NBuffers.scala 157:92:@23508.4]
  wire  _T_368; // @[NBuffers.scala 153:105:@23520.4]
  wire  _T_372; // @[NBuffers.scala 157:92:@23530.4]
  wire  _T_375; // @[NBuffers.scala 157:92:@23536.4]
  wire  _T_381; // @[NBuffers.scala 157:92:@23548.4]
  wire  _T_384; // @[NBuffers.scala 157:92:@23554.4]
  wire  _T_405; // @[Mux.scala 19:72:@23573.4]
  wire  _T_407; // @[Mux.scala 19:72:@23574.4]
  wire  _T_409; // @[Mux.scala 19:72:@23575.4]
  wire  _T_411; // @[Mux.scala 19:72:@23576.4]
  wire  _T_413; // @[Mux.scala 19:72:@23577.4]
  wire  _T_415; // @[Mux.scala 19:72:@23578.4]
  wire  _T_417; // @[Mux.scala 19:72:@23579.4]
  wire  _T_418; // @[Mux.scala 19:72:@23580.4]
  wire  _T_419; // @[Mux.scala 19:72:@23581.4]
  wire  _T_420; // @[Mux.scala 19:72:@23582.4]
  wire  _T_421; // @[Mux.scala 19:72:@23583.4]
  wire  _T_422; // @[Mux.scala 19:72:@23584.4]
  wire  _T_442; // @[Mux.scala 19:72:@23596.4]
  wire  _T_444; // @[Mux.scala 19:72:@23597.4]
  wire  _T_446; // @[Mux.scala 19:72:@23598.4]
  wire  _T_448; // @[Mux.scala 19:72:@23599.4]
  wire  _T_450; // @[Mux.scala 19:72:@23600.4]
  wire  _T_452; // @[Mux.scala 19:72:@23601.4]
  wire  _T_454; // @[Mux.scala 19:72:@23602.4]
  wire  _T_455; // @[Mux.scala 19:72:@23603.4]
  wire  _T_456; // @[Mux.scala 19:72:@23604.4]
  wire  _T_457; // @[Mux.scala 19:72:@23605.4]
  wire  _T_458; // @[Mux.scala 19:72:@23606.4]
  wire  _T_459; // @[Mux.scala 19:72:@23607.4]
  wire  _T_516; // @[Mux.scala 19:72:@23642.4]
  wire  _T_518; // @[Mux.scala 19:72:@23643.4]
  wire  _T_520; // @[Mux.scala 19:72:@23644.4]
  wire  _T_522; // @[Mux.scala 19:72:@23645.4]
  wire  _T_524; // @[Mux.scala 19:72:@23646.4]
  wire  _T_526; // @[Mux.scala 19:72:@23647.4]
  wire  _T_528; // @[Mux.scala 19:72:@23648.4]
  wire  _T_529; // @[Mux.scala 19:72:@23649.4]
  wire  _T_530; // @[Mux.scala 19:72:@23650.4]
  wire  _T_531; // @[Mux.scala 19:72:@23651.4]
  wire  _T_532; // @[Mux.scala 19:72:@23652.4]
  wire  _T_533; // @[Mux.scala 19:72:@23653.4]
  wire  _T_553; // @[Mux.scala 19:72:@23665.4]
  wire  _T_555; // @[Mux.scala 19:72:@23666.4]
  wire  _T_557; // @[Mux.scala 19:72:@23667.4]
  wire  _T_559; // @[Mux.scala 19:72:@23668.4]
  wire  _T_561; // @[Mux.scala 19:72:@23669.4]
  wire  _T_563; // @[Mux.scala 19:72:@23670.4]
  wire  _T_565; // @[Mux.scala 19:72:@23671.4]
  wire  _T_566; // @[Mux.scala 19:72:@23672.4]
  wire  _T_567; // @[Mux.scala 19:72:@23673.4]
  wire  _T_568; // @[Mux.scala 19:72:@23674.4]
  wire  _T_569; // @[Mux.scala 19:72:@23675.4]
  wire  _T_570; // @[Mux.scala 19:72:@23676.4]
  NBufController_3 ctrl ( // @[NBuffers.scala 83:20:@22933.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sEn_2(ctrl_io_sEn_2),
    .io_sEn_3(ctrl_io_sEn_3),
    .io_sEn_4(ctrl_io_sEn_4),
    .io_sEn_5(ctrl_io_sEn_5),
    .io_sEn_6(ctrl_io_sEn_6),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_sDone_2(ctrl_io_sDone_2),
    .io_sDone_3(ctrl_io_sDone_3),
    .io_sDone_4(ctrl_io_sDone_4),
    .io_sDone_5(ctrl_io_sDone_5),
    .io_sDone_6(ctrl_io_sDone_6),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1),
    .io_statesInR_2(ctrl_io_statesInR_2),
    .io_statesInR_3(ctrl_io_statesInR_3),
    .io_statesInR_4(ctrl_io_statesInR_4),
    .io_statesInR_5(ctrl_io_statesInR_5),
    .io_statesInR_6(ctrl_io_statesInR_6)
  );
  FF_20 FF ( // @[NBuffers.scala 146:23:@22950.4]
    .clock(FF_clock),
    .reset(FF_reset),
    .io_rPort_4_output_0(FF_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_io_rPort_3_output_0),
    .io_rPort_1_output_0(FF_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_io_wPort_0_en_0)
  );
  FF_20 FF_1 ( // @[NBuffers.scala 146:23:@22991.4]
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_rPort_4_output_0(FF_1_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_1_io_rPort_3_output_0),
    .io_rPort_1_output_0(FF_1_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_1_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_1_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_1_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_1_io_wPort_0_en_0)
  );
  FF_20 FF_2 ( // @[NBuffers.scala 146:23:@23032.4]
    .clock(FF_2_clock),
    .reset(FF_2_reset),
    .io_rPort_4_output_0(FF_2_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_2_io_rPort_3_output_0),
    .io_rPort_1_output_0(FF_2_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_2_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_2_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_2_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_2_io_wPort_0_en_0)
  );
  FF_20 FF_3 ( // @[NBuffers.scala 146:23:@23073.4]
    .clock(FF_3_clock),
    .reset(FF_3_reset),
    .io_rPort_4_output_0(FF_3_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_3_io_rPort_3_output_0),
    .io_rPort_1_output_0(FF_3_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_3_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_3_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_3_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_3_io_wPort_0_en_0)
  );
  FF_20 FF_4 ( // @[NBuffers.scala 146:23:@23114.4]
    .clock(FF_4_clock),
    .reset(FF_4_reset),
    .io_rPort_4_output_0(FF_4_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_4_io_rPort_3_output_0),
    .io_rPort_1_output_0(FF_4_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_4_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_4_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_4_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_4_io_wPort_0_en_0)
  );
  FF_20 FF_5 ( // @[NBuffers.scala 146:23:@23155.4]
    .clock(FF_5_clock),
    .reset(FF_5_reset),
    .io_rPort_4_output_0(FF_5_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_5_io_rPort_3_output_0),
    .io_rPort_1_output_0(FF_5_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_5_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_5_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_5_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_5_io_wPort_0_en_0)
  );
  FF_20 FF_6 ( // @[NBuffers.scala 146:23:@23196.4]
    .clock(FF_6_clock),
    .reset(FF_6_reset),
    .io_rPort_4_output_0(FF_6_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_6_io_rPort_3_output_0),
    .io_rPort_1_output_0(FF_6_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_6_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_6_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_6_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_6_io_wPort_0_en_0)
  );
  assign _T_236 = ctrl_io_statesInW_0 == 4'h0; // @[NBuffers.scala 153:105:@23244.4]
  assign _T_240 = ctrl_io_statesInR_1 == 4'h0; // @[NBuffers.scala 157:92:@23254.4]
  assign _T_243 = ctrl_io_statesInR_2 == 4'h0; // @[NBuffers.scala 157:92:@23260.4]
  assign _T_249 = ctrl_io_statesInR_4 == 4'h0; // @[NBuffers.scala 157:92:@23272.4]
  assign _T_252 = ctrl_io_statesInR_5 == 4'h0; // @[NBuffers.scala 157:92:@23278.4]
  assign _T_258 = ctrl_io_statesInW_0 == 4'h1; // @[NBuffers.scala 153:105:@23290.4]
  assign _T_262 = ctrl_io_statesInR_1 == 4'h1; // @[NBuffers.scala 157:92:@23300.4]
  assign _T_265 = ctrl_io_statesInR_2 == 4'h1; // @[NBuffers.scala 157:92:@23306.4]
  assign _T_271 = ctrl_io_statesInR_4 == 4'h1; // @[NBuffers.scala 157:92:@23318.4]
  assign _T_274 = ctrl_io_statesInR_5 == 4'h1; // @[NBuffers.scala 157:92:@23324.4]
  assign _T_280 = ctrl_io_statesInW_0 == 4'h2; // @[NBuffers.scala 153:105:@23336.4]
  assign _T_284 = ctrl_io_statesInR_1 == 4'h2; // @[NBuffers.scala 157:92:@23346.4]
  assign _T_287 = ctrl_io_statesInR_2 == 4'h2; // @[NBuffers.scala 157:92:@23352.4]
  assign _T_293 = ctrl_io_statesInR_4 == 4'h2; // @[NBuffers.scala 157:92:@23364.4]
  assign _T_296 = ctrl_io_statesInR_5 == 4'h2; // @[NBuffers.scala 157:92:@23370.4]
  assign _T_302 = ctrl_io_statesInW_0 == 4'h3; // @[NBuffers.scala 153:105:@23382.4]
  assign _T_306 = ctrl_io_statesInR_1 == 4'h3; // @[NBuffers.scala 157:92:@23392.4]
  assign _T_309 = ctrl_io_statesInR_2 == 4'h3; // @[NBuffers.scala 157:92:@23398.4]
  assign _T_315 = ctrl_io_statesInR_4 == 4'h3; // @[NBuffers.scala 157:92:@23410.4]
  assign _T_318 = ctrl_io_statesInR_5 == 4'h3; // @[NBuffers.scala 157:92:@23416.4]
  assign _T_324 = ctrl_io_statesInW_0 == 4'h4; // @[NBuffers.scala 153:105:@23428.4]
  assign _T_328 = ctrl_io_statesInR_1 == 4'h4; // @[NBuffers.scala 157:92:@23438.4]
  assign _T_331 = ctrl_io_statesInR_2 == 4'h4; // @[NBuffers.scala 157:92:@23444.4]
  assign _T_337 = ctrl_io_statesInR_4 == 4'h4; // @[NBuffers.scala 157:92:@23456.4]
  assign _T_340 = ctrl_io_statesInR_5 == 4'h4; // @[NBuffers.scala 157:92:@23462.4]
  assign _T_346 = ctrl_io_statesInW_0 == 4'h5; // @[NBuffers.scala 153:105:@23474.4]
  assign _T_350 = ctrl_io_statesInR_1 == 4'h5; // @[NBuffers.scala 157:92:@23484.4]
  assign _T_353 = ctrl_io_statesInR_2 == 4'h5; // @[NBuffers.scala 157:92:@23490.4]
  assign _T_359 = ctrl_io_statesInR_4 == 4'h5; // @[NBuffers.scala 157:92:@23502.4]
  assign _T_362 = ctrl_io_statesInR_5 == 4'h5; // @[NBuffers.scala 157:92:@23508.4]
  assign _T_368 = ctrl_io_statesInW_0 == 4'h6; // @[NBuffers.scala 153:105:@23520.4]
  assign _T_372 = ctrl_io_statesInR_1 == 4'h6; // @[NBuffers.scala 157:92:@23530.4]
  assign _T_375 = ctrl_io_statesInR_2 == 4'h6; // @[NBuffers.scala 157:92:@23536.4]
  assign _T_381 = ctrl_io_statesInR_4 == 4'h6; // @[NBuffers.scala 157:92:@23548.4]
  assign _T_384 = ctrl_io_statesInR_5 == 4'h6; // @[NBuffers.scala 157:92:@23554.4]
  assign _T_405 = _T_240 ? FF_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@23573.4]
  assign _T_407 = _T_262 ? FF_1_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@23574.4]
  assign _T_409 = _T_284 ? FF_2_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@23575.4]
  assign _T_411 = _T_306 ? FF_3_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@23576.4]
  assign _T_413 = _T_328 ? FF_4_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@23577.4]
  assign _T_415 = _T_350 ? FF_5_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@23578.4]
  assign _T_417 = _T_372 ? FF_6_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@23579.4]
  assign _T_418 = _T_405 | _T_407; // @[Mux.scala 19:72:@23580.4]
  assign _T_419 = _T_418 | _T_409; // @[Mux.scala 19:72:@23581.4]
  assign _T_420 = _T_419 | _T_411; // @[Mux.scala 19:72:@23582.4]
  assign _T_421 = _T_420 | _T_413; // @[Mux.scala 19:72:@23583.4]
  assign _T_422 = _T_421 | _T_415; // @[Mux.scala 19:72:@23584.4]
  assign _T_442 = _T_243 ? FF_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@23596.4]
  assign _T_444 = _T_265 ? FF_1_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@23597.4]
  assign _T_446 = _T_287 ? FF_2_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@23598.4]
  assign _T_448 = _T_309 ? FF_3_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@23599.4]
  assign _T_450 = _T_331 ? FF_4_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@23600.4]
  assign _T_452 = _T_353 ? FF_5_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@23601.4]
  assign _T_454 = _T_375 ? FF_6_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@23602.4]
  assign _T_455 = _T_442 | _T_444; // @[Mux.scala 19:72:@23603.4]
  assign _T_456 = _T_455 | _T_446; // @[Mux.scala 19:72:@23604.4]
  assign _T_457 = _T_456 | _T_448; // @[Mux.scala 19:72:@23605.4]
  assign _T_458 = _T_457 | _T_450; // @[Mux.scala 19:72:@23606.4]
  assign _T_459 = _T_458 | _T_452; // @[Mux.scala 19:72:@23607.4]
  assign _T_516 = _T_249 ? FF_io_rPort_3_output_0 : 1'h0; // @[Mux.scala 19:72:@23642.4]
  assign _T_518 = _T_271 ? FF_1_io_rPort_3_output_0 : 1'h0; // @[Mux.scala 19:72:@23643.4]
  assign _T_520 = _T_293 ? FF_2_io_rPort_3_output_0 : 1'h0; // @[Mux.scala 19:72:@23644.4]
  assign _T_522 = _T_315 ? FF_3_io_rPort_3_output_0 : 1'h0; // @[Mux.scala 19:72:@23645.4]
  assign _T_524 = _T_337 ? FF_4_io_rPort_3_output_0 : 1'h0; // @[Mux.scala 19:72:@23646.4]
  assign _T_526 = _T_359 ? FF_5_io_rPort_3_output_0 : 1'h0; // @[Mux.scala 19:72:@23647.4]
  assign _T_528 = _T_381 ? FF_6_io_rPort_3_output_0 : 1'h0; // @[Mux.scala 19:72:@23648.4]
  assign _T_529 = _T_516 | _T_518; // @[Mux.scala 19:72:@23649.4]
  assign _T_530 = _T_529 | _T_520; // @[Mux.scala 19:72:@23650.4]
  assign _T_531 = _T_530 | _T_522; // @[Mux.scala 19:72:@23651.4]
  assign _T_532 = _T_531 | _T_524; // @[Mux.scala 19:72:@23652.4]
  assign _T_533 = _T_532 | _T_526; // @[Mux.scala 19:72:@23653.4]
  assign _T_553 = _T_252 ? FF_io_rPort_4_output_0 : 1'h0; // @[Mux.scala 19:72:@23665.4]
  assign _T_555 = _T_274 ? FF_1_io_rPort_4_output_0 : 1'h0; // @[Mux.scala 19:72:@23666.4]
  assign _T_557 = _T_296 ? FF_2_io_rPort_4_output_0 : 1'h0; // @[Mux.scala 19:72:@23667.4]
  assign _T_559 = _T_318 ? FF_3_io_rPort_4_output_0 : 1'h0; // @[Mux.scala 19:72:@23668.4]
  assign _T_561 = _T_340 ? FF_4_io_rPort_4_output_0 : 1'h0; // @[Mux.scala 19:72:@23669.4]
  assign _T_563 = _T_362 ? FF_5_io_rPort_4_output_0 : 1'h0; // @[Mux.scala 19:72:@23670.4]
  assign _T_565 = _T_384 ? FF_6_io_rPort_4_output_0 : 1'h0; // @[Mux.scala 19:72:@23671.4]
  assign _T_566 = _T_553 | _T_555; // @[Mux.scala 19:72:@23672.4]
  assign _T_567 = _T_566 | _T_557; // @[Mux.scala 19:72:@23673.4]
  assign _T_568 = _T_567 | _T_559; // @[Mux.scala 19:72:@23674.4]
  assign _T_569 = _T_568 | _T_561; // @[Mux.scala 19:72:@23675.4]
  assign _T_570 = _T_569 | _T_563; // @[Mux.scala 19:72:@23676.4]
  assign io_rPort_4_output_0 = _T_570 | _T_565; // @[NBuffers.scala 163:66:@23680.4]
  assign io_rPort_3_output_0 = _T_533 | _T_528; // @[NBuffers.scala 163:66:@23657.4]
  assign io_rPort_1_output_0 = _T_459 | _T_454; // @[NBuffers.scala 163:66:@23611.4]
  assign io_rPort_0_output_0 = _T_422 | _T_417; // @[NBuffers.scala 163:66:@23588.4]
  assign ctrl_clock = clock; // @[:@22934.4]
  assign ctrl_reset = reset; // @[:@22935.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@22936.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@22938.4]
  assign ctrl_io_sEn_2 = io_sEn_2; // @[NBuffers.scala 85:20:@22940.4]
  assign ctrl_io_sEn_3 = io_sEn_3; // @[NBuffers.scala 85:20:@22942.4]
  assign ctrl_io_sEn_4 = io_sEn_4; // @[NBuffers.scala 85:20:@22944.4]
  assign ctrl_io_sEn_5 = io_sEn_5; // @[NBuffers.scala 85:20:@22946.4]
  assign ctrl_io_sEn_6 = io_sEn_6; // @[NBuffers.scala 85:20:@22948.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@22937.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@22939.4]
  assign ctrl_io_sDone_2 = io_sDone_2; // @[NBuffers.scala 86:22:@22941.4]
  assign ctrl_io_sDone_3 = io_sDone_3; // @[NBuffers.scala 86:22:@22943.4]
  assign ctrl_io_sDone_4 = io_sDone_4; // @[NBuffers.scala 86:22:@22945.4]
  assign ctrl_io_sDone_5 = io_sDone_5; // @[NBuffers.scala 86:22:@22947.4]
  assign ctrl_io_sDone_6 = io_sDone_6; // @[NBuffers.scala 86:22:@22949.4]
  assign FF_clock = clock; // @[:@22951.4]
  assign FF_reset = reset; // @[:@22952.4]
  assign FF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@23247.4]
  assign FF_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@23248.4]
  assign FF_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_236; // @[MemPrimitives.scala 37:29:@23253.4]
  assign FF_1_clock = clock; // @[:@22992.4]
  assign FF_1_reset = reset; // @[:@22993.4]
  assign FF_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@23293.4]
  assign FF_1_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@23294.4]
  assign FF_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_258; // @[MemPrimitives.scala 37:29:@23299.4]
  assign FF_2_clock = clock; // @[:@23033.4]
  assign FF_2_reset = reset; // @[:@23034.4]
  assign FF_2_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@23339.4]
  assign FF_2_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@23340.4]
  assign FF_2_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_280; // @[MemPrimitives.scala 37:29:@23345.4]
  assign FF_3_clock = clock; // @[:@23074.4]
  assign FF_3_reset = reset; // @[:@23075.4]
  assign FF_3_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@23385.4]
  assign FF_3_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@23386.4]
  assign FF_3_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_302; // @[MemPrimitives.scala 37:29:@23391.4]
  assign FF_4_clock = clock; // @[:@23115.4]
  assign FF_4_reset = reset; // @[:@23116.4]
  assign FF_4_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@23431.4]
  assign FF_4_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@23432.4]
  assign FF_4_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_324; // @[MemPrimitives.scala 37:29:@23437.4]
  assign FF_5_clock = clock; // @[:@23156.4]
  assign FF_5_reset = reset; // @[:@23157.4]
  assign FF_5_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@23477.4]
  assign FF_5_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@23478.4]
  assign FF_5_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_346; // @[MemPrimitives.scala 37:29:@23483.4]
  assign FF_6_clock = clock; // @[:@23197.4]
  assign FF_6_reset = reset; // @[:@23198.4]
  assign FF_6_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@23523.4]
  assign FF_6_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@23524.4]
  assign FF_6_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_368; // @[MemPrimitives.scala 37:29:@23529.4]
endmodule
module b552_chain( // @[:@23705.2]
  input   clock, // @[:@23706.4]
  input   reset, // @[:@23707.4]
  output  io_rPort_4_output_0, // @[:@23708.4]
  output  io_rPort_3_output_0, // @[:@23708.4]
  output  io_rPort_1_output_0, // @[:@23708.4]
  output  io_rPort_0_output_0, // @[:@23708.4]
  input   io_wPort_0_data_0, // @[:@23708.4]
  input   io_wPort_0_reset, // @[:@23708.4]
  input   io_wPort_0_en_0, // @[:@23708.4]
  input   io_sEn_0, // @[:@23708.4]
  input   io_sEn_1, // @[:@23708.4]
  input   io_sEn_2, // @[:@23708.4]
  input   io_sEn_3, // @[:@23708.4]
  input   io_sEn_4, // @[:@23708.4]
  input   io_sEn_5, // @[:@23708.4]
  input   io_sEn_6, // @[:@23708.4]
  input   io_sDone_0, // @[:@23708.4]
  input   io_sDone_1, // @[:@23708.4]
  input   io_sDone_2, // @[:@23708.4]
  input   io_sDone_3, // @[:@23708.4]
  input   io_sDone_4, // @[:@23708.4]
  input   io_sDone_5, // @[:@23708.4]
  input   io_sDone_6 // @[:@23708.4]
);
  wire  nbufFF_clock; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_reset; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_rPort_4_output_0; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_rPort_3_output_0; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_rPort_1_output_0; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_rPort_0_output_0; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_wPort_0_data_0; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_wPort_0_reset; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_wPort_0_en_0; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_sEn_0; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_sEn_1; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_sEn_2; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_sEn_3; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_sEn_4; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_sEn_5; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_sEn_6; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_sDone_0; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_sDone_1; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_sDone_2; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_sDone_3; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_sDone_4; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_sDone_5; // @[NBuffers.scala 298:22:@23716.4]
  wire  nbufFF_io_sDone_6; // @[NBuffers.scala 298:22:@23716.4]
  NBuf_3 nbufFF ( // @[NBuffers.scala 298:22:@23716.4]
    .clock(nbufFF_clock),
    .reset(nbufFF_reset),
    .io_rPort_4_output_0(nbufFF_io_rPort_4_output_0),
    .io_rPort_3_output_0(nbufFF_io_rPort_3_output_0),
    .io_rPort_1_output_0(nbufFF_io_rPort_1_output_0),
    .io_rPort_0_output_0(nbufFF_io_rPort_0_output_0),
    .io_wPort_0_data_0(nbufFF_io_wPort_0_data_0),
    .io_wPort_0_reset(nbufFF_io_wPort_0_reset),
    .io_wPort_0_en_0(nbufFF_io_wPort_0_en_0),
    .io_sEn_0(nbufFF_io_sEn_0),
    .io_sEn_1(nbufFF_io_sEn_1),
    .io_sEn_2(nbufFF_io_sEn_2),
    .io_sEn_3(nbufFF_io_sEn_3),
    .io_sEn_4(nbufFF_io_sEn_4),
    .io_sEn_5(nbufFF_io_sEn_5),
    .io_sEn_6(nbufFF_io_sEn_6),
    .io_sDone_0(nbufFF_io_sDone_0),
    .io_sDone_1(nbufFF_io_sDone_1),
    .io_sDone_2(nbufFF_io_sDone_2),
    .io_sDone_3(nbufFF_io_sDone_3),
    .io_sDone_4(nbufFF_io_sDone_4),
    .io_sDone_5(nbufFF_io_sDone_5),
    .io_sDone_6(nbufFF_io_sDone_6)
  );
  assign io_rPort_4_output_0 = nbufFF_io_rPort_4_output_0; // @[NBuffers.scala 299:6:@23768.4]
  assign io_rPort_3_output_0 = nbufFF_io_rPort_3_output_0; // @[NBuffers.scala 299:6:@23763.4]
  assign io_rPort_1_output_0 = nbufFF_io_rPort_1_output_0; // @[NBuffers.scala 299:6:@23753.4]
  assign io_rPort_0_output_0 = nbufFF_io_rPort_0_output_0; // @[NBuffers.scala 299:6:@23748.4]
  assign nbufFF_clock = clock; // @[:@23717.4]
  assign nbufFF_reset = reset; // @[:@23718.4]
  assign nbufFF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[NBuffers.scala 299:6:@23745.4]
  assign nbufFF_io_wPort_0_reset = io_wPort_0_reset; // @[NBuffers.scala 299:6:@23744.4]
  assign nbufFF_io_wPort_0_en_0 = io_wPort_0_en_0; // @[NBuffers.scala 299:6:@23741.4]
  assign nbufFF_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 299:6:@23726.4]
  assign nbufFF_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 299:6:@23727.4]
  assign nbufFF_io_sEn_2 = io_sEn_2; // @[NBuffers.scala 299:6:@23728.4]
  assign nbufFF_io_sEn_3 = io_sEn_3; // @[NBuffers.scala 299:6:@23729.4]
  assign nbufFF_io_sEn_4 = io_sEn_4; // @[NBuffers.scala 299:6:@23730.4]
  assign nbufFF_io_sEn_5 = io_sEn_5; // @[NBuffers.scala 299:6:@23731.4]
  assign nbufFF_io_sEn_6 = io_sEn_6; // @[NBuffers.scala 299:6:@23732.4]
  assign nbufFF_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 299:6:@23719.4]
  assign nbufFF_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 299:6:@23720.4]
  assign nbufFF_io_sDone_2 = io_sDone_2; // @[NBuffers.scala 299:6:@23721.4]
  assign nbufFF_io_sDone_3 = io_sDone_3; // @[NBuffers.scala 299:6:@23722.4]
  assign nbufFF_io_sDone_4 = io_sDone_4; // @[NBuffers.scala 299:6:@23723.4]
  assign nbufFF_io_sDone_5 = io_sDone_5; // @[NBuffers.scala 299:6:@23724.4]
  assign nbufFF_io_sDone_6 = io_sDone_6; // @[NBuffers.scala 299:6:@23725.4]
endmodule
module RetimeWrapper_249( // @[:@24747.2]
  input         clock, // @[:@24748.4]
  input         reset, // @[:@24749.4]
  input         io_flow, // @[:@24750.4]
  input  [31:0] io_in, // @[:@24750.4]
  output [31:0] io_out // @[:@24750.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@24752.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@24752.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@24752.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@24752.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@24752.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@24752.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@24752.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24765.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24764.4]
  assign sr_init = 32'h5; // @[RetimeShiftRegister.scala 19:16:@24763.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24762.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24761.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@24759.4]
endmodule
module NBufCtr_25( // @[:@24767.2]
  input         clock, // @[:@24768.4]
  input         reset, // @[:@24769.4]
  input         io_input_countUp, // @[:@24770.4]
  input         io_input_enable, // @[:@24770.4]
  output [31:0] io_output_count // @[:@24770.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@24807.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@24807.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@24807.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@24812.4 package.scala 96:25:@24813.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@24773.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@24774.4]
  wire  _T_21; // @[Counter.scala 49:55:@24775.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@24776.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@24777.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@24778.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@24779.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@24780.4]
  wire  _T_33; // @[Counter.scala 51:52:@24784.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@24785.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@24786.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@24787.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@24788.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@24789.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@24790.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@24791.4]
  wire  _T_45; // @[Counter.scala 52:70:@24792.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@24794.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@24795.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@24796.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@24797.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@24798.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@24799.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@24802.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@24803.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@24805.4]
  RetimeWrapper_249 RetimeWrapper ( // @[package.scala 93:22:@24807.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@24812.4 package.scala 96:25:@24813.4]
  assign _T_18 = {{1'd0}, _T_66}; // @[Counter.scala 49:32:@24773.4]
  assign _T_19 = _T_18[31:0]; // @[Counter.scala 49:32:@24774.4]
  assign _T_21 = _T_19 >= 32'h6; // @[Counter.scala 49:55:@24775.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@24776.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 49:91:@24777.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 49:91:@24778.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@24779.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@24780.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@24784.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@24785.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@24786.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@24787.4]
  assign _T_39 = _T_33 ? 32'h5 : _T_38; // @[Counter.scala 51:47:@24788.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@24789.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@24790.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@24791.4]
  assign _T_45 = _T_43 >= 32'h6; // @[Counter.scala 52:70:@24792.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@24794.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@24795.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@24796.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@24797.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@24798.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@24799.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@24802.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@24803.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@24805.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@24815.4]
  assign RetimeWrapper_clock = clock; // @[:@24808.4]
  assign RetimeWrapper_reset = reset; // @[:@24809.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@24811.4]
  assign RetimeWrapper_io_in = reset ? 32'h5 : _T_62; // @[package.scala 94:16:@24810.4]
endmodule
module NBufCtr_26( // @[:@24849.2]
  input         clock, // @[:@24850.4]
  input         reset, // @[:@24851.4]
  input         io_input_countUp, // @[:@24852.4]
  input         io_input_enable, // @[:@24852.4]
  output [31:0] io_output_count // @[:@24852.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@24889.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@24889.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@24889.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@24889.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@24889.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@24894.4 package.scala 96:25:@24895.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@24855.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@24856.4]
  wire  _T_21; // @[Counter.scala 49:55:@24857.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@24858.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@24859.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@24860.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@24861.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@24862.4]
  wire  _T_33; // @[Counter.scala 51:52:@24866.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@24867.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@24868.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@24869.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@24870.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@24871.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@24872.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@24873.4]
  wire  _T_45; // @[Counter.scala 52:70:@24874.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@24876.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@24877.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@24878.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@24879.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@24880.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@24881.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@24884.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@24885.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@24887.4]
  RetimeWrapper_249 RetimeWrapper ( // @[package.scala 93:22:@24889.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@24894.4 package.scala 96:25:@24895.4]
  assign _T_18 = _T_66 + 32'h5; // @[Counter.scala 49:32:@24855.4]
  assign _T_19 = _T_66 + 32'h5; // @[Counter.scala 49:32:@24856.4]
  assign _T_21 = _T_19 >= 32'h6; // @[Counter.scala 49:55:@24857.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@24858.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 49:91:@24859.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 49:91:@24860.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@24861.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@24862.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@24866.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@24867.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@24868.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@24869.4]
  assign _T_39 = _T_33 ? 32'h5 : _T_38; // @[Counter.scala 51:47:@24870.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@24871.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@24872.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@24873.4]
  assign _T_45 = _T_43 >= 32'h6; // @[Counter.scala 52:70:@24874.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@24876.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@24877.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@24878.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@24879.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@24880.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@24881.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@24884.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@24885.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@24887.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@24897.4]
  assign RetimeWrapper_clock = clock; // @[:@24890.4]
  assign RetimeWrapper_reset = reset; // @[:@24891.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@24893.4]
  assign RetimeWrapper_io_in = reset ? 32'h5 : _T_62; // @[package.scala 94:16:@24892.4]
endmodule
module NBufCtr_28( // @[:@25013.2]
  input         clock, // @[:@25014.4]
  input         reset, // @[:@25015.4]
  input         io_input_countUp, // @[:@25016.4]
  input         io_input_enable, // @[:@25016.4]
  output [31:0] io_output_count // @[:@25016.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@25053.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@25053.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@25053.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@25053.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@25053.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@25058.4 package.scala 96:25:@25059.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@25019.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@25020.4]
  wire  _T_21; // @[Counter.scala 49:55:@25021.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@25022.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@25023.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@25024.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@25025.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@25026.4]
  wire  _T_33; // @[Counter.scala 51:52:@25030.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@25031.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@25032.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@25033.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@25034.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@25035.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@25044.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@25045.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@25048.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@25049.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@25051.4]
  RetimeWrapper_249 RetimeWrapper ( // @[package.scala 93:22:@25053.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@25058.4 package.scala 96:25:@25059.4]
  assign _T_18 = _T_66 + 32'h1; // @[Counter.scala 49:32:@25019.4]
  assign _T_19 = _T_66 + 32'h1; // @[Counter.scala 49:32:@25020.4]
  assign _T_21 = _T_19 >= 32'h6; // @[Counter.scala 49:55:@25021.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@25022.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 49:91:@25023.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 49:91:@25024.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@25025.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@25026.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@25030.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@25031.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@25032.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@25033.4]
  assign _T_39 = _T_33 ? 32'h5 : _T_38; // @[Counter.scala 51:47:@25034.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@25035.4]
  assign _T_53 = {{1'd0}, _T_27}; // @[Counter.scala 52:107:@25044.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@25045.4]
  assign _T_58 = _T_21 ? _T_54 : _T_19; // @[Counter.scala 52:45:@25048.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@25049.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@25051.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@25061.4]
  assign RetimeWrapper_clock = clock; // @[:@25054.4]
  assign RetimeWrapper_reset = reset; // @[:@25055.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@25057.4]
  assign RetimeWrapper_io_in = reset ? 32'h5 : _T_62; // @[package.scala 94:16:@25056.4]
endmodule
module NBufCtr_29( // @[:@25095.2]
  input   clock, // @[:@25096.4]
  input   reset, // @[:@25097.4]
  input   io_input_countUp, // @[:@25098.4]
  input   io_input_enable // @[:@25098.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@25135.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@25135.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@25135.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@25135.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@25135.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@25140.4 package.scala 96:25:@25141.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@25104.4]
  wire  _T_33; // @[Counter.scala 51:52:@25112.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@25113.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@25114.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@25115.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@25116.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@25117.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@25118.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@25119.4]
  wire  _T_45; // @[Counter.scala 52:70:@25120.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@25122.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@25123.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@25124.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@25125.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@25126.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@25127.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@25130.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@25131.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@25133.4]
  RetimeWrapper_249 RetimeWrapper ( // @[package.scala 93:22:@25135.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@25140.4 package.scala 96:25:@25141.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@25104.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@25112.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@25113.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@25114.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@25115.4]
  assign _T_39 = _T_33 ? 32'h5 : _T_38; // @[Counter.scala 51:47:@25116.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@25117.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@25118.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@25119.4]
  assign _T_45 = _T_43 >= 32'h6; // @[Counter.scala 52:70:@25120.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@25122.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@25123.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@25124.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@25125.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@25126.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@25127.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@25130.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@25131.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@25133.4]
  assign RetimeWrapper_clock = clock; // @[:@25136.4]
  assign RetimeWrapper_reset = reset; // @[:@25137.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@25139.4]
  assign RetimeWrapper_io_in = reset ? 32'h5 : _T_62; // @[package.scala 94:16:@25138.4]
endmodule
module NBufCtr_30( // @[:@25177.2]
  input   clock, // @[:@25178.4]
  input   reset, // @[:@25179.4]
  input   io_input_countUp, // @[:@25180.4]
  input   io_input_enable // @[:@25180.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@25217.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@25217.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@25217.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@25217.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@25217.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@25222.4 package.scala 96:25:@25223.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@25186.4]
  wire  _T_33; // @[Counter.scala 51:52:@25194.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@25195.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@25196.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@25197.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@25198.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@25199.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@25200.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@25201.4]
  wire  _T_45; // @[Counter.scala 52:70:@25202.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@25204.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@25205.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@25206.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@25207.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@25208.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@25209.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@25212.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@25213.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@25215.4]
  RetimeWrapper_249 RetimeWrapper ( // @[package.scala 93:22:@25217.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@25222.4 package.scala 96:25:@25223.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@25186.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@25194.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@25195.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@25196.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@25197.4]
  assign _T_39 = _T_33 ? 32'h5 : _T_38; // @[Counter.scala 51:47:@25198.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@25199.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@25200.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@25201.4]
  assign _T_45 = _T_43 >= 32'h6; // @[Counter.scala 52:70:@25202.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@25204.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@25205.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@25206.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@25207.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@25208.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@25209.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@25212.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@25213.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@25215.4]
  assign RetimeWrapper_clock = clock; // @[:@25218.4]
  assign RetimeWrapper_reset = reset; // @[:@25219.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@25221.4]
  assign RetimeWrapper_io_in = reset ? 32'h5 : _T_62; // @[package.scala 94:16:@25220.4]
endmodule
module NBufCtr_31( // @[:@25259.2]
  input   clock, // @[:@25260.4]
  input   reset, // @[:@25261.4]
  input   io_input_countUp, // @[:@25262.4]
  input   io_input_enable // @[:@25262.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@25299.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@25299.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@25299.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@25299.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@25299.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@25304.4 package.scala 96:25:@25305.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@25268.4]
  wire  _T_33; // @[Counter.scala 51:52:@25276.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@25277.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@25278.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@25279.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@25280.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@25281.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@25282.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@25283.4]
  wire  _T_45; // @[Counter.scala 52:70:@25284.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@25286.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@25287.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@25288.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@25289.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@25290.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@25291.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@25294.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@25295.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@25297.4]
  RetimeWrapper_249 RetimeWrapper ( // @[package.scala 93:22:@25299.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@25304.4 package.scala 96:25:@25305.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@25268.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@25276.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@25277.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@25278.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@25279.4]
  assign _T_39 = _T_33 ? 32'h5 : _T_38; // @[Counter.scala 51:47:@25280.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@25281.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@25282.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@25283.4]
  assign _T_45 = _T_43 >= 32'h6; // @[Counter.scala 52:70:@25284.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@25286.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@25287.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@25288.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@25289.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@25290.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@25291.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@25294.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@25295.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@25297.4]
  assign RetimeWrapper_clock = clock; // @[:@25300.4]
  assign RetimeWrapper_reset = reset; // @[:@25301.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@25303.4]
  assign RetimeWrapper_io_in = reset ? 32'h5 : _T_62; // @[package.scala 94:16:@25302.4]
endmodule
module NBufController_5( // @[:@25391.2]
  input        clock, // @[:@25392.4]
  input        reset, // @[:@25393.4]
  input        io_sEn_0, // @[:@25394.4]
  input        io_sEn_1, // @[:@25394.4]
  input        io_sEn_2, // @[:@25394.4]
  input        io_sEn_3, // @[:@25394.4]
  input        io_sEn_4, // @[:@25394.4]
  input        io_sEn_5, // @[:@25394.4]
  input        io_sDone_0, // @[:@25394.4]
  input        io_sDone_1, // @[:@25394.4]
  input        io_sDone_2, // @[:@25394.4]
  input        io_sDone_3, // @[:@25394.4]
  input        io_sDone_4, // @[:@25394.4]
  input        io_sDone_5, // @[:@25394.4]
  output [3:0] io_statesInW_0, // @[:@25394.4]
  output [3:0] io_statesInW_1, // @[:@25394.4]
  output [3:0] io_statesInR_1, // @[:@25394.4]
  output [3:0] io_statesInR_5 // @[:@25394.4]
);
  wire  sEn_latch_0_clock; // @[NBuffers.scala 21:52:@25396.4]
  wire  sEn_latch_0_reset; // @[NBuffers.scala 21:52:@25396.4]
  wire  sEn_latch_0_io_input_set; // @[NBuffers.scala 21:52:@25396.4]
  wire  sEn_latch_0_io_input_reset; // @[NBuffers.scala 21:52:@25396.4]
  wire  sEn_latch_0_io_input_asyn_reset; // @[NBuffers.scala 21:52:@25396.4]
  wire  sEn_latch_0_io_output; // @[NBuffers.scala 21:52:@25396.4]
  wire  sEn_latch_1_clock; // @[NBuffers.scala 21:52:@25399.4]
  wire  sEn_latch_1_reset; // @[NBuffers.scala 21:52:@25399.4]
  wire  sEn_latch_1_io_input_set; // @[NBuffers.scala 21:52:@25399.4]
  wire  sEn_latch_1_io_input_reset; // @[NBuffers.scala 21:52:@25399.4]
  wire  sEn_latch_1_io_input_asyn_reset; // @[NBuffers.scala 21:52:@25399.4]
  wire  sEn_latch_1_io_output; // @[NBuffers.scala 21:52:@25399.4]
  wire  sEn_latch_2_clock; // @[NBuffers.scala 21:52:@25402.4]
  wire  sEn_latch_2_reset; // @[NBuffers.scala 21:52:@25402.4]
  wire  sEn_latch_2_io_input_set; // @[NBuffers.scala 21:52:@25402.4]
  wire  sEn_latch_2_io_input_reset; // @[NBuffers.scala 21:52:@25402.4]
  wire  sEn_latch_2_io_input_asyn_reset; // @[NBuffers.scala 21:52:@25402.4]
  wire  sEn_latch_2_io_output; // @[NBuffers.scala 21:52:@25402.4]
  wire  sEn_latch_3_clock; // @[NBuffers.scala 21:52:@25405.4]
  wire  sEn_latch_3_reset; // @[NBuffers.scala 21:52:@25405.4]
  wire  sEn_latch_3_io_input_set; // @[NBuffers.scala 21:52:@25405.4]
  wire  sEn_latch_3_io_input_reset; // @[NBuffers.scala 21:52:@25405.4]
  wire  sEn_latch_3_io_input_asyn_reset; // @[NBuffers.scala 21:52:@25405.4]
  wire  sEn_latch_3_io_output; // @[NBuffers.scala 21:52:@25405.4]
  wire  sEn_latch_4_clock; // @[NBuffers.scala 21:52:@25408.4]
  wire  sEn_latch_4_reset; // @[NBuffers.scala 21:52:@25408.4]
  wire  sEn_latch_4_io_input_set; // @[NBuffers.scala 21:52:@25408.4]
  wire  sEn_latch_4_io_input_reset; // @[NBuffers.scala 21:52:@25408.4]
  wire  sEn_latch_4_io_input_asyn_reset; // @[NBuffers.scala 21:52:@25408.4]
  wire  sEn_latch_4_io_output; // @[NBuffers.scala 21:52:@25408.4]
  wire  sEn_latch_5_clock; // @[NBuffers.scala 21:52:@25411.4]
  wire  sEn_latch_5_reset; // @[NBuffers.scala 21:52:@25411.4]
  wire  sEn_latch_5_io_input_set; // @[NBuffers.scala 21:52:@25411.4]
  wire  sEn_latch_5_io_input_reset; // @[NBuffers.scala 21:52:@25411.4]
  wire  sEn_latch_5_io_input_asyn_reset; // @[NBuffers.scala 21:52:@25411.4]
  wire  sEn_latch_5_io_output; // @[NBuffers.scala 21:52:@25411.4]
  wire  sDone_latch_0_clock; // @[NBuffers.scala 22:54:@25414.4]
  wire  sDone_latch_0_reset; // @[NBuffers.scala 22:54:@25414.4]
  wire  sDone_latch_0_io_input_set; // @[NBuffers.scala 22:54:@25414.4]
  wire  sDone_latch_0_io_input_reset; // @[NBuffers.scala 22:54:@25414.4]
  wire  sDone_latch_0_io_input_asyn_reset; // @[NBuffers.scala 22:54:@25414.4]
  wire  sDone_latch_0_io_output; // @[NBuffers.scala 22:54:@25414.4]
  wire  sDone_latch_1_clock; // @[NBuffers.scala 22:54:@25417.4]
  wire  sDone_latch_1_reset; // @[NBuffers.scala 22:54:@25417.4]
  wire  sDone_latch_1_io_input_set; // @[NBuffers.scala 22:54:@25417.4]
  wire  sDone_latch_1_io_input_reset; // @[NBuffers.scala 22:54:@25417.4]
  wire  sDone_latch_1_io_input_asyn_reset; // @[NBuffers.scala 22:54:@25417.4]
  wire  sDone_latch_1_io_output; // @[NBuffers.scala 22:54:@25417.4]
  wire  sDone_latch_2_clock; // @[NBuffers.scala 22:54:@25420.4]
  wire  sDone_latch_2_reset; // @[NBuffers.scala 22:54:@25420.4]
  wire  sDone_latch_2_io_input_set; // @[NBuffers.scala 22:54:@25420.4]
  wire  sDone_latch_2_io_input_reset; // @[NBuffers.scala 22:54:@25420.4]
  wire  sDone_latch_2_io_input_asyn_reset; // @[NBuffers.scala 22:54:@25420.4]
  wire  sDone_latch_2_io_output; // @[NBuffers.scala 22:54:@25420.4]
  wire  sDone_latch_3_clock; // @[NBuffers.scala 22:54:@25423.4]
  wire  sDone_latch_3_reset; // @[NBuffers.scala 22:54:@25423.4]
  wire  sDone_latch_3_io_input_set; // @[NBuffers.scala 22:54:@25423.4]
  wire  sDone_latch_3_io_input_reset; // @[NBuffers.scala 22:54:@25423.4]
  wire  sDone_latch_3_io_input_asyn_reset; // @[NBuffers.scala 22:54:@25423.4]
  wire  sDone_latch_3_io_output; // @[NBuffers.scala 22:54:@25423.4]
  wire  sDone_latch_4_clock; // @[NBuffers.scala 22:54:@25426.4]
  wire  sDone_latch_4_reset; // @[NBuffers.scala 22:54:@25426.4]
  wire  sDone_latch_4_io_input_set; // @[NBuffers.scala 22:54:@25426.4]
  wire  sDone_latch_4_io_input_reset; // @[NBuffers.scala 22:54:@25426.4]
  wire  sDone_latch_4_io_input_asyn_reset; // @[NBuffers.scala 22:54:@25426.4]
  wire  sDone_latch_4_io_output; // @[NBuffers.scala 22:54:@25426.4]
  wire  sDone_latch_5_clock; // @[NBuffers.scala 22:54:@25429.4]
  wire  sDone_latch_5_reset; // @[NBuffers.scala 22:54:@25429.4]
  wire  sDone_latch_5_io_input_set; // @[NBuffers.scala 22:54:@25429.4]
  wire  sDone_latch_5_io_input_reset; // @[NBuffers.scala 22:54:@25429.4]
  wire  sDone_latch_5_io_input_asyn_reset; // @[NBuffers.scala 22:54:@25429.4]
  wire  sDone_latch_5_io_output; // @[NBuffers.scala 22:54:@25429.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@25436.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@25436.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@25436.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@25436.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@25436.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@25444.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@25444.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@25444.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@25444.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@25444.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@25453.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@25453.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@25453.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@25453.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@25453.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@25461.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@25461.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@25461.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@25461.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@25461.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@25472.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@25472.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@25472.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@25472.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@25472.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@25480.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@25480.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@25480.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@25480.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@25480.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@25489.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@25489.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@25489.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@25489.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@25489.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@25497.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@25497.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@25497.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@25497.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@25497.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@25508.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@25508.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@25508.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@25508.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@25508.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@25516.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@25516.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@25516.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@25516.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@25516.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@25525.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@25525.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@25525.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@25525.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@25525.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@25533.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@25533.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@25533.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@25533.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@25533.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@25544.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@25544.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@25544.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@25544.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@25544.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@25552.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@25552.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@25552.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@25552.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@25552.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@25561.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@25561.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@25561.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@25561.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@25561.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@25569.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@25569.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@25569.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@25569.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@25569.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@25580.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@25580.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@25580.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@25580.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@25580.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@25588.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@25588.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@25588.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@25588.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@25588.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@25597.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@25597.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@25597.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@25597.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@25597.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@25605.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@25605.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@25605.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@25605.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@25605.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@25616.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@25616.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@25616.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@25616.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@25616.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@25624.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@25624.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@25624.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@25624.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@25624.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@25633.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@25633.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@25633.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@25633.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@25633.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@25641.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@25641.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@25641.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@25641.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@25641.4]
  wire  NBufCtr_clock; // @[NBuffers.scala 40:19:@25678.4]
  wire  NBufCtr_reset; // @[NBuffers.scala 40:19:@25678.4]
  wire  NBufCtr_io_input_countUp; // @[NBuffers.scala 40:19:@25678.4]
  wire  NBufCtr_io_input_enable; // @[NBuffers.scala 40:19:@25678.4]
  wire [31:0] NBufCtr_io_output_count; // @[NBuffers.scala 40:19:@25678.4]
  wire  NBufCtr_1_clock; // @[NBuffers.scala 40:19:@25689.4]
  wire  NBufCtr_1_reset; // @[NBuffers.scala 40:19:@25689.4]
  wire  NBufCtr_1_io_input_countUp; // @[NBuffers.scala 40:19:@25689.4]
  wire  NBufCtr_1_io_input_enable; // @[NBuffers.scala 40:19:@25689.4]
  wire [31:0] NBufCtr_1_io_output_count; // @[NBuffers.scala 40:19:@25689.4]
  wire  statesInR_0_clock; // @[NBuffers.scala 50:19:@25700.4]
  wire  statesInR_0_reset; // @[NBuffers.scala 50:19:@25700.4]
  wire  statesInR_0_io_input_countUp; // @[NBuffers.scala 50:19:@25700.4]
  wire  statesInR_0_io_input_enable; // @[NBuffers.scala 50:19:@25700.4]
  wire [31:0] statesInR_0_io_output_count; // @[NBuffers.scala 50:19:@25700.4]
  wire  statesInR_1_clock; // @[NBuffers.scala 50:19:@25711.4]
  wire  statesInR_1_reset; // @[NBuffers.scala 50:19:@25711.4]
  wire  statesInR_1_io_input_countUp; // @[NBuffers.scala 50:19:@25711.4]
  wire  statesInR_1_io_input_enable; // @[NBuffers.scala 50:19:@25711.4]
  wire [31:0] statesInR_1_io_output_count; // @[NBuffers.scala 50:19:@25711.4]
  wire  statesInR_2_clock; // @[NBuffers.scala 50:19:@25722.4]
  wire  statesInR_2_reset; // @[NBuffers.scala 50:19:@25722.4]
  wire  statesInR_2_io_input_countUp; // @[NBuffers.scala 50:19:@25722.4]
  wire  statesInR_2_io_input_enable; // @[NBuffers.scala 50:19:@25722.4]
  wire  statesInR_3_clock; // @[NBuffers.scala 50:19:@25733.4]
  wire  statesInR_3_reset; // @[NBuffers.scala 50:19:@25733.4]
  wire  statesInR_3_io_input_countUp; // @[NBuffers.scala 50:19:@25733.4]
  wire  statesInR_3_io_input_enable; // @[NBuffers.scala 50:19:@25733.4]
  wire  statesInR_4_clock; // @[NBuffers.scala 50:19:@25744.4]
  wire  statesInR_4_reset; // @[NBuffers.scala 50:19:@25744.4]
  wire  statesInR_4_io_input_countUp; // @[NBuffers.scala 50:19:@25744.4]
  wire  statesInR_4_io_input_enable; // @[NBuffers.scala 50:19:@25744.4]
  wire  statesInR_5_clock; // @[NBuffers.scala 50:19:@25755.4]
  wire  statesInR_5_reset; // @[NBuffers.scala 50:19:@25755.4]
  wire  statesInR_5_io_input_countUp; // @[NBuffers.scala 50:19:@25755.4]
  wire  statesInR_5_io_input_enable; // @[NBuffers.scala 50:19:@25755.4]
  wire [31:0] statesInR_5_io_output_count; // @[NBuffers.scala 50:19:@25755.4]
  wire  _T_33; // @[NBuffers.scala 26:46:@25433.4]
  wire  _T_48; // @[NBuffers.scala 26:46:@25469.4]
  wire  _T_63; // @[NBuffers.scala 26:46:@25505.4]
  wire  _T_78; // @[NBuffers.scala 26:46:@25541.4]
  wire  _T_93; // @[NBuffers.scala 26:46:@25577.4]
  wire  _T_108; // @[NBuffers.scala 26:46:@25613.4]
  wire  _T_122; // @[NBuffers.scala 33:64:@25649.4]
  wire  _T_123; // @[NBuffers.scala 33:64:@25650.4]
  wire  _T_124; // @[NBuffers.scala 33:64:@25651.4]
  wire  _T_125; // @[NBuffers.scala 33:64:@25652.4]
  wire  anyEnabled; // @[NBuffers.scala 33:64:@25653.4]
  wire  _T_126; // @[NBuffers.scala 34:124:@25654.4]
  wire  _T_127; // @[NBuffers.scala 34:104:@25655.4]
  wire  _T_128; // @[NBuffers.scala 34:124:@25656.4]
  wire  _T_129; // @[NBuffers.scala 34:104:@25657.4]
  wire  _T_130; // @[NBuffers.scala 34:124:@25658.4]
  wire  _T_131; // @[NBuffers.scala 34:104:@25659.4]
  wire  _T_132; // @[NBuffers.scala 34:124:@25660.4]
  wire  _T_133; // @[NBuffers.scala 34:104:@25661.4]
  wire  _T_134; // @[NBuffers.scala 34:124:@25662.4]
  wire  _T_135; // @[NBuffers.scala 34:104:@25663.4]
  wire  _T_136; // @[NBuffers.scala 34:124:@25664.4]
  wire  _T_137; // @[NBuffers.scala 34:104:@25665.4]
  wire  _T_138; // @[NBuffers.scala 34:150:@25666.4]
  wire  _T_139; // @[NBuffers.scala 34:150:@25667.4]
  wire  _T_140; // @[NBuffers.scala 34:150:@25668.4]
  wire  _T_141; // @[NBuffers.scala 34:150:@25669.4]
  wire  _T_142; // @[NBuffers.scala 34:150:@25670.4]
  wire  _T_143; // @[NBuffers.scala 34:154:@25671.4]
  wire  _T_145; // @[package.scala 100:49:@25672.4]
  reg  _T_148; // @[package.scala 48:56:@25673.4]
  reg [31:0] _RAND_0;
  SRFF sEn_latch_0 ( // @[NBuffers.scala 21:52:@25396.4]
    .clock(sEn_latch_0_clock),
    .reset(sEn_latch_0_reset),
    .io_input_set(sEn_latch_0_io_input_set),
    .io_input_reset(sEn_latch_0_io_input_reset),
    .io_input_asyn_reset(sEn_latch_0_io_input_asyn_reset),
    .io_output(sEn_latch_0_io_output)
  );
  SRFF sEn_latch_1 ( // @[NBuffers.scala 21:52:@25399.4]
    .clock(sEn_latch_1_clock),
    .reset(sEn_latch_1_reset),
    .io_input_set(sEn_latch_1_io_input_set),
    .io_input_reset(sEn_latch_1_io_input_reset),
    .io_input_asyn_reset(sEn_latch_1_io_input_asyn_reset),
    .io_output(sEn_latch_1_io_output)
  );
  SRFF sEn_latch_2 ( // @[NBuffers.scala 21:52:@25402.4]
    .clock(sEn_latch_2_clock),
    .reset(sEn_latch_2_reset),
    .io_input_set(sEn_latch_2_io_input_set),
    .io_input_reset(sEn_latch_2_io_input_reset),
    .io_input_asyn_reset(sEn_latch_2_io_input_asyn_reset),
    .io_output(sEn_latch_2_io_output)
  );
  SRFF sEn_latch_3 ( // @[NBuffers.scala 21:52:@25405.4]
    .clock(sEn_latch_3_clock),
    .reset(sEn_latch_3_reset),
    .io_input_set(sEn_latch_3_io_input_set),
    .io_input_reset(sEn_latch_3_io_input_reset),
    .io_input_asyn_reset(sEn_latch_3_io_input_asyn_reset),
    .io_output(sEn_latch_3_io_output)
  );
  SRFF sEn_latch_4 ( // @[NBuffers.scala 21:52:@25408.4]
    .clock(sEn_latch_4_clock),
    .reset(sEn_latch_4_reset),
    .io_input_set(sEn_latch_4_io_input_set),
    .io_input_reset(sEn_latch_4_io_input_reset),
    .io_input_asyn_reset(sEn_latch_4_io_input_asyn_reset),
    .io_output(sEn_latch_4_io_output)
  );
  SRFF sEn_latch_5 ( // @[NBuffers.scala 21:52:@25411.4]
    .clock(sEn_latch_5_clock),
    .reset(sEn_latch_5_reset),
    .io_input_set(sEn_latch_5_io_input_set),
    .io_input_reset(sEn_latch_5_io_input_reset),
    .io_input_asyn_reset(sEn_latch_5_io_input_asyn_reset),
    .io_output(sEn_latch_5_io_output)
  );
  SRFF sDone_latch_0 ( // @[NBuffers.scala 22:54:@25414.4]
    .clock(sDone_latch_0_clock),
    .reset(sDone_latch_0_reset),
    .io_input_set(sDone_latch_0_io_input_set),
    .io_input_reset(sDone_latch_0_io_input_reset),
    .io_input_asyn_reset(sDone_latch_0_io_input_asyn_reset),
    .io_output(sDone_latch_0_io_output)
  );
  SRFF sDone_latch_1 ( // @[NBuffers.scala 22:54:@25417.4]
    .clock(sDone_latch_1_clock),
    .reset(sDone_latch_1_reset),
    .io_input_set(sDone_latch_1_io_input_set),
    .io_input_reset(sDone_latch_1_io_input_reset),
    .io_input_asyn_reset(sDone_latch_1_io_input_asyn_reset),
    .io_output(sDone_latch_1_io_output)
  );
  SRFF sDone_latch_2 ( // @[NBuffers.scala 22:54:@25420.4]
    .clock(sDone_latch_2_clock),
    .reset(sDone_latch_2_reset),
    .io_input_set(sDone_latch_2_io_input_set),
    .io_input_reset(sDone_latch_2_io_input_reset),
    .io_input_asyn_reset(sDone_latch_2_io_input_asyn_reset),
    .io_output(sDone_latch_2_io_output)
  );
  SRFF sDone_latch_3 ( // @[NBuffers.scala 22:54:@25423.4]
    .clock(sDone_latch_3_clock),
    .reset(sDone_latch_3_reset),
    .io_input_set(sDone_latch_3_io_input_set),
    .io_input_reset(sDone_latch_3_io_input_reset),
    .io_input_asyn_reset(sDone_latch_3_io_input_asyn_reset),
    .io_output(sDone_latch_3_io_output)
  );
  SRFF sDone_latch_4 ( // @[NBuffers.scala 22:54:@25426.4]
    .clock(sDone_latch_4_clock),
    .reset(sDone_latch_4_reset),
    .io_input_set(sDone_latch_4_io_input_set),
    .io_input_reset(sDone_latch_4_io_input_reset),
    .io_input_asyn_reset(sDone_latch_4_io_input_asyn_reset),
    .io_output(sDone_latch_4_io_output)
  );
  SRFF sDone_latch_5 ( // @[NBuffers.scala 22:54:@25429.4]
    .clock(sDone_latch_5_clock),
    .reset(sDone_latch_5_reset),
    .io_input_set(sDone_latch_5_io_input_set),
    .io_input_reset(sDone_latch_5_io_input_reset),
    .io_input_asyn_reset(sDone_latch_5_io_input_asyn_reset),
    .io_output(sDone_latch_5_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@25436.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@25444.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@25453.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@25461.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@25472.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@25480.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@25489.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@25497.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@25508.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@25516.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@25525.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 ( // @[package.scala 93:22:@25533.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper RetimeWrapper_12 ( // @[package.scala 93:22:@25544.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 ( // @[package.scala 93:22:@25552.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@25561.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@25569.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 ( // @[package.scala 93:22:@25580.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper RetimeWrapper_17 ( // @[package.scala 93:22:@25588.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 ( // @[package.scala 93:22:@25597.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper RetimeWrapper_19 ( // @[package.scala 93:22:@25605.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper RetimeWrapper_20 ( // @[package.scala 93:22:@25616.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper RetimeWrapper_21 ( // @[package.scala 93:22:@25624.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper RetimeWrapper_22 ( // @[package.scala 93:22:@25633.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper RetimeWrapper_23 ( // @[package.scala 93:22:@25641.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  NBufCtr_25 NBufCtr ( // @[NBuffers.scala 40:19:@25678.4]
    .clock(NBufCtr_clock),
    .reset(NBufCtr_reset),
    .io_input_countUp(NBufCtr_io_input_countUp),
    .io_input_enable(NBufCtr_io_input_enable),
    .io_output_count(NBufCtr_io_output_count)
  );
  NBufCtr_26 NBufCtr_1 ( // @[NBuffers.scala 40:19:@25689.4]
    .clock(NBufCtr_1_clock),
    .reset(NBufCtr_1_reset),
    .io_input_countUp(NBufCtr_1_io_input_countUp),
    .io_input_enable(NBufCtr_1_io_input_enable),
    .io_output_count(NBufCtr_1_io_output_count)
  );
  NBufCtr_25 statesInR_0 ( // @[NBuffers.scala 50:19:@25700.4]
    .clock(statesInR_0_clock),
    .reset(statesInR_0_reset),
    .io_input_countUp(statesInR_0_io_input_countUp),
    .io_input_enable(statesInR_0_io_input_enable),
    .io_output_count(statesInR_0_io_output_count)
  );
  NBufCtr_28 statesInR_1 ( // @[NBuffers.scala 50:19:@25711.4]
    .clock(statesInR_1_clock),
    .reset(statesInR_1_reset),
    .io_input_countUp(statesInR_1_io_input_countUp),
    .io_input_enable(statesInR_1_io_input_enable),
    .io_output_count(statesInR_1_io_output_count)
  );
  NBufCtr_29 statesInR_2 ( // @[NBuffers.scala 50:19:@25722.4]
    .clock(statesInR_2_clock),
    .reset(statesInR_2_reset),
    .io_input_countUp(statesInR_2_io_input_countUp),
    .io_input_enable(statesInR_2_io_input_enable)
  );
  NBufCtr_30 statesInR_3 ( // @[NBuffers.scala 50:19:@25733.4]
    .clock(statesInR_3_clock),
    .reset(statesInR_3_reset),
    .io_input_countUp(statesInR_3_io_input_countUp),
    .io_input_enable(statesInR_3_io_input_enable)
  );
  NBufCtr_31 statesInR_4 ( // @[NBuffers.scala 50:19:@25744.4]
    .clock(statesInR_4_clock),
    .reset(statesInR_4_reset),
    .io_input_countUp(statesInR_4_io_input_countUp),
    .io_input_enable(statesInR_4_io_input_enable)
  );
  NBufCtr_26 statesInR_5 ( // @[NBuffers.scala 50:19:@25755.4]
    .clock(statesInR_5_clock),
    .reset(statesInR_5_reset),
    .io_input_countUp(statesInR_5_io_input_countUp),
    .io_input_enable(statesInR_5_io_input_enable),
    .io_output_count(statesInR_5_io_output_count)
  );
  assign _T_33 = io_sDone_0 == 1'h0; // @[NBuffers.scala 26:46:@25433.4]
  assign _T_48 = io_sDone_1 == 1'h0; // @[NBuffers.scala 26:46:@25469.4]
  assign _T_63 = io_sDone_2 == 1'h0; // @[NBuffers.scala 26:46:@25505.4]
  assign _T_78 = io_sDone_3 == 1'h0; // @[NBuffers.scala 26:46:@25541.4]
  assign _T_93 = io_sDone_4 == 1'h0; // @[NBuffers.scala 26:46:@25577.4]
  assign _T_108 = io_sDone_5 == 1'h0; // @[NBuffers.scala 26:46:@25613.4]
  assign _T_122 = sEn_latch_0_io_output | sEn_latch_1_io_output; // @[NBuffers.scala 33:64:@25649.4]
  assign _T_123 = _T_122 | sEn_latch_2_io_output; // @[NBuffers.scala 33:64:@25650.4]
  assign _T_124 = _T_123 | sEn_latch_3_io_output; // @[NBuffers.scala 33:64:@25651.4]
  assign _T_125 = _T_124 | sEn_latch_4_io_output; // @[NBuffers.scala 33:64:@25652.4]
  assign anyEnabled = _T_125 | sEn_latch_5_io_output; // @[NBuffers.scala 33:64:@25653.4]
  assign _T_126 = sDone_latch_0_io_output | io_sDone_0; // @[NBuffers.scala 34:124:@25654.4]
  assign _T_127 = sEn_latch_0_io_output == _T_126; // @[NBuffers.scala 34:104:@25655.4]
  assign _T_128 = sDone_latch_1_io_output | io_sDone_1; // @[NBuffers.scala 34:124:@25656.4]
  assign _T_129 = sEn_latch_1_io_output == _T_128; // @[NBuffers.scala 34:104:@25657.4]
  assign _T_130 = sDone_latch_2_io_output | io_sDone_2; // @[NBuffers.scala 34:124:@25658.4]
  assign _T_131 = sEn_latch_2_io_output == _T_130; // @[NBuffers.scala 34:104:@25659.4]
  assign _T_132 = sDone_latch_3_io_output | io_sDone_3; // @[NBuffers.scala 34:124:@25660.4]
  assign _T_133 = sEn_latch_3_io_output == _T_132; // @[NBuffers.scala 34:104:@25661.4]
  assign _T_134 = sDone_latch_4_io_output | io_sDone_4; // @[NBuffers.scala 34:124:@25662.4]
  assign _T_135 = sEn_latch_4_io_output == _T_134; // @[NBuffers.scala 34:104:@25663.4]
  assign _T_136 = sDone_latch_5_io_output | io_sDone_5; // @[NBuffers.scala 34:124:@25664.4]
  assign _T_137 = sEn_latch_5_io_output == _T_136; // @[NBuffers.scala 34:104:@25665.4]
  assign _T_138 = _T_127 & _T_129; // @[NBuffers.scala 34:150:@25666.4]
  assign _T_139 = _T_138 & _T_131; // @[NBuffers.scala 34:150:@25667.4]
  assign _T_140 = _T_139 & _T_133; // @[NBuffers.scala 34:150:@25668.4]
  assign _T_141 = _T_140 & _T_135; // @[NBuffers.scala 34:150:@25669.4]
  assign _T_142 = _T_141 & _T_137; // @[NBuffers.scala 34:150:@25670.4]
  assign _T_143 = _T_142 & anyEnabled; // @[NBuffers.scala 34:154:@25671.4]
  assign _T_145 = _T_143 == 1'h0; // @[package.scala 100:49:@25672.4]
  assign io_statesInW_0 = NBufCtr_io_output_count[3:0]; // @[NBuffers.scala 44:21:@25688.4]
  assign io_statesInW_1 = NBufCtr_1_io_output_count[3:0]; // @[NBuffers.scala 44:21:@25699.4]
  assign io_statesInR_1 = statesInR_1_io_output_count[3:0]; // @[NBuffers.scala 54:21:@25721.4]
  assign io_statesInR_5 = statesInR_5_io_output_count[3:0]; // @[NBuffers.scala 54:21:@25765.4]
  assign sEn_latch_0_clock = clock; // @[:@25397.4]
  assign sEn_latch_0_reset = reset; // @[:@25398.4]
  assign sEn_latch_0_io_input_set = io_sEn_0 & _T_33; // @[NBuffers.scala 26:31:@25435.4]
  assign sEn_latch_0_io_input_reset = RetimeWrapper_io_out; // @[NBuffers.scala 27:33:@25443.4]
  assign sEn_latch_0_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[NBuffers.scala 28:38:@25451.4]
  assign sEn_latch_1_clock = clock; // @[:@25400.4]
  assign sEn_latch_1_reset = reset; // @[:@25401.4]
  assign sEn_latch_1_io_input_set = io_sEn_1 & _T_48; // @[NBuffers.scala 26:31:@25471.4]
  assign sEn_latch_1_io_input_reset = RetimeWrapper_4_io_out; // @[NBuffers.scala 27:33:@25479.4]
  assign sEn_latch_1_io_input_asyn_reset = RetimeWrapper_5_io_out; // @[NBuffers.scala 28:38:@25487.4]
  assign sEn_latch_2_clock = clock; // @[:@25403.4]
  assign sEn_latch_2_reset = reset; // @[:@25404.4]
  assign sEn_latch_2_io_input_set = io_sEn_2 & _T_63; // @[NBuffers.scala 26:31:@25507.4]
  assign sEn_latch_2_io_input_reset = RetimeWrapper_8_io_out; // @[NBuffers.scala 27:33:@25515.4]
  assign sEn_latch_2_io_input_asyn_reset = RetimeWrapper_9_io_out; // @[NBuffers.scala 28:38:@25523.4]
  assign sEn_latch_3_clock = clock; // @[:@25406.4]
  assign sEn_latch_3_reset = reset; // @[:@25407.4]
  assign sEn_latch_3_io_input_set = io_sEn_3 & _T_78; // @[NBuffers.scala 26:31:@25543.4]
  assign sEn_latch_3_io_input_reset = RetimeWrapper_12_io_out; // @[NBuffers.scala 27:33:@25551.4]
  assign sEn_latch_3_io_input_asyn_reset = RetimeWrapper_13_io_out; // @[NBuffers.scala 28:38:@25559.4]
  assign sEn_latch_4_clock = clock; // @[:@25409.4]
  assign sEn_latch_4_reset = reset; // @[:@25410.4]
  assign sEn_latch_4_io_input_set = io_sEn_4 & _T_93; // @[NBuffers.scala 26:31:@25579.4]
  assign sEn_latch_4_io_input_reset = RetimeWrapper_16_io_out; // @[NBuffers.scala 27:33:@25587.4]
  assign sEn_latch_4_io_input_asyn_reset = RetimeWrapper_17_io_out; // @[NBuffers.scala 28:38:@25595.4]
  assign sEn_latch_5_clock = clock; // @[:@25412.4]
  assign sEn_latch_5_reset = reset; // @[:@25413.4]
  assign sEn_latch_5_io_input_set = io_sEn_5 & _T_108; // @[NBuffers.scala 26:31:@25615.4]
  assign sEn_latch_5_io_input_reset = RetimeWrapper_20_io_out; // @[NBuffers.scala 27:33:@25623.4]
  assign sEn_latch_5_io_input_asyn_reset = RetimeWrapper_21_io_out; // @[NBuffers.scala 28:38:@25631.4]
  assign sDone_latch_0_clock = clock; // @[:@25415.4]
  assign sDone_latch_0_reset = reset; // @[:@25416.4]
  assign sDone_latch_0_io_input_set = io_sDone_0; // @[NBuffers.scala 29:33:@25452.4]
  assign sDone_latch_0_io_input_reset = RetimeWrapper_2_io_out; // @[NBuffers.scala 30:35:@25460.4]
  assign sDone_latch_0_io_input_asyn_reset = RetimeWrapper_3_io_out; // @[NBuffers.scala 31:40:@25468.4]
  assign sDone_latch_1_clock = clock; // @[:@25418.4]
  assign sDone_latch_1_reset = reset; // @[:@25419.4]
  assign sDone_latch_1_io_input_set = io_sDone_1; // @[NBuffers.scala 29:33:@25488.4]
  assign sDone_latch_1_io_input_reset = RetimeWrapper_6_io_out; // @[NBuffers.scala 30:35:@25496.4]
  assign sDone_latch_1_io_input_asyn_reset = RetimeWrapper_7_io_out; // @[NBuffers.scala 31:40:@25504.4]
  assign sDone_latch_2_clock = clock; // @[:@25421.4]
  assign sDone_latch_2_reset = reset; // @[:@25422.4]
  assign sDone_latch_2_io_input_set = io_sDone_2; // @[NBuffers.scala 29:33:@25524.4]
  assign sDone_latch_2_io_input_reset = RetimeWrapper_10_io_out; // @[NBuffers.scala 30:35:@25532.4]
  assign sDone_latch_2_io_input_asyn_reset = RetimeWrapper_11_io_out; // @[NBuffers.scala 31:40:@25540.4]
  assign sDone_latch_3_clock = clock; // @[:@25424.4]
  assign sDone_latch_3_reset = reset; // @[:@25425.4]
  assign sDone_latch_3_io_input_set = io_sDone_3; // @[NBuffers.scala 29:33:@25560.4]
  assign sDone_latch_3_io_input_reset = RetimeWrapper_14_io_out; // @[NBuffers.scala 30:35:@25568.4]
  assign sDone_latch_3_io_input_asyn_reset = RetimeWrapper_15_io_out; // @[NBuffers.scala 31:40:@25576.4]
  assign sDone_latch_4_clock = clock; // @[:@25427.4]
  assign sDone_latch_4_reset = reset; // @[:@25428.4]
  assign sDone_latch_4_io_input_set = io_sDone_4; // @[NBuffers.scala 29:33:@25596.4]
  assign sDone_latch_4_io_input_reset = RetimeWrapper_18_io_out; // @[NBuffers.scala 30:35:@25604.4]
  assign sDone_latch_4_io_input_asyn_reset = RetimeWrapper_19_io_out; // @[NBuffers.scala 31:40:@25612.4]
  assign sDone_latch_5_clock = clock; // @[:@25430.4]
  assign sDone_latch_5_reset = reset; // @[:@25431.4]
  assign sDone_latch_5_io_input_set = io_sDone_5; // @[NBuffers.scala 29:33:@25632.4]
  assign sDone_latch_5_io_input_reset = RetimeWrapper_22_io_out; // @[NBuffers.scala 30:35:@25640.4]
  assign sDone_latch_5_io_input_asyn_reset = RetimeWrapper_23_io_out; // @[NBuffers.scala 31:40:@25648.4]
  assign RetimeWrapper_clock = clock; // @[:@25437.4]
  assign RetimeWrapper_reset = reset; // @[:@25438.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@25440.4]
  assign RetimeWrapper_io_in = _T_143 & _T_148; // @[package.scala 94:16:@25439.4]
  assign RetimeWrapper_1_clock = clock; // @[:@25445.4]
  assign RetimeWrapper_1_reset = reset; // @[:@25446.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@25448.4]
  assign RetimeWrapper_1_io_in = reset; // @[package.scala 94:16:@25447.4]
  assign RetimeWrapper_2_clock = clock; // @[:@25454.4]
  assign RetimeWrapper_2_reset = reset; // @[:@25455.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@25457.4]
  assign RetimeWrapper_2_io_in = _T_143 & _T_148; // @[package.scala 94:16:@25456.4]
  assign RetimeWrapper_3_clock = clock; // @[:@25462.4]
  assign RetimeWrapper_3_reset = reset; // @[:@25463.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@25465.4]
  assign RetimeWrapper_3_io_in = reset; // @[package.scala 94:16:@25464.4]
  assign RetimeWrapper_4_clock = clock; // @[:@25473.4]
  assign RetimeWrapper_4_reset = reset; // @[:@25474.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@25476.4]
  assign RetimeWrapper_4_io_in = _T_143 & _T_148; // @[package.scala 94:16:@25475.4]
  assign RetimeWrapper_5_clock = clock; // @[:@25481.4]
  assign RetimeWrapper_5_reset = reset; // @[:@25482.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@25484.4]
  assign RetimeWrapper_5_io_in = reset; // @[package.scala 94:16:@25483.4]
  assign RetimeWrapper_6_clock = clock; // @[:@25490.4]
  assign RetimeWrapper_6_reset = reset; // @[:@25491.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@25493.4]
  assign RetimeWrapper_6_io_in = _T_143 & _T_148; // @[package.scala 94:16:@25492.4]
  assign RetimeWrapper_7_clock = clock; // @[:@25498.4]
  assign RetimeWrapper_7_reset = reset; // @[:@25499.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@25501.4]
  assign RetimeWrapper_7_io_in = reset; // @[package.scala 94:16:@25500.4]
  assign RetimeWrapper_8_clock = clock; // @[:@25509.4]
  assign RetimeWrapper_8_reset = reset; // @[:@25510.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@25512.4]
  assign RetimeWrapper_8_io_in = _T_143 & _T_148; // @[package.scala 94:16:@25511.4]
  assign RetimeWrapper_9_clock = clock; // @[:@25517.4]
  assign RetimeWrapper_9_reset = reset; // @[:@25518.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@25520.4]
  assign RetimeWrapper_9_io_in = reset; // @[package.scala 94:16:@25519.4]
  assign RetimeWrapper_10_clock = clock; // @[:@25526.4]
  assign RetimeWrapper_10_reset = reset; // @[:@25527.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@25529.4]
  assign RetimeWrapper_10_io_in = _T_143 & _T_148; // @[package.scala 94:16:@25528.4]
  assign RetimeWrapper_11_clock = clock; // @[:@25534.4]
  assign RetimeWrapper_11_reset = reset; // @[:@25535.4]
  assign RetimeWrapper_11_io_flow = 1'h1; // @[package.scala 95:18:@25537.4]
  assign RetimeWrapper_11_io_in = reset; // @[package.scala 94:16:@25536.4]
  assign RetimeWrapper_12_clock = clock; // @[:@25545.4]
  assign RetimeWrapper_12_reset = reset; // @[:@25546.4]
  assign RetimeWrapper_12_io_flow = 1'h1; // @[package.scala 95:18:@25548.4]
  assign RetimeWrapper_12_io_in = _T_143 & _T_148; // @[package.scala 94:16:@25547.4]
  assign RetimeWrapper_13_clock = clock; // @[:@25553.4]
  assign RetimeWrapper_13_reset = reset; // @[:@25554.4]
  assign RetimeWrapper_13_io_flow = 1'h1; // @[package.scala 95:18:@25556.4]
  assign RetimeWrapper_13_io_in = reset; // @[package.scala 94:16:@25555.4]
  assign RetimeWrapper_14_clock = clock; // @[:@25562.4]
  assign RetimeWrapper_14_reset = reset; // @[:@25563.4]
  assign RetimeWrapper_14_io_flow = 1'h1; // @[package.scala 95:18:@25565.4]
  assign RetimeWrapper_14_io_in = _T_143 & _T_148; // @[package.scala 94:16:@25564.4]
  assign RetimeWrapper_15_clock = clock; // @[:@25570.4]
  assign RetimeWrapper_15_reset = reset; // @[:@25571.4]
  assign RetimeWrapper_15_io_flow = 1'h1; // @[package.scala 95:18:@25573.4]
  assign RetimeWrapper_15_io_in = reset; // @[package.scala 94:16:@25572.4]
  assign RetimeWrapper_16_clock = clock; // @[:@25581.4]
  assign RetimeWrapper_16_reset = reset; // @[:@25582.4]
  assign RetimeWrapper_16_io_flow = 1'h1; // @[package.scala 95:18:@25584.4]
  assign RetimeWrapper_16_io_in = _T_143 & _T_148; // @[package.scala 94:16:@25583.4]
  assign RetimeWrapper_17_clock = clock; // @[:@25589.4]
  assign RetimeWrapper_17_reset = reset; // @[:@25590.4]
  assign RetimeWrapper_17_io_flow = 1'h1; // @[package.scala 95:18:@25592.4]
  assign RetimeWrapper_17_io_in = reset; // @[package.scala 94:16:@25591.4]
  assign RetimeWrapper_18_clock = clock; // @[:@25598.4]
  assign RetimeWrapper_18_reset = reset; // @[:@25599.4]
  assign RetimeWrapper_18_io_flow = 1'h1; // @[package.scala 95:18:@25601.4]
  assign RetimeWrapper_18_io_in = _T_143 & _T_148; // @[package.scala 94:16:@25600.4]
  assign RetimeWrapper_19_clock = clock; // @[:@25606.4]
  assign RetimeWrapper_19_reset = reset; // @[:@25607.4]
  assign RetimeWrapper_19_io_flow = 1'h1; // @[package.scala 95:18:@25609.4]
  assign RetimeWrapper_19_io_in = reset; // @[package.scala 94:16:@25608.4]
  assign RetimeWrapper_20_clock = clock; // @[:@25617.4]
  assign RetimeWrapper_20_reset = reset; // @[:@25618.4]
  assign RetimeWrapper_20_io_flow = 1'h1; // @[package.scala 95:18:@25620.4]
  assign RetimeWrapper_20_io_in = _T_143 & _T_148; // @[package.scala 94:16:@25619.4]
  assign RetimeWrapper_21_clock = clock; // @[:@25625.4]
  assign RetimeWrapper_21_reset = reset; // @[:@25626.4]
  assign RetimeWrapper_21_io_flow = 1'h1; // @[package.scala 95:18:@25628.4]
  assign RetimeWrapper_21_io_in = reset; // @[package.scala 94:16:@25627.4]
  assign RetimeWrapper_22_clock = clock; // @[:@25634.4]
  assign RetimeWrapper_22_reset = reset; // @[:@25635.4]
  assign RetimeWrapper_22_io_flow = 1'h1; // @[package.scala 95:18:@25637.4]
  assign RetimeWrapper_22_io_in = _T_143 & _T_148; // @[package.scala 94:16:@25636.4]
  assign RetimeWrapper_23_clock = clock; // @[:@25642.4]
  assign RetimeWrapper_23_reset = reset; // @[:@25643.4]
  assign RetimeWrapper_23_io_flow = 1'h1; // @[package.scala 95:18:@25645.4]
  assign RetimeWrapper_23_io_in = reset; // @[package.scala 94:16:@25644.4]
  assign NBufCtr_clock = clock; // @[:@25679.4]
  assign NBufCtr_reset = reset; // @[:@25680.4]
  assign NBufCtr_io_input_countUp = 1'h0; // @[NBuffers.scala 43:24:@25687.4]
  assign NBufCtr_io_input_enable = _T_143 & _T_148; // @[NBuffers.scala 42:23:@25686.4]
  assign NBufCtr_1_clock = clock; // @[:@25690.4]
  assign NBufCtr_1_reset = reset; // @[:@25691.4]
  assign NBufCtr_1_io_input_countUp = 1'h0; // @[NBuffers.scala 43:24:@25698.4]
  assign NBufCtr_1_io_input_enable = _T_143 & _T_148; // @[NBuffers.scala 42:23:@25697.4]
  assign statesInR_0_clock = clock; // @[:@25701.4]
  assign statesInR_0_reset = reset; // @[:@25702.4]
  assign statesInR_0_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@25709.4]
  assign statesInR_0_io_input_enable = _T_143 & _T_148; // @[NBuffers.scala 52:23:@25708.4]
  assign statesInR_1_clock = clock; // @[:@25712.4]
  assign statesInR_1_reset = reset; // @[:@25713.4]
  assign statesInR_1_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@25720.4]
  assign statesInR_1_io_input_enable = _T_143 & _T_148; // @[NBuffers.scala 52:23:@25719.4]
  assign statesInR_2_clock = clock; // @[:@25723.4]
  assign statesInR_2_reset = reset; // @[:@25724.4]
  assign statesInR_2_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@25731.4]
  assign statesInR_2_io_input_enable = _T_143 & _T_148; // @[NBuffers.scala 52:23:@25730.4]
  assign statesInR_3_clock = clock; // @[:@25734.4]
  assign statesInR_3_reset = reset; // @[:@25735.4]
  assign statesInR_3_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@25742.4]
  assign statesInR_3_io_input_enable = _T_143 & _T_148; // @[NBuffers.scala 52:23:@25741.4]
  assign statesInR_4_clock = clock; // @[:@25745.4]
  assign statesInR_4_reset = reset; // @[:@25746.4]
  assign statesInR_4_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@25753.4]
  assign statesInR_4_io_input_enable = _T_143 & _T_148; // @[NBuffers.scala 52:23:@25752.4]
  assign statesInR_5_clock = clock; // @[:@25756.4]
  assign statesInR_5_reset = reset; // @[:@25757.4]
  assign statesInR_5_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@25764.4]
  assign statesInR_5_io_input_enable = _T_143 & _T_148; // @[NBuffers.scala 52:23:@25763.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_148 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_148 <= 1'h0;
    end else begin
      _T_148 <= _T_145;
    end
  end
endmodule
module SRAM_10( // @[:@25906.2]
  input         clock, // @[:@25907.4]
  input         reset, // @[:@25908.4]
  input  [1:0]  io_rPort_0_ofs_0, // @[:@25909.4]
  input         io_rPort_0_en_0, // @[:@25909.4]
  input         io_rPort_0_backpressure, // @[:@25909.4]
  output [31:0] io_rPort_0_output_0, // @[:@25909.4]
  input  [1:0]  io_wPort_1_ofs_0, // @[:@25909.4]
  input  [31:0] io_wPort_1_data_0, // @[:@25909.4]
  input         io_wPort_1_en_0, // @[:@25909.4]
  input  [1:0]  io_wPort_0_ofs_0, // @[:@25909.4]
  input  [31:0] io_wPort_0_data_0, // @[:@25909.4]
  input         io_wPort_0_en_0 // @[:@25909.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@25931.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@25931.4]
  wire [1:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@25931.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@25931.4]
  wire [1:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@25931.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@25931.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@25931.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@25931.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@25961.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@25961.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@25975.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@25975.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@25975.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@25975.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@25975.4]
  wire [34:0] _T_106; // @[Cat.scala 30:58:@25950.4]
  wire [34:0] _T_108; // @[Cat.scala 30:58:@25952.4]
  wire [34:0] _T_109; // @[Mux.scala 31:69:@25953.4]
  wire  _T_115; // @[MemPrimitives.scala 126:35:@25965.4]
  wire [3:0] _T_117; // @[Cat.scala 30:58:@25967.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@25931.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@25961.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@25975.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_106 = {io_wPort_0_en_0,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@25950.4]
  assign _T_108 = {io_wPort_1_en_0,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@25952.4]
  assign _T_109 = io_wPort_0_en_0 ? _T_106 : _T_108; // @[Mux.scala 31:69:@25953.4]
  assign _T_115 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@25965.4]
  assign _T_117 = {_T_115,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@25967.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@25982.4]
  assign Mem1D_clock = clock; // @[:@25932.4]
  assign Mem1D_reset = reset; // @[:@25933.4]
  assign Mem1D_io_r_ofs_0 = _T_117[1:0]; // @[MemPrimitives.scala 131:28:@25971.4]
  assign Mem1D_io_r_backpressure = _T_117[2]; // @[MemPrimitives.scala 132:32:@25972.4]
  assign Mem1D_io_w_ofs_0 = _T_109[1:0]; // @[MemPrimitives.scala 94:28:@25957.4]
  assign Mem1D_io_w_data_0 = _T_109[33:2]; // @[MemPrimitives.scala 95:29:@25958.4]
  assign Mem1D_io_w_en_0 = _T_109[34]; // @[MemPrimitives.scala 96:27:@25959.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@25964.4]
  assign RetimeWrapper_clock = clock; // @[:@25976.4]
  assign RetimeWrapper_reset = reset; // @[:@25977.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@25979.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@25978.4]
endmodule
module x554_tmp_0( // @[:@27069.2]
  input         clock, // @[:@27070.4]
  input         reset, // @[:@27071.4]
  input  [1:0]  io_rPort_0_ofs_0, // @[:@27072.4]
  input         io_rPort_0_en_0, // @[:@27072.4]
  output [31:0] io_rPort_0_output_0, // @[:@27072.4]
  input  [1:0]  io_wPort_1_ofs_0, // @[:@27072.4]
  input  [31:0] io_wPort_1_data_0, // @[:@27072.4]
  input         io_wPort_1_en_0, // @[:@27072.4]
  input  [1:0]  io_wPort_0_ofs_0, // @[:@27072.4]
  input  [31:0] io_wPort_0_data_0, // @[:@27072.4]
  input         io_wPort_0_en_0, // @[:@27072.4]
  input         io_sEn_0, // @[:@27072.4]
  input         io_sEn_1, // @[:@27072.4]
  input         io_sEn_2, // @[:@27072.4]
  input         io_sEn_3, // @[:@27072.4]
  input         io_sEn_4, // @[:@27072.4]
  input         io_sEn_5, // @[:@27072.4]
  input         io_sDone_0, // @[:@27072.4]
  input         io_sDone_1, // @[:@27072.4]
  input         io_sDone_2, // @[:@27072.4]
  input         io_sDone_3, // @[:@27072.4]
  input         io_sDone_4, // @[:@27072.4]
  input         io_sDone_5 // @[:@27072.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@27082.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@27082.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@27082.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@27082.4]
  wire  ctrl_io_sEn_2; // @[NBuffers.scala 83:20:@27082.4]
  wire  ctrl_io_sEn_3; // @[NBuffers.scala 83:20:@27082.4]
  wire  ctrl_io_sEn_4; // @[NBuffers.scala 83:20:@27082.4]
  wire  ctrl_io_sEn_5; // @[NBuffers.scala 83:20:@27082.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@27082.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@27082.4]
  wire  ctrl_io_sDone_2; // @[NBuffers.scala 83:20:@27082.4]
  wire  ctrl_io_sDone_3; // @[NBuffers.scala 83:20:@27082.4]
  wire  ctrl_io_sDone_4; // @[NBuffers.scala 83:20:@27082.4]
  wire  ctrl_io_sDone_5; // @[NBuffers.scala 83:20:@27082.4]
  wire [3:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@27082.4]
  wire [3:0] ctrl_io_statesInW_1; // @[NBuffers.scala 83:20:@27082.4]
  wire [3:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@27082.4]
  wire [3:0] ctrl_io_statesInR_5; // @[NBuffers.scala 83:20:@27082.4]
  wire  SRAM_clock; // @[NBuffers.scala 94:23:@27097.4]
  wire  SRAM_reset; // @[NBuffers.scala 94:23:@27097.4]
  wire [1:0] SRAM_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@27097.4]
  wire  SRAM_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@27097.4]
  wire  SRAM_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@27097.4]
  wire [31:0] SRAM_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@27097.4]
  wire [1:0] SRAM_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@27097.4]
  wire [31:0] SRAM_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@27097.4]
  wire  SRAM_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@27097.4]
  wire [1:0] SRAM_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@27097.4]
  wire [31:0] SRAM_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@27097.4]
  wire  SRAM_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@27097.4]
  wire  SRAM_1_clock; // @[NBuffers.scala 94:23:@27120.4]
  wire  SRAM_1_reset; // @[NBuffers.scala 94:23:@27120.4]
  wire [1:0] SRAM_1_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@27120.4]
  wire  SRAM_1_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@27120.4]
  wire  SRAM_1_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@27120.4]
  wire [31:0] SRAM_1_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@27120.4]
  wire [1:0] SRAM_1_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@27120.4]
  wire [31:0] SRAM_1_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@27120.4]
  wire  SRAM_1_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@27120.4]
  wire [1:0] SRAM_1_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@27120.4]
  wire [31:0] SRAM_1_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@27120.4]
  wire  SRAM_1_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@27120.4]
  wire  SRAM_2_clock; // @[NBuffers.scala 94:23:@27143.4]
  wire  SRAM_2_reset; // @[NBuffers.scala 94:23:@27143.4]
  wire [1:0] SRAM_2_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@27143.4]
  wire  SRAM_2_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@27143.4]
  wire  SRAM_2_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@27143.4]
  wire [31:0] SRAM_2_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@27143.4]
  wire [1:0] SRAM_2_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@27143.4]
  wire [31:0] SRAM_2_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@27143.4]
  wire  SRAM_2_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@27143.4]
  wire [1:0] SRAM_2_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@27143.4]
  wire [31:0] SRAM_2_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@27143.4]
  wire  SRAM_2_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@27143.4]
  wire  SRAM_3_clock; // @[NBuffers.scala 94:23:@27166.4]
  wire  SRAM_3_reset; // @[NBuffers.scala 94:23:@27166.4]
  wire [1:0] SRAM_3_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@27166.4]
  wire  SRAM_3_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@27166.4]
  wire  SRAM_3_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@27166.4]
  wire [31:0] SRAM_3_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@27166.4]
  wire [1:0] SRAM_3_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@27166.4]
  wire [31:0] SRAM_3_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@27166.4]
  wire  SRAM_3_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@27166.4]
  wire [1:0] SRAM_3_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@27166.4]
  wire [31:0] SRAM_3_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@27166.4]
  wire  SRAM_3_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@27166.4]
  wire  SRAM_4_clock; // @[NBuffers.scala 94:23:@27189.4]
  wire  SRAM_4_reset; // @[NBuffers.scala 94:23:@27189.4]
  wire [1:0] SRAM_4_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@27189.4]
  wire  SRAM_4_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@27189.4]
  wire  SRAM_4_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@27189.4]
  wire [31:0] SRAM_4_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@27189.4]
  wire [1:0] SRAM_4_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@27189.4]
  wire [31:0] SRAM_4_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@27189.4]
  wire  SRAM_4_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@27189.4]
  wire [1:0] SRAM_4_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@27189.4]
  wire [31:0] SRAM_4_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@27189.4]
  wire  SRAM_4_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@27189.4]
  wire  SRAM_5_clock; // @[NBuffers.scala 94:23:@27212.4]
  wire  SRAM_5_reset; // @[NBuffers.scala 94:23:@27212.4]
  wire [1:0] SRAM_5_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@27212.4]
  wire  SRAM_5_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@27212.4]
  wire  SRAM_5_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@27212.4]
  wire [31:0] SRAM_5_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@27212.4]
  wire [1:0] SRAM_5_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@27212.4]
  wire [31:0] SRAM_5_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@27212.4]
  wire  SRAM_5_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@27212.4]
  wire [1:0] SRAM_5_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@27212.4]
  wire [31:0] SRAM_5_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@27212.4]
  wire  SRAM_5_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@27212.4]
  wire  _T_148; // @[NBuffers.scala 104:105:@27235.4]
  wire  _T_152; // @[NBuffers.scala 104:105:@27245.4]
  wire  _T_156; // @[NBuffers.scala 108:92:@27255.4]
  wire  _T_159; // @[NBuffers.scala 104:105:@27261.4]
  wire  _T_163; // @[NBuffers.scala 104:105:@27271.4]
  wire  _T_167; // @[NBuffers.scala 108:92:@27281.4]
  wire  _T_170; // @[NBuffers.scala 104:105:@27287.4]
  wire  _T_174; // @[NBuffers.scala 104:105:@27297.4]
  wire  _T_178; // @[NBuffers.scala 108:92:@27307.4]
  wire  _T_181; // @[NBuffers.scala 104:105:@27313.4]
  wire  _T_185; // @[NBuffers.scala 104:105:@27323.4]
  wire  _T_189; // @[NBuffers.scala 108:92:@27333.4]
  wire  _T_192; // @[NBuffers.scala 104:105:@27339.4]
  wire  _T_196; // @[NBuffers.scala 104:105:@27349.4]
  wire  _T_200; // @[NBuffers.scala 108:92:@27359.4]
  wire  _T_203; // @[NBuffers.scala 104:105:@27365.4]
  wire  _T_207; // @[NBuffers.scala 104:105:@27375.4]
  wire  _T_211; // @[NBuffers.scala 108:92:@27385.4]
  wire [31:0] _T_227; // @[Mux.scala 19:72:@27397.4]
  wire [31:0] _T_229; // @[Mux.scala 19:72:@27398.4]
  wire [31:0] _T_231; // @[Mux.scala 19:72:@27399.4]
  wire [31:0] _T_233; // @[Mux.scala 19:72:@27400.4]
  wire [31:0] _T_235; // @[Mux.scala 19:72:@27401.4]
  wire [31:0] _T_237; // @[Mux.scala 19:72:@27402.4]
  wire [31:0] _T_238; // @[Mux.scala 19:72:@27403.4]
  wire [31:0] _T_239; // @[Mux.scala 19:72:@27404.4]
  wire [31:0] _T_240; // @[Mux.scala 19:72:@27405.4]
  wire [31:0] _T_241; // @[Mux.scala 19:72:@27406.4]
  NBufController_5 ctrl ( // @[NBuffers.scala 83:20:@27082.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sEn_2(ctrl_io_sEn_2),
    .io_sEn_3(ctrl_io_sEn_3),
    .io_sEn_4(ctrl_io_sEn_4),
    .io_sEn_5(ctrl_io_sEn_5),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_sDone_2(ctrl_io_sDone_2),
    .io_sDone_3(ctrl_io_sDone_3),
    .io_sDone_4(ctrl_io_sDone_4),
    .io_sDone_5(ctrl_io_sDone_5),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInW_1(ctrl_io_statesInW_1),
    .io_statesInR_1(ctrl_io_statesInR_1),
    .io_statesInR_5(ctrl_io_statesInR_5)
  );
  SRAM_10 SRAM ( // @[NBuffers.scala 94:23:@27097.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_rPort_0_ofs_0(SRAM_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_1 ( // @[NBuffers.scala 94:23:@27120.4]
    .clock(SRAM_1_clock),
    .reset(SRAM_1_reset),
    .io_rPort_0_ofs_0(SRAM_1_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_1_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_1_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_1_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_1_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_1_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_1_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_1_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_1_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_2 ( // @[NBuffers.scala 94:23:@27143.4]
    .clock(SRAM_2_clock),
    .reset(SRAM_2_reset),
    .io_rPort_0_ofs_0(SRAM_2_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_2_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_2_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_2_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_2_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_2_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_2_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_2_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_2_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_2_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_3 ( // @[NBuffers.scala 94:23:@27166.4]
    .clock(SRAM_3_clock),
    .reset(SRAM_3_reset),
    .io_rPort_0_ofs_0(SRAM_3_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_3_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_3_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_3_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_3_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_3_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_3_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_3_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_3_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_3_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_4 ( // @[NBuffers.scala 94:23:@27189.4]
    .clock(SRAM_4_clock),
    .reset(SRAM_4_reset),
    .io_rPort_0_ofs_0(SRAM_4_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_4_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_4_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_4_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_4_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_4_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_4_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_4_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_4_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_4_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_5 ( // @[NBuffers.scala 94:23:@27212.4]
    .clock(SRAM_5_clock),
    .reset(SRAM_5_reset),
    .io_rPort_0_ofs_0(SRAM_5_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_5_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_5_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_5_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_5_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_5_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_5_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_5_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_5_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_5_io_wPort_0_en_0)
  );
  assign _T_148 = ctrl_io_statesInW_0 == 4'h0; // @[NBuffers.scala 104:105:@27235.4]
  assign _T_152 = ctrl_io_statesInW_1 == 4'h0; // @[NBuffers.scala 104:105:@27245.4]
  assign _T_156 = ctrl_io_statesInR_1 == 4'h0; // @[NBuffers.scala 108:92:@27255.4]
  assign _T_159 = ctrl_io_statesInW_0 == 4'h1; // @[NBuffers.scala 104:105:@27261.4]
  assign _T_163 = ctrl_io_statesInW_1 == 4'h1; // @[NBuffers.scala 104:105:@27271.4]
  assign _T_167 = ctrl_io_statesInR_1 == 4'h1; // @[NBuffers.scala 108:92:@27281.4]
  assign _T_170 = ctrl_io_statesInW_0 == 4'h2; // @[NBuffers.scala 104:105:@27287.4]
  assign _T_174 = ctrl_io_statesInW_1 == 4'h2; // @[NBuffers.scala 104:105:@27297.4]
  assign _T_178 = ctrl_io_statesInR_1 == 4'h2; // @[NBuffers.scala 108:92:@27307.4]
  assign _T_181 = ctrl_io_statesInW_0 == 4'h3; // @[NBuffers.scala 104:105:@27313.4]
  assign _T_185 = ctrl_io_statesInW_1 == 4'h3; // @[NBuffers.scala 104:105:@27323.4]
  assign _T_189 = ctrl_io_statesInR_1 == 4'h3; // @[NBuffers.scala 108:92:@27333.4]
  assign _T_192 = ctrl_io_statesInW_0 == 4'h4; // @[NBuffers.scala 104:105:@27339.4]
  assign _T_196 = ctrl_io_statesInW_1 == 4'h4; // @[NBuffers.scala 104:105:@27349.4]
  assign _T_200 = ctrl_io_statesInR_1 == 4'h4; // @[NBuffers.scala 108:92:@27359.4]
  assign _T_203 = ctrl_io_statesInW_0 == 4'h5; // @[NBuffers.scala 104:105:@27365.4]
  assign _T_207 = ctrl_io_statesInW_1 == 4'h5; // @[NBuffers.scala 104:105:@27375.4]
  assign _T_211 = ctrl_io_statesInR_1 == 4'h5; // @[NBuffers.scala 108:92:@27385.4]
  assign _T_227 = _T_156 ? SRAM_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@27397.4]
  assign _T_229 = _T_167 ? SRAM_1_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@27398.4]
  assign _T_231 = _T_178 ? SRAM_2_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@27399.4]
  assign _T_233 = _T_189 ? SRAM_3_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@27400.4]
  assign _T_235 = _T_200 ? SRAM_4_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@27401.4]
  assign _T_237 = _T_211 ? SRAM_5_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@27402.4]
  assign _T_238 = _T_227 | _T_229; // @[Mux.scala 19:72:@27403.4]
  assign _T_239 = _T_238 | _T_231; // @[Mux.scala 19:72:@27404.4]
  assign _T_240 = _T_239 | _T_233; // @[Mux.scala 19:72:@27405.4]
  assign _T_241 = _T_240 | _T_235; // @[Mux.scala 19:72:@27406.4]
  assign io_rPort_0_output_0 = _T_241 | _T_237; // @[NBuffers.scala 115:66:@27410.4]
  assign ctrl_clock = clock; // @[:@27083.4]
  assign ctrl_reset = reset; // @[:@27084.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@27085.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@27087.4]
  assign ctrl_io_sEn_2 = io_sEn_2; // @[NBuffers.scala 85:20:@27089.4]
  assign ctrl_io_sEn_3 = io_sEn_3; // @[NBuffers.scala 85:20:@27091.4]
  assign ctrl_io_sEn_4 = io_sEn_4; // @[NBuffers.scala 85:20:@27093.4]
  assign ctrl_io_sEn_5 = io_sEn_5; // @[NBuffers.scala 85:20:@27095.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@27086.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@27088.4]
  assign ctrl_io_sDone_2 = io_sDone_2; // @[NBuffers.scala 86:22:@27090.4]
  assign ctrl_io_sDone_3 = io_sDone_3; // @[NBuffers.scala 86:22:@27092.4]
  assign ctrl_io_sDone_4 = io_sDone_4; // @[NBuffers.scala 86:22:@27094.4]
  assign ctrl_io_sDone_5 = io_sDone_5; // @[NBuffers.scala 86:22:@27096.4]
  assign SRAM_clock = clock; // @[:@27098.4]
  assign SRAM_reset = reset; // @[:@27099.4]
  assign SRAM_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@27257.4]
  assign SRAM_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_156; // @[MemPrimitives.scala 43:33:@27259.4]
  assign SRAM_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@27260.4]
  assign SRAM_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@27247.4]
  assign SRAM_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@27248.4]
  assign SRAM_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_152; // @[MemPrimitives.scala 37:29:@27254.4]
  assign SRAM_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@27237.4]
  assign SRAM_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@27238.4]
  assign SRAM_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_148; // @[MemPrimitives.scala 37:29:@27244.4]
  assign SRAM_1_clock = clock; // @[:@27121.4]
  assign SRAM_1_reset = reset; // @[:@27122.4]
  assign SRAM_1_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@27283.4]
  assign SRAM_1_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_167; // @[MemPrimitives.scala 43:33:@27285.4]
  assign SRAM_1_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@27286.4]
  assign SRAM_1_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@27273.4]
  assign SRAM_1_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@27274.4]
  assign SRAM_1_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_163; // @[MemPrimitives.scala 37:29:@27280.4]
  assign SRAM_1_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@27263.4]
  assign SRAM_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@27264.4]
  assign SRAM_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_159; // @[MemPrimitives.scala 37:29:@27270.4]
  assign SRAM_2_clock = clock; // @[:@27144.4]
  assign SRAM_2_reset = reset; // @[:@27145.4]
  assign SRAM_2_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@27309.4]
  assign SRAM_2_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_178; // @[MemPrimitives.scala 43:33:@27311.4]
  assign SRAM_2_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@27312.4]
  assign SRAM_2_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@27299.4]
  assign SRAM_2_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@27300.4]
  assign SRAM_2_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_174; // @[MemPrimitives.scala 37:29:@27306.4]
  assign SRAM_2_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@27289.4]
  assign SRAM_2_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@27290.4]
  assign SRAM_2_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_170; // @[MemPrimitives.scala 37:29:@27296.4]
  assign SRAM_3_clock = clock; // @[:@27167.4]
  assign SRAM_3_reset = reset; // @[:@27168.4]
  assign SRAM_3_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@27335.4]
  assign SRAM_3_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_189; // @[MemPrimitives.scala 43:33:@27337.4]
  assign SRAM_3_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@27338.4]
  assign SRAM_3_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@27325.4]
  assign SRAM_3_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@27326.4]
  assign SRAM_3_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_185; // @[MemPrimitives.scala 37:29:@27332.4]
  assign SRAM_3_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@27315.4]
  assign SRAM_3_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@27316.4]
  assign SRAM_3_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_181; // @[MemPrimitives.scala 37:29:@27322.4]
  assign SRAM_4_clock = clock; // @[:@27190.4]
  assign SRAM_4_reset = reset; // @[:@27191.4]
  assign SRAM_4_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@27361.4]
  assign SRAM_4_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_200; // @[MemPrimitives.scala 43:33:@27363.4]
  assign SRAM_4_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@27364.4]
  assign SRAM_4_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@27351.4]
  assign SRAM_4_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@27352.4]
  assign SRAM_4_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_196; // @[MemPrimitives.scala 37:29:@27358.4]
  assign SRAM_4_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@27341.4]
  assign SRAM_4_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@27342.4]
  assign SRAM_4_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_192; // @[MemPrimitives.scala 37:29:@27348.4]
  assign SRAM_5_clock = clock; // @[:@27213.4]
  assign SRAM_5_reset = reset; // @[:@27214.4]
  assign SRAM_5_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@27387.4]
  assign SRAM_5_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_211; // @[MemPrimitives.scala 43:33:@27389.4]
  assign SRAM_5_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@27390.4]
  assign SRAM_5_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@27377.4]
  assign SRAM_5_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@27378.4]
  assign SRAM_5_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_207; // @[MemPrimitives.scala 37:29:@27384.4]
  assign SRAM_5_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@27367.4]
  assign SRAM_5_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@27368.4]
  assign SRAM_5_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_203; // @[MemPrimitives.scala 37:29:@27374.4]
endmodule
module x557_tmp_3( // @[:@37872.2]
  input         clock, // @[:@37873.4]
  input         reset, // @[:@37874.4]
  input  [1:0]  io_rPort_0_ofs_0, // @[:@37875.4]
  input         io_rPort_0_en_0, // @[:@37875.4]
  output [31:0] io_rPort_0_output_0, // @[:@37875.4]
  input  [1:0]  io_wPort_1_ofs_0, // @[:@37875.4]
  input  [31:0] io_wPort_1_data_0, // @[:@37875.4]
  input         io_wPort_1_en_0, // @[:@37875.4]
  input  [1:0]  io_wPort_0_ofs_0, // @[:@37875.4]
  input  [31:0] io_wPort_0_data_0, // @[:@37875.4]
  input         io_wPort_0_en_0, // @[:@37875.4]
  input         io_sEn_0, // @[:@37875.4]
  input         io_sEn_1, // @[:@37875.4]
  input         io_sEn_2, // @[:@37875.4]
  input         io_sEn_3, // @[:@37875.4]
  input         io_sEn_4, // @[:@37875.4]
  input         io_sEn_5, // @[:@37875.4]
  input         io_sDone_0, // @[:@37875.4]
  input         io_sDone_1, // @[:@37875.4]
  input         io_sDone_2, // @[:@37875.4]
  input         io_sDone_3, // @[:@37875.4]
  input         io_sDone_4, // @[:@37875.4]
  input         io_sDone_5 // @[:@37875.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@37885.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@37885.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@37885.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@37885.4]
  wire  ctrl_io_sEn_2; // @[NBuffers.scala 83:20:@37885.4]
  wire  ctrl_io_sEn_3; // @[NBuffers.scala 83:20:@37885.4]
  wire  ctrl_io_sEn_4; // @[NBuffers.scala 83:20:@37885.4]
  wire  ctrl_io_sEn_5; // @[NBuffers.scala 83:20:@37885.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@37885.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@37885.4]
  wire  ctrl_io_sDone_2; // @[NBuffers.scala 83:20:@37885.4]
  wire  ctrl_io_sDone_3; // @[NBuffers.scala 83:20:@37885.4]
  wire  ctrl_io_sDone_4; // @[NBuffers.scala 83:20:@37885.4]
  wire  ctrl_io_sDone_5; // @[NBuffers.scala 83:20:@37885.4]
  wire [3:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@37885.4]
  wire [3:0] ctrl_io_statesInW_1; // @[NBuffers.scala 83:20:@37885.4]
  wire [3:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@37885.4]
  wire [3:0] ctrl_io_statesInR_5; // @[NBuffers.scala 83:20:@37885.4]
  wire  SRAM_clock; // @[NBuffers.scala 94:23:@37900.4]
  wire  SRAM_reset; // @[NBuffers.scala 94:23:@37900.4]
  wire [1:0] SRAM_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@37900.4]
  wire  SRAM_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@37900.4]
  wire  SRAM_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@37900.4]
  wire [31:0] SRAM_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@37900.4]
  wire [1:0] SRAM_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@37900.4]
  wire [31:0] SRAM_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@37900.4]
  wire  SRAM_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@37900.4]
  wire [1:0] SRAM_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@37900.4]
  wire [31:0] SRAM_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@37900.4]
  wire  SRAM_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@37900.4]
  wire  SRAM_1_clock; // @[NBuffers.scala 94:23:@37923.4]
  wire  SRAM_1_reset; // @[NBuffers.scala 94:23:@37923.4]
  wire [1:0] SRAM_1_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@37923.4]
  wire  SRAM_1_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@37923.4]
  wire  SRAM_1_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@37923.4]
  wire [31:0] SRAM_1_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@37923.4]
  wire [1:0] SRAM_1_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@37923.4]
  wire [31:0] SRAM_1_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@37923.4]
  wire  SRAM_1_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@37923.4]
  wire [1:0] SRAM_1_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@37923.4]
  wire [31:0] SRAM_1_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@37923.4]
  wire  SRAM_1_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@37923.4]
  wire  SRAM_2_clock; // @[NBuffers.scala 94:23:@37946.4]
  wire  SRAM_2_reset; // @[NBuffers.scala 94:23:@37946.4]
  wire [1:0] SRAM_2_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@37946.4]
  wire  SRAM_2_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@37946.4]
  wire  SRAM_2_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@37946.4]
  wire [31:0] SRAM_2_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@37946.4]
  wire [1:0] SRAM_2_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@37946.4]
  wire [31:0] SRAM_2_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@37946.4]
  wire  SRAM_2_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@37946.4]
  wire [1:0] SRAM_2_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@37946.4]
  wire [31:0] SRAM_2_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@37946.4]
  wire  SRAM_2_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@37946.4]
  wire  SRAM_3_clock; // @[NBuffers.scala 94:23:@37969.4]
  wire  SRAM_3_reset; // @[NBuffers.scala 94:23:@37969.4]
  wire [1:0] SRAM_3_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@37969.4]
  wire  SRAM_3_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@37969.4]
  wire  SRAM_3_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@37969.4]
  wire [31:0] SRAM_3_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@37969.4]
  wire [1:0] SRAM_3_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@37969.4]
  wire [31:0] SRAM_3_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@37969.4]
  wire  SRAM_3_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@37969.4]
  wire [1:0] SRAM_3_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@37969.4]
  wire [31:0] SRAM_3_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@37969.4]
  wire  SRAM_3_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@37969.4]
  wire  SRAM_4_clock; // @[NBuffers.scala 94:23:@37992.4]
  wire  SRAM_4_reset; // @[NBuffers.scala 94:23:@37992.4]
  wire [1:0] SRAM_4_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@37992.4]
  wire  SRAM_4_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@37992.4]
  wire  SRAM_4_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@37992.4]
  wire [31:0] SRAM_4_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@37992.4]
  wire [1:0] SRAM_4_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@37992.4]
  wire [31:0] SRAM_4_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@37992.4]
  wire  SRAM_4_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@37992.4]
  wire [1:0] SRAM_4_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@37992.4]
  wire [31:0] SRAM_4_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@37992.4]
  wire  SRAM_4_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@37992.4]
  wire  SRAM_5_clock; // @[NBuffers.scala 94:23:@38015.4]
  wire  SRAM_5_reset; // @[NBuffers.scala 94:23:@38015.4]
  wire [1:0] SRAM_5_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@38015.4]
  wire  SRAM_5_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@38015.4]
  wire  SRAM_5_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@38015.4]
  wire [31:0] SRAM_5_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@38015.4]
  wire [1:0] SRAM_5_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@38015.4]
  wire [31:0] SRAM_5_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@38015.4]
  wire  SRAM_5_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@38015.4]
  wire [1:0] SRAM_5_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@38015.4]
  wire [31:0] SRAM_5_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@38015.4]
  wire  SRAM_5_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@38015.4]
  wire  _T_148; // @[NBuffers.scala 104:105:@38038.4]
  wire  _T_152; // @[NBuffers.scala 104:105:@38048.4]
  wire  _T_156; // @[NBuffers.scala 108:92:@38058.4]
  wire  _T_159; // @[NBuffers.scala 104:105:@38064.4]
  wire  _T_163; // @[NBuffers.scala 104:105:@38074.4]
  wire  _T_167; // @[NBuffers.scala 108:92:@38084.4]
  wire  _T_170; // @[NBuffers.scala 104:105:@38090.4]
  wire  _T_174; // @[NBuffers.scala 104:105:@38100.4]
  wire  _T_178; // @[NBuffers.scala 108:92:@38110.4]
  wire  _T_181; // @[NBuffers.scala 104:105:@38116.4]
  wire  _T_185; // @[NBuffers.scala 104:105:@38126.4]
  wire  _T_189; // @[NBuffers.scala 108:92:@38136.4]
  wire  _T_192; // @[NBuffers.scala 104:105:@38142.4]
  wire  _T_196; // @[NBuffers.scala 104:105:@38152.4]
  wire  _T_200; // @[NBuffers.scala 108:92:@38162.4]
  wire  _T_203; // @[NBuffers.scala 104:105:@38168.4]
  wire  _T_207; // @[NBuffers.scala 104:105:@38178.4]
  wire  _T_211; // @[NBuffers.scala 108:92:@38188.4]
  wire [31:0] _T_227; // @[Mux.scala 19:72:@38200.4]
  wire [31:0] _T_229; // @[Mux.scala 19:72:@38201.4]
  wire [31:0] _T_231; // @[Mux.scala 19:72:@38202.4]
  wire [31:0] _T_233; // @[Mux.scala 19:72:@38203.4]
  wire [31:0] _T_235; // @[Mux.scala 19:72:@38204.4]
  wire [31:0] _T_237; // @[Mux.scala 19:72:@38205.4]
  wire [31:0] _T_238; // @[Mux.scala 19:72:@38206.4]
  wire [31:0] _T_239; // @[Mux.scala 19:72:@38207.4]
  wire [31:0] _T_240; // @[Mux.scala 19:72:@38208.4]
  wire [31:0] _T_241; // @[Mux.scala 19:72:@38209.4]
  NBufController_5 ctrl ( // @[NBuffers.scala 83:20:@37885.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sEn_2(ctrl_io_sEn_2),
    .io_sEn_3(ctrl_io_sEn_3),
    .io_sEn_4(ctrl_io_sEn_4),
    .io_sEn_5(ctrl_io_sEn_5),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_sDone_2(ctrl_io_sDone_2),
    .io_sDone_3(ctrl_io_sDone_3),
    .io_sDone_4(ctrl_io_sDone_4),
    .io_sDone_5(ctrl_io_sDone_5),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInW_1(ctrl_io_statesInW_1),
    .io_statesInR_1(ctrl_io_statesInR_1),
    .io_statesInR_5(ctrl_io_statesInR_5)
  );
  SRAM_10 SRAM ( // @[NBuffers.scala 94:23:@37900.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_rPort_0_ofs_0(SRAM_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_1 ( // @[NBuffers.scala 94:23:@37923.4]
    .clock(SRAM_1_clock),
    .reset(SRAM_1_reset),
    .io_rPort_0_ofs_0(SRAM_1_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_1_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_1_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_1_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_1_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_1_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_1_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_1_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_1_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_2 ( // @[NBuffers.scala 94:23:@37946.4]
    .clock(SRAM_2_clock),
    .reset(SRAM_2_reset),
    .io_rPort_0_ofs_0(SRAM_2_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_2_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_2_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_2_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_2_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_2_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_2_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_2_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_2_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_2_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_3 ( // @[NBuffers.scala 94:23:@37969.4]
    .clock(SRAM_3_clock),
    .reset(SRAM_3_reset),
    .io_rPort_0_ofs_0(SRAM_3_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_3_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_3_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_3_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_3_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_3_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_3_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_3_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_3_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_3_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_4 ( // @[NBuffers.scala 94:23:@37992.4]
    .clock(SRAM_4_clock),
    .reset(SRAM_4_reset),
    .io_rPort_0_ofs_0(SRAM_4_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_4_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_4_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_4_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_4_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_4_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_4_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_4_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_4_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_4_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_5 ( // @[NBuffers.scala 94:23:@38015.4]
    .clock(SRAM_5_clock),
    .reset(SRAM_5_reset),
    .io_rPort_0_ofs_0(SRAM_5_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_5_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_5_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_5_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_5_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_5_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_5_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_5_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_5_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_5_io_wPort_0_en_0)
  );
  assign _T_148 = ctrl_io_statesInW_0 == 4'h0; // @[NBuffers.scala 104:105:@38038.4]
  assign _T_152 = ctrl_io_statesInW_1 == 4'h0; // @[NBuffers.scala 104:105:@38048.4]
  assign _T_156 = ctrl_io_statesInR_5 == 4'h0; // @[NBuffers.scala 108:92:@38058.4]
  assign _T_159 = ctrl_io_statesInW_0 == 4'h1; // @[NBuffers.scala 104:105:@38064.4]
  assign _T_163 = ctrl_io_statesInW_1 == 4'h1; // @[NBuffers.scala 104:105:@38074.4]
  assign _T_167 = ctrl_io_statesInR_5 == 4'h1; // @[NBuffers.scala 108:92:@38084.4]
  assign _T_170 = ctrl_io_statesInW_0 == 4'h2; // @[NBuffers.scala 104:105:@38090.4]
  assign _T_174 = ctrl_io_statesInW_1 == 4'h2; // @[NBuffers.scala 104:105:@38100.4]
  assign _T_178 = ctrl_io_statesInR_5 == 4'h2; // @[NBuffers.scala 108:92:@38110.4]
  assign _T_181 = ctrl_io_statesInW_0 == 4'h3; // @[NBuffers.scala 104:105:@38116.4]
  assign _T_185 = ctrl_io_statesInW_1 == 4'h3; // @[NBuffers.scala 104:105:@38126.4]
  assign _T_189 = ctrl_io_statesInR_5 == 4'h3; // @[NBuffers.scala 108:92:@38136.4]
  assign _T_192 = ctrl_io_statesInW_0 == 4'h4; // @[NBuffers.scala 104:105:@38142.4]
  assign _T_196 = ctrl_io_statesInW_1 == 4'h4; // @[NBuffers.scala 104:105:@38152.4]
  assign _T_200 = ctrl_io_statesInR_5 == 4'h4; // @[NBuffers.scala 108:92:@38162.4]
  assign _T_203 = ctrl_io_statesInW_0 == 4'h5; // @[NBuffers.scala 104:105:@38168.4]
  assign _T_207 = ctrl_io_statesInW_1 == 4'h5; // @[NBuffers.scala 104:105:@38178.4]
  assign _T_211 = ctrl_io_statesInR_5 == 4'h5; // @[NBuffers.scala 108:92:@38188.4]
  assign _T_227 = _T_156 ? SRAM_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@38200.4]
  assign _T_229 = _T_167 ? SRAM_1_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@38201.4]
  assign _T_231 = _T_178 ? SRAM_2_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@38202.4]
  assign _T_233 = _T_189 ? SRAM_3_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@38203.4]
  assign _T_235 = _T_200 ? SRAM_4_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@38204.4]
  assign _T_237 = _T_211 ? SRAM_5_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@38205.4]
  assign _T_238 = _T_227 | _T_229; // @[Mux.scala 19:72:@38206.4]
  assign _T_239 = _T_238 | _T_231; // @[Mux.scala 19:72:@38207.4]
  assign _T_240 = _T_239 | _T_233; // @[Mux.scala 19:72:@38208.4]
  assign _T_241 = _T_240 | _T_235; // @[Mux.scala 19:72:@38209.4]
  assign io_rPort_0_output_0 = _T_241 | _T_237; // @[NBuffers.scala 115:66:@38213.4]
  assign ctrl_clock = clock; // @[:@37886.4]
  assign ctrl_reset = reset; // @[:@37887.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@37888.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@37890.4]
  assign ctrl_io_sEn_2 = io_sEn_2; // @[NBuffers.scala 85:20:@37892.4]
  assign ctrl_io_sEn_3 = io_sEn_3; // @[NBuffers.scala 85:20:@37894.4]
  assign ctrl_io_sEn_4 = io_sEn_4; // @[NBuffers.scala 85:20:@37896.4]
  assign ctrl_io_sEn_5 = io_sEn_5; // @[NBuffers.scala 85:20:@37898.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@37889.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@37891.4]
  assign ctrl_io_sDone_2 = io_sDone_2; // @[NBuffers.scala 86:22:@37893.4]
  assign ctrl_io_sDone_3 = io_sDone_3; // @[NBuffers.scala 86:22:@37895.4]
  assign ctrl_io_sDone_4 = io_sDone_4; // @[NBuffers.scala 86:22:@37897.4]
  assign ctrl_io_sDone_5 = io_sDone_5; // @[NBuffers.scala 86:22:@37899.4]
  assign SRAM_clock = clock; // @[:@37901.4]
  assign SRAM_reset = reset; // @[:@37902.4]
  assign SRAM_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@38060.4]
  assign SRAM_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_156; // @[MemPrimitives.scala 43:33:@38062.4]
  assign SRAM_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@38063.4]
  assign SRAM_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@38050.4]
  assign SRAM_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@38051.4]
  assign SRAM_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_152; // @[MemPrimitives.scala 37:29:@38057.4]
  assign SRAM_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@38040.4]
  assign SRAM_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@38041.4]
  assign SRAM_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_148; // @[MemPrimitives.scala 37:29:@38047.4]
  assign SRAM_1_clock = clock; // @[:@37924.4]
  assign SRAM_1_reset = reset; // @[:@37925.4]
  assign SRAM_1_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@38086.4]
  assign SRAM_1_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_167; // @[MemPrimitives.scala 43:33:@38088.4]
  assign SRAM_1_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@38089.4]
  assign SRAM_1_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@38076.4]
  assign SRAM_1_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@38077.4]
  assign SRAM_1_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_163; // @[MemPrimitives.scala 37:29:@38083.4]
  assign SRAM_1_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@38066.4]
  assign SRAM_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@38067.4]
  assign SRAM_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_159; // @[MemPrimitives.scala 37:29:@38073.4]
  assign SRAM_2_clock = clock; // @[:@37947.4]
  assign SRAM_2_reset = reset; // @[:@37948.4]
  assign SRAM_2_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@38112.4]
  assign SRAM_2_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_178; // @[MemPrimitives.scala 43:33:@38114.4]
  assign SRAM_2_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@38115.4]
  assign SRAM_2_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@38102.4]
  assign SRAM_2_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@38103.4]
  assign SRAM_2_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_174; // @[MemPrimitives.scala 37:29:@38109.4]
  assign SRAM_2_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@38092.4]
  assign SRAM_2_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@38093.4]
  assign SRAM_2_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_170; // @[MemPrimitives.scala 37:29:@38099.4]
  assign SRAM_3_clock = clock; // @[:@37970.4]
  assign SRAM_3_reset = reset; // @[:@37971.4]
  assign SRAM_3_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@38138.4]
  assign SRAM_3_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_189; // @[MemPrimitives.scala 43:33:@38140.4]
  assign SRAM_3_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@38141.4]
  assign SRAM_3_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@38128.4]
  assign SRAM_3_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@38129.4]
  assign SRAM_3_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_185; // @[MemPrimitives.scala 37:29:@38135.4]
  assign SRAM_3_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@38118.4]
  assign SRAM_3_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@38119.4]
  assign SRAM_3_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_181; // @[MemPrimitives.scala 37:29:@38125.4]
  assign SRAM_4_clock = clock; // @[:@37993.4]
  assign SRAM_4_reset = reset; // @[:@37994.4]
  assign SRAM_4_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@38164.4]
  assign SRAM_4_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_200; // @[MemPrimitives.scala 43:33:@38166.4]
  assign SRAM_4_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@38167.4]
  assign SRAM_4_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@38154.4]
  assign SRAM_4_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@38155.4]
  assign SRAM_4_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_196; // @[MemPrimitives.scala 37:29:@38161.4]
  assign SRAM_4_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@38144.4]
  assign SRAM_4_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@38145.4]
  assign SRAM_4_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_192; // @[MemPrimitives.scala 37:29:@38151.4]
  assign SRAM_5_clock = clock; // @[:@38016.4]
  assign SRAM_5_reset = reset; // @[:@38017.4]
  assign SRAM_5_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@38190.4]
  assign SRAM_5_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_211; // @[MemPrimitives.scala 43:33:@38192.4]
  assign SRAM_5_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@38193.4]
  assign SRAM_5_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@38180.4]
  assign SRAM_5_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@38181.4]
  assign SRAM_5_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_207; // @[MemPrimitives.scala 37:29:@38187.4]
  assign SRAM_5_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@38170.4]
  assign SRAM_5_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@38171.4]
  assign SRAM_5_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_203; // @[MemPrimitives.scala 37:29:@38177.4]
endmodule
module NBufController_9( // @[:@40031.2]
  input        clock, // @[:@40032.4]
  input        reset, // @[:@40033.4]
  input        io_sEn_0, // @[:@40034.4]
  input        io_sEn_1, // @[:@40034.4]
  input        io_sEn_2, // @[:@40034.4]
  input        io_sEn_3, // @[:@40034.4]
  input        io_sEn_4, // @[:@40034.4]
  input        io_sEn_5, // @[:@40034.4]
  input        io_sEn_6, // @[:@40034.4]
  input        io_sDone_0, // @[:@40034.4]
  input        io_sDone_1, // @[:@40034.4]
  input        io_sDone_2, // @[:@40034.4]
  input        io_sDone_3, // @[:@40034.4]
  input        io_sDone_4, // @[:@40034.4]
  input        io_sDone_5, // @[:@40034.4]
  input        io_sDone_6, // @[:@40034.4]
  output [3:0] io_statesInW_0, // @[:@40034.4]
  output [3:0] io_statesInW_1, // @[:@40034.4]
  output [3:0] io_statesInR_6 // @[:@40034.4]
);
  wire  sEn_latch_0_clock; // @[NBuffers.scala 21:52:@40036.4]
  wire  sEn_latch_0_reset; // @[NBuffers.scala 21:52:@40036.4]
  wire  sEn_latch_0_io_input_set; // @[NBuffers.scala 21:52:@40036.4]
  wire  sEn_latch_0_io_input_reset; // @[NBuffers.scala 21:52:@40036.4]
  wire  sEn_latch_0_io_input_asyn_reset; // @[NBuffers.scala 21:52:@40036.4]
  wire  sEn_latch_0_io_output; // @[NBuffers.scala 21:52:@40036.4]
  wire  sEn_latch_1_clock; // @[NBuffers.scala 21:52:@40039.4]
  wire  sEn_latch_1_reset; // @[NBuffers.scala 21:52:@40039.4]
  wire  sEn_latch_1_io_input_set; // @[NBuffers.scala 21:52:@40039.4]
  wire  sEn_latch_1_io_input_reset; // @[NBuffers.scala 21:52:@40039.4]
  wire  sEn_latch_1_io_input_asyn_reset; // @[NBuffers.scala 21:52:@40039.4]
  wire  sEn_latch_1_io_output; // @[NBuffers.scala 21:52:@40039.4]
  wire  sEn_latch_2_clock; // @[NBuffers.scala 21:52:@40042.4]
  wire  sEn_latch_2_reset; // @[NBuffers.scala 21:52:@40042.4]
  wire  sEn_latch_2_io_input_set; // @[NBuffers.scala 21:52:@40042.4]
  wire  sEn_latch_2_io_input_reset; // @[NBuffers.scala 21:52:@40042.4]
  wire  sEn_latch_2_io_input_asyn_reset; // @[NBuffers.scala 21:52:@40042.4]
  wire  sEn_latch_2_io_output; // @[NBuffers.scala 21:52:@40042.4]
  wire  sEn_latch_3_clock; // @[NBuffers.scala 21:52:@40045.4]
  wire  sEn_latch_3_reset; // @[NBuffers.scala 21:52:@40045.4]
  wire  sEn_latch_3_io_input_set; // @[NBuffers.scala 21:52:@40045.4]
  wire  sEn_latch_3_io_input_reset; // @[NBuffers.scala 21:52:@40045.4]
  wire  sEn_latch_3_io_input_asyn_reset; // @[NBuffers.scala 21:52:@40045.4]
  wire  sEn_latch_3_io_output; // @[NBuffers.scala 21:52:@40045.4]
  wire  sEn_latch_4_clock; // @[NBuffers.scala 21:52:@40048.4]
  wire  sEn_latch_4_reset; // @[NBuffers.scala 21:52:@40048.4]
  wire  sEn_latch_4_io_input_set; // @[NBuffers.scala 21:52:@40048.4]
  wire  sEn_latch_4_io_input_reset; // @[NBuffers.scala 21:52:@40048.4]
  wire  sEn_latch_4_io_input_asyn_reset; // @[NBuffers.scala 21:52:@40048.4]
  wire  sEn_latch_4_io_output; // @[NBuffers.scala 21:52:@40048.4]
  wire  sEn_latch_5_clock; // @[NBuffers.scala 21:52:@40051.4]
  wire  sEn_latch_5_reset; // @[NBuffers.scala 21:52:@40051.4]
  wire  sEn_latch_5_io_input_set; // @[NBuffers.scala 21:52:@40051.4]
  wire  sEn_latch_5_io_input_reset; // @[NBuffers.scala 21:52:@40051.4]
  wire  sEn_latch_5_io_input_asyn_reset; // @[NBuffers.scala 21:52:@40051.4]
  wire  sEn_latch_5_io_output; // @[NBuffers.scala 21:52:@40051.4]
  wire  sEn_latch_6_clock; // @[NBuffers.scala 21:52:@40054.4]
  wire  sEn_latch_6_reset; // @[NBuffers.scala 21:52:@40054.4]
  wire  sEn_latch_6_io_input_set; // @[NBuffers.scala 21:52:@40054.4]
  wire  sEn_latch_6_io_input_reset; // @[NBuffers.scala 21:52:@40054.4]
  wire  sEn_latch_6_io_input_asyn_reset; // @[NBuffers.scala 21:52:@40054.4]
  wire  sEn_latch_6_io_output; // @[NBuffers.scala 21:52:@40054.4]
  wire  sDone_latch_0_clock; // @[NBuffers.scala 22:54:@40057.4]
  wire  sDone_latch_0_reset; // @[NBuffers.scala 22:54:@40057.4]
  wire  sDone_latch_0_io_input_set; // @[NBuffers.scala 22:54:@40057.4]
  wire  sDone_latch_0_io_input_reset; // @[NBuffers.scala 22:54:@40057.4]
  wire  sDone_latch_0_io_input_asyn_reset; // @[NBuffers.scala 22:54:@40057.4]
  wire  sDone_latch_0_io_output; // @[NBuffers.scala 22:54:@40057.4]
  wire  sDone_latch_1_clock; // @[NBuffers.scala 22:54:@40060.4]
  wire  sDone_latch_1_reset; // @[NBuffers.scala 22:54:@40060.4]
  wire  sDone_latch_1_io_input_set; // @[NBuffers.scala 22:54:@40060.4]
  wire  sDone_latch_1_io_input_reset; // @[NBuffers.scala 22:54:@40060.4]
  wire  sDone_latch_1_io_input_asyn_reset; // @[NBuffers.scala 22:54:@40060.4]
  wire  sDone_latch_1_io_output; // @[NBuffers.scala 22:54:@40060.4]
  wire  sDone_latch_2_clock; // @[NBuffers.scala 22:54:@40063.4]
  wire  sDone_latch_2_reset; // @[NBuffers.scala 22:54:@40063.4]
  wire  sDone_latch_2_io_input_set; // @[NBuffers.scala 22:54:@40063.4]
  wire  sDone_latch_2_io_input_reset; // @[NBuffers.scala 22:54:@40063.4]
  wire  sDone_latch_2_io_input_asyn_reset; // @[NBuffers.scala 22:54:@40063.4]
  wire  sDone_latch_2_io_output; // @[NBuffers.scala 22:54:@40063.4]
  wire  sDone_latch_3_clock; // @[NBuffers.scala 22:54:@40066.4]
  wire  sDone_latch_3_reset; // @[NBuffers.scala 22:54:@40066.4]
  wire  sDone_latch_3_io_input_set; // @[NBuffers.scala 22:54:@40066.4]
  wire  sDone_latch_3_io_input_reset; // @[NBuffers.scala 22:54:@40066.4]
  wire  sDone_latch_3_io_input_asyn_reset; // @[NBuffers.scala 22:54:@40066.4]
  wire  sDone_latch_3_io_output; // @[NBuffers.scala 22:54:@40066.4]
  wire  sDone_latch_4_clock; // @[NBuffers.scala 22:54:@40069.4]
  wire  sDone_latch_4_reset; // @[NBuffers.scala 22:54:@40069.4]
  wire  sDone_latch_4_io_input_set; // @[NBuffers.scala 22:54:@40069.4]
  wire  sDone_latch_4_io_input_reset; // @[NBuffers.scala 22:54:@40069.4]
  wire  sDone_latch_4_io_input_asyn_reset; // @[NBuffers.scala 22:54:@40069.4]
  wire  sDone_latch_4_io_output; // @[NBuffers.scala 22:54:@40069.4]
  wire  sDone_latch_5_clock; // @[NBuffers.scala 22:54:@40072.4]
  wire  sDone_latch_5_reset; // @[NBuffers.scala 22:54:@40072.4]
  wire  sDone_latch_5_io_input_set; // @[NBuffers.scala 22:54:@40072.4]
  wire  sDone_latch_5_io_input_reset; // @[NBuffers.scala 22:54:@40072.4]
  wire  sDone_latch_5_io_input_asyn_reset; // @[NBuffers.scala 22:54:@40072.4]
  wire  sDone_latch_5_io_output; // @[NBuffers.scala 22:54:@40072.4]
  wire  sDone_latch_6_clock; // @[NBuffers.scala 22:54:@40075.4]
  wire  sDone_latch_6_reset; // @[NBuffers.scala 22:54:@40075.4]
  wire  sDone_latch_6_io_input_set; // @[NBuffers.scala 22:54:@40075.4]
  wire  sDone_latch_6_io_input_reset; // @[NBuffers.scala 22:54:@40075.4]
  wire  sDone_latch_6_io_input_asyn_reset; // @[NBuffers.scala 22:54:@40075.4]
  wire  sDone_latch_6_io_output; // @[NBuffers.scala 22:54:@40075.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@40082.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@40082.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@40082.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@40082.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@40082.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@40090.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@40090.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@40090.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@40090.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@40090.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@40099.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@40099.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@40099.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@40099.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@40099.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@40107.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@40107.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@40107.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@40107.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@40107.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@40118.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@40118.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@40118.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@40118.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@40118.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@40126.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@40126.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@40126.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@40126.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@40126.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@40135.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@40135.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@40135.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@40135.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@40135.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@40143.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@40143.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@40143.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@40143.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@40143.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@40154.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@40154.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@40154.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@40154.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@40154.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@40162.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@40162.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@40162.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@40162.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@40162.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@40171.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@40171.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@40171.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@40171.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@40171.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@40179.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@40179.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@40179.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@40179.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@40179.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@40190.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@40190.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@40190.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@40190.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@40190.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@40198.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@40198.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@40198.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@40198.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@40198.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@40207.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@40207.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@40207.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@40207.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@40207.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@40215.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@40215.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@40215.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@40215.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@40215.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@40226.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@40226.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@40226.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@40226.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@40226.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@40234.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@40234.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@40234.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@40234.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@40234.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@40243.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@40243.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@40243.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@40243.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@40243.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@40251.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@40251.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@40251.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@40251.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@40251.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@40262.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@40262.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@40262.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@40262.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@40262.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@40270.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@40270.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@40270.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@40270.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@40270.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@40279.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@40279.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@40279.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@40279.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@40279.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@40287.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@40287.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@40287.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@40287.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@40287.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@40298.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@40298.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@40298.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@40298.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@40298.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@40306.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@40306.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@40306.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@40306.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@40306.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@40315.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@40315.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@40315.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@40315.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@40315.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@40323.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@40323.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@40323.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@40323.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@40323.4]
  wire  NBufCtr_clock; // @[NBuffers.scala 40:19:@40364.4]
  wire  NBufCtr_reset; // @[NBuffers.scala 40:19:@40364.4]
  wire  NBufCtr_io_input_countUp; // @[NBuffers.scala 40:19:@40364.4]
  wire  NBufCtr_io_input_enable; // @[NBuffers.scala 40:19:@40364.4]
  wire [31:0] NBufCtr_io_output_count; // @[NBuffers.scala 40:19:@40364.4]
  wire  NBufCtr_1_clock; // @[NBuffers.scala 40:19:@40375.4]
  wire  NBufCtr_1_reset; // @[NBuffers.scala 40:19:@40375.4]
  wire  NBufCtr_1_io_input_countUp; // @[NBuffers.scala 40:19:@40375.4]
  wire  NBufCtr_1_io_input_enable; // @[NBuffers.scala 40:19:@40375.4]
  wire [31:0] NBufCtr_1_io_output_count; // @[NBuffers.scala 40:19:@40375.4]
  wire  statesInR_0_clock; // @[NBuffers.scala 50:19:@40386.4]
  wire  statesInR_0_reset; // @[NBuffers.scala 50:19:@40386.4]
  wire  statesInR_0_io_input_countUp; // @[NBuffers.scala 50:19:@40386.4]
  wire  statesInR_0_io_input_enable; // @[NBuffers.scala 50:19:@40386.4]
  wire [31:0] statesInR_0_io_output_count; // @[NBuffers.scala 50:19:@40386.4]
  wire  statesInR_1_clock; // @[NBuffers.scala 50:19:@40397.4]
  wire  statesInR_1_reset; // @[NBuffers.scala 50:19:@40397.4]
  wire  statesInR_1_io_input_countUp; // @[NBuffers.scala 50:19:@40397.4]
  wire  statesInR_1_io_input_enable; // @[NBuffers.scala 50:19:@40397.4]
  wire [31:0] statesInR_1_io_output_count; // @[NBuffers.scala 50:19:@40397.4]
  wire  statesInR_2_clock; // @[NBuffers.scala 50:19:@40408.4]
  wire  statesInR_2_reset; // @[NBuffers.scala 50:19:@40408.4]
  wire  statesInR_2_io_input_countUp; // @[NBuffers.scala 50:19:@40408.4]
  wire  statesInR_2_io_input_enable; // @[NBuffers.scala 50:19:@40408.4]
  wire [31:0] statesInR_2_io_output_count; // @[NBuffers.scala 50:19:@40408.4]
  wire  statesInR_3_clock; // @[NBuffers.scala 50:19:@40419.4]
  wire  statesInR_3_reset; // @[NBuffers.scala 50:19:@40419.4]
  wire  statesInR_3_io_input_countUp; // @[NBuffers.scala 50:19:@40419.4]
  wire  statesInR_3_io_input_enable; // @[NBuffers.scala 50:19:@40419.4]
  wire [31:0] statesInR_3_io_output_count; // @[NBuffers.scala 50:19:@40419.4]
  wire  statesInR_4_clock; // @[NBuffers.scala 50:19:@40430.4]
  wire  statesInR_4_reset; // @[NBuffers.scala 50:19:@40430.4]
  wire  statesInR_4_io_input_countUp; // @[NBuffers.scala 50:19:@40430.4]
  wire  statesInR_4_io_input_enable; // @[NBuffers.scala 50:19:@40430.4]
  wire [31:0] statesInR_4_io_output_count; // @[NBuffers.scala 50:19:@40430.4]
  wire  statesInR_5_clock; // @[NBuffers.scala 50:19:@40441.4]
  wire  statesInR_5_reset; // @[NBuffers.scala 50:19:@40441.4]
  wire  statesInR_5_io_input_countUp; // @[NBuffers.scala 50:19:@40441.4]
  wire  statesInR_5_io_input_enable; // @[NBuffers.scala 50:19:@40441.4]
  wire [31:0] statesInR_5_io_output_count; // @[NBuffers.scala 50:19:@40441.4]
  wire  statesInR_6_clock; // @[NBuffers.scala 50:19:@40452.4]
  wire  statesInR_6_reset; // @[NBuffers.scala 50:19:@40452.4]
  wire  statesInR_6_io_input_countUp; // @[NBuffers.scala 50:19:@40452.4]
  wire  statesInR_6_io_input_enable; // @[NBuffers.scala 50:19:@40452.4]
  wire [31:0] statesInR_6_io_output_count; // @[NBuffers.scala 50:19:@40452.4]
  wire  _T_33; // @[NBuffers.scala 26:46:@40079.4]
  wire  _T_48; // @[NBuffers.scala 26:46:@40115.4]
  wire  _T_63; // @[NBuffers.scala 26:46:@40151.4]
  wire  _T_78; // @[NBuffers.scala 26:46:@40187.4]
  wire  _T_93; // @[NBuffers.scala 26:46:@40223.4]
  wire  _T_108; // @[NBuffers.scala 26:46:@40259.4]
  wire  _T_123; // @[NBuffers.scala 26:46:@40295.4]
  wire  _T_137; // @[NBuffers.scala 33:64:@40331.4]
  wire  _T_138; // @[NBuffers.scala 33:64:@40332.4]
  wire  _T_139; // @[NBuffers.scala 33:64:@40333.4]
  wire  _T_140; // @[NBuffers.scala 33:64:@40334.4]
  wire  _T_141; // @[NBuffers.scala 33:64:@40335.4]
  wire  anyEnabled; // @[NBuffers.scala 33:64:@40336.4]
  wire  _T_142; // @[NBuffers.scala 34:124:@40337.4]
  wire  _T_143; // @[NBuffers.scala 34:104:@40338.4]
  wire  _T_144; // @[NBuffers.scala 34:124:@40339.4]
  wire  _T_145; // @[NBuffers.scala 34:104:@40340.4]
  wire  _T_146; // @[NBuffers.scala 34:124:@40341.4]
  wire  _T_147; // @[NBuffers.scala 34:104:@40342.4]
  wire  _T_148; // @[NBuffers.scala 34:124:@40343.4]
  wire  _T_149; // @[NBuffers.scala 34:104:@40344.4]
  wire  _T_150; // @[NBuffers.scala 34:124:@40345.4]
  wire  _T_151; // @[NBuffers.scala 34:104:@40346.4]
  wire  _T_152; // @[NBuffers.scala 34:124:@40347.4]
  wire  _T_153; // @[NBuffers.scala 34:104:@40348.4]
  wire  _T_154; // @[NBuffers.scala 34:124:@40349.4]
  wire  _T_155; // @[NBuffers.scala 34:104:@40350.4]
  wire  _T_156; // @[NBuffers.scala 34:150:@40351.4]
  wire  _T_157; // @[NBuffers.scala 34:150:@40352.4]
  wire  _T_158; // @[NBuffers.scala 34:150:@40353.4]
  wire  _T_159; // @[NBuffers.scala 34:150:@40354.4]
  wire  _T_160; // @[NBuffers.scala 34:150:@40355.4]
  wire  _T_161; // @[NBuffers.scala 34:150:@40356.4]
  wire  _T_162; // @[NBuffers.scala 34:154:@40357.4]
  wire  _T_164; // @[package.scala 100:49:@40358.4]
  reg  _T_167; // @[package.scala 48:56:@40359.4]
  reg [31:0] _RAND_0;
  SRFF sEn_latch_0 ( // @[NBuffers.scala 21:52:@40036.4]
    .clock(sEn_latch_0_clock),
    .reset(sEn_latch_0_reset),
    .io_input_set(sEn_latch_0_io_input_set),
    .io_input_reset(sEn_latch_0_io_input_reset),
    .io_input_asyn_reset(sEn_latch_0_io_input_asyn_reset),
    .io_output(sEn_latch_0_io_output)
  );
  SRFF sEn_latch_1 ( // @[NBuffers.scala 21:52:@40039.4]
    .clock(sEn_latch_1_clock),
    .reset(sEn_latch_1_reset),
    .io_input_set(sEn_latch_1_io_input_set),
    .io_input_reset(sEn_latch_1_io_input_reset),
    .io_input_asyn_reset(sEn_latch_1_io_input_asyn_reset),
    .io_output(sEn_latch_1_io_output)
  );
  SRFF sEn_latch_2 ( // @[NBuffers.scala 21:52:@40042.4]
    .clock(sEn_latch_2_clock),
    .reset(sEn_latch_2_reset),
    .io_input_set(sEn_latch_2_io_input_set),
    .io_input_reset(sEn_latch_2_io_input_reset),
    .io_input_asyn_reset(sEn_latch_2_io_input_asyn_reset),
    .io_output(sEn_latch_2_io_output)
  );
  SRFF sEn_latch_3 ( // @[NBuffers.scala 21:52:@40045.4]
    .clock(sEn_latch_3_clock),
    .reset(sEn_latch_3_reset),
    .io_input_set(sEn_latch_3_io_input_set),
    .io_input_reset(sEn_latch_3_io_input_reset),
    .io_input_asyn_reset(sEn_latch_3_io_input_asyn_reset),
    .io_output(sEn_latch_3_io_output)
  );
  SRFF sEn_latch_4 ( // @[NBuffers.scala 21:52:@40048.4]
    .clock(sEn_latch_4_clock),
    .reset(sEn_latch_4_reset),
    .io_input_set(sEn_latch_4_io_input_set),
    .io_input_reset(sEn_latch_4_io_input_reset),
    .io_input_asyn_reset(sEn_latch_4_io_input_asyn_reset),
    .io_output(sEn_latch_4_io_output)
  );
  SRFF sEn_latch_5 ( // @[NBuffers.scala 21:52:@40051.4]
    .clock(sEn_latch_5_clock),
    .reset(sEn_latch_5_reset),
    .io_input_set(sEn_latch_5_io_input_set),
    .io_input_reset(sEn_latch_5_io_input_reset),
    .io_input_asyn_reset(sEn_latch_5_io_input_asyn_reset),
    .io_output(sEn_latch_5_io_output)
  );
  SRFF sEn_latch_6 ( // @[NBuffers.scala 21:52:@40054.4]
    .clock(sEn_latch_6_clock),
    .reset(sEn_latch_6_reset),
    .io_input_set(sEn_latch_6_io_input_set),
    .io_input_reset(sEn_latch_6_io_input_reset),
    .io_input_asyn_reset(sEn_latch_6_io_input_asyn_reset),
    .io_output(sEn_latch_6_io_output)
  );
  SRFF sDone_latch_0 ( // @[NBuffers.scala 22:54:@40057.4]
    .clock(sDone_latch_0_clock),
    .reset(sDone_latch_0_reset),
    .io_input_set(sDone_latch_0_io_input_set),
    .io_input_reset(sDone_latch_0_io_input_reset),
    .io_input_asyn_reset(sDone_latch_0_io_input_asyn_reset),
    .io_output(sDone_latch_0_io_output)
  );
  SRFF sDone_latch_1 ( // @[NBuffers.scala 22:54:@40060.4]
    .clock(sDone_latch_1_clock),
    .reset(sDone_latch_1_reset),
    .io_input_set(sDone_latch_1_io_input_set),
    .io_input_reset(sDone_latch_1_io_input_reset),
    .io_input_asyn_reset(sDone_latch_1_io_input_asyn_reset),
    .io_output(sDone_latch_1_io_output)
  );
  SRFF sDone_latch_2 ( // @[NBuffers.scala 22:54:@40063.4]
    .clock(sDone_latch_2_clock),
    .reset(sDone_latch_2_reset),
    .io_input_set(sDone_latch_2_io_input_set),
    .io_input_reset(sDone_latch_2_io_input_reset),
    .io_input_asyn_reset(sDone_latch_2_io_input_asyn_reset),
    .io_output(sDone_latch_2_io_output)
  );
  SRFF sDone_latch_3 ( // @[NBuffers.scala 22:54:@40066.4]
    .clock(sDone_latch_3_clock),
    .reset(sDone_latch_3_reset),
    .io_input_set(sDone_latch_3_io_input_set),
    .io_input_reset(sDone_latch_3_io_input_reset),
    .io_input_asyn_reset(sDone_latch_3_io_input_asyn_reset),
    .io_output(sDone_latch_3_io_output)
  );
  SRFF sDone_latch_4 ( // @[NBuffers.scala 22:54:@40069.4]
    .clock(sDone_latch_4_clock),
    .reset(sDone_latch_4_reset),
    .io_input_set(sDone_latch_4_io_input_set),
    .io_input_reset(sDone_latch_4_io_input_reset),
    .io_input_asyn_reset(sDone_latch_4_io_input_asyn_reset),
    .io_output(sDone_latch_4_io_output)
  );
  SRFF sDone_latch_5 ( // @[NBuffers.scala 22:54:@40072.4]
    .clock(sDone_latch_5_clock),
    .reset(sDone_latch_5_reset),
    .io_input_set(sDone_latch_5_io_input_set),
    .io_input_reset(sDone_latch_5_io_input_reset),
    .io_input_asyn_reset(sDone_latch_5_io_input_asyn_reset),
    .io_output(sDone_latch_5_io_output)
  );
  SRFF sDone_latch_6 ( // @[NBuffers.scala 22:54:@40075.4]
    .clock(sDone_latch_6_clock),
    .reset(sDone_latch_6_reset),
    .io_input_set(sDone_latch_6_io_input_set),
    .io_input_reset(sDone_latch_6_io_input_reset),
    .io_input_asyn_reset(sDone_latch_6_io_input_asyn_reset),
    .io_output(sDone_latch_6_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@40082.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@40090.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@40099.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@40107.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@40118.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@40126.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@40135.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@40143.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@40154.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@40162.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@40171.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 ( // @[package.scala 93:22:@40179.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper RetimeWrapper_12 ( // @[package.scala 93:22:@40190.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 ( // @[package.scala 93:22:@40198.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@40207.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@40215.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 ( // @[package.scala 93:22:@40226.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper RetimeWrapper_17 ( // @[package.scala 93:22:@40234.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 ( // @[package.scala 93:22:@40243.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper RetimeWrapper_19 ( // @[package.scala 93:22:@40251.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper RetimeWrapper_20 ( // @[package.scala 93:22:@40262.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper RetimeWrapper_21 ( // @[package.scala 93:22:@40270.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper RetimeWrapper_22 ( // @[package.scala 93:22:@40279.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper RetimeWrapper_23 ( // @[package.scala 93:22:@40287.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper RetimeWrapper_24 ( // @[package.scala 93:22:@40298.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@40306.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper RetimeWrapper_26 ( // @[package.scala 93:22:@40315.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper RetimeWrapper_27 ( // @[package.scala 93:22:@40323.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  NBufCtr_9 NBufCtr ( // @[NBuffers.scala 40:19:@40364.4]
    .clock(NBufCtr_clock),
    .reset(NBufCtr_reset),
    .io_input_countUp(NBufCtr_io_input_countUp),
    .io_input_enable(NBufCtr_io_input_enable),
    .io_output_count(NBufCtr_io_output_count)
  );
  NBufCtr_15 NBufCtr_1 ( // @[NBuffers.scala 40:19:@40375.4]
    .clock(NBufCtr_1_clock),
    .reset(NBufCtr_1_reset),
    .io_input_countUp(NBufCtr_1_io_input_countUp),
    .io_input_enable(NBufCtr_1_io_input_enable),
    .io_output_count(NBufCtr_1_io_output_count)
  );
  NBufCtr_9 statesInR_0 ( // @[NBuffers.scala 50:19:@40386.4]
    .clock(statesInR_0_clock),
    .reset(statesInR_0_reset),
    .io_input_countUp(statesInR_0_io_input_countUp),
    .io_input_enable(statesInR_0_io_input_enable),
    .io_output_count(statesInR_0_io_output_count)
  );
  NBufCtr_11 statesInR_1 ( // @[NBuffers.scala 50:19:@40397.4]
    .clock(statesInR_1_clock),
    .reset(statesInR_1_reset),
    .io_input_countUp(statesInR_1_io_input_countUp),
    .io_input_enable(statesInR_1_io_input_enable),
    .io_output_count(statesInR_1_io_output_count)
  );
  NBufCtr_12 statesInR_2 ( // @[NBuffers.scala 50:19:@40408.4]
    .clock(statesInR_2_clock),
    .reset(statesInR_2_reset),
    .io_input_countUp(statesInR_2_io_input_countUp),
    .io_input_enable(statesInR_2_io_input_enable),
    .io_output_count(statesInR_2_io_output_count)
  );
  NBufCtr_13 statesInR_3 ( // @[NBuffers.scala 50:19:@40419.4]
    .clock(statesInR_3_clock),
    .reset(statesInR_3_reset),
    .io_input_countUp(statesInR_3_io_input_countUp),
    .io_input_enable(statesInR_3_io_input_enable),
    .io_output_count(statesInR_3_io_output_count)
  );
  NBufCtr_14 statesInR_4 ( // @[NBuffers.scala 50:19:@40430.4]
    .clock(statesInR_4_clock),
    .reset(statesInR_4_reset),
    .io_input_countUp(statesInR_4_io_input_countUp),
    .io_input_enable(statesInR_4_io_input_enable),
    .io_output_count(statesInR_4_io_output_count)
  );
  NBufCtr_15 statesInR_5 ( // @[NBuffers.scala 50:19:@40441.4]
    .clock(statesInR_5_clock),
    .reset(statesInR_5_reset),
    .io_input_countUp(statesInR_5_io_input_countUp),
    .io_input_enable(statesInR_5_io_input_enable),
    .io_output_count(statesInR_5_io_output_count)
  );
  NBufCtr_16 statesInR_6 ( // @[NBuffers.scala 50:19:@40452.4]
    .clock(statesInR_6_clock),
    .reset(statesInR_6_reset),
    .io_input_countUp(statesInR_6_io_input_countUp),
    .io_input_enable(statesInR_6_io_input_enable),
    .io_output_count(statesInR_6_io_output_count)
  );
  assign _T_33 = io_sDone_0 == 1'h0; // @[NBuffers.scala 26:46:@40079.4]
  assign _T_48 = io_sDone_1 == 1'h0; // @[NBuffers.scala 26:46:@40115.4]
  assign _T_63 = io_sDone_2 == 1'h0; // @[NBuffers.scala 26:46:@40151.4]
  assign _T_78 = io_sDone_3 == 1'h0; // @[NBuffers.scala 26:46:@40187.4]
  assign _T_93 = io_sDone_4 == 1'h0; // @[NBuffers.scala 26:46:@40223.4]
  assign _T_108 = io_sDone_5 == 1'h0; // @[NBuffers.scala 26:46:@40259.4]
  assign _T_123 = io_sDone_6 == 1'h0; // @[NBuffers.scala 26:46:@40295.4]
  assign _T_137 = sEn_latch_0_io_output | sEn_latch_1_io_output; // @[NBuffers.scala 33:64:@40331.4]
  assign _T_138 = _T_137 | sEn_latch_2_io_output; // @[NBuffers.scala 33:64:@40332.4]
  assign _T_139 = _T_138 | sEn_latch_3_io_output; // @[NBuffers.scala 33:64:@40333.4]
  assign _T_140 = _T_139 | sEn_latch_4_io_output; // @[NBuffers.scala 33:64:@40334.4]
  assign _T_141 = _T_140 | sEn_latch_5_io_output; // @[NBuffers.scala 33:64:@40335.4]
  assign anyEnabled = _T_141 | sEn_latch_6_io_output; // @[NBuffers.scala 33:64:@40336.4]
  assign _T_142 = sDone_latch_0_io_output | io_sDone_0; // @[NBuffers.scala 34:124:@40337.4]
  assign _T_143 = sEn_latch_0_io_output == _T_142; // @[NBuffers.scala 34:104:@40338.4]
  assign _T_144 = sDone_latch_1_io_output | io_sDone_1; // @[NBuffers.scala 34:124:@40339.4]
  assign _T_145 = sEn_latch_1_io_output == _T_144; // @[NBuffers.scala 34:104:@40340.4]
  assign _T_146 = sDone_latch_2_io_output | io_sDone_2; // @[NBuffers.scala 34:124:@40341.4]
  assign _T_147 = sEn_latch_2_io_output == _T_146; // @[NBuffers.scala 34:104:@40342.4]
  assign _T_148 = sDone_latch_3_io_output | io_sDone_3; // @[NBuffers.scala 34:124:@40343.4]
  assign _T_149 = sEn_latch_3_io_output == _T_148; // @[NBuffers.scala 34:104:@40344.4]
  assign _T_150 = sDone_latch_4_io_output | io_sDone_4; // @[NBuffers.scala 34:124:@40345.4]
  assign _T_151 = sEn_latch_4_io_output == _T_150; // @[NBuffers.scala 34:104:@40346.4]
  assign _T_152 = sDone_latch_5_io_output | io_sDone_5; // @[NBuffers.scala 34:124:@40347.4]
  assign _T_153 = sEn_latch_5_io_output == _T_152; // @[NBuffers.scala 34:104:@40348.4]
  assign _T_154 = sDone_latch_6_io_output | io_sDone_6; // @[NBuffers.scala 34:124:@40349.4]
  assign _T_155 = sEn_latch_6_io_output == _T_154; // @[NBuffers.scala 34:104:@40350.4]
  assign _T_156 = _T_143 & _T_145; // @[NBuffers.scala 34:150:@40351.4]
  assign _T_157 = _T_156 & _T_147; // @[NBuffers.scala 34:150:@40352.4]
  assign _T_158 = _T_157 & _T_149; // @[NBuffers.scala 34:150:@40353.4]
  assign _T_159 = _T_158 & _T_151; // @[NBuffers.scala 34:150:@40354.4]
  assign _T_160 = _T_159 & _T_153; // @[NBuffers.scala 34:150:@40355.4]
  assign _T_161 = _T_160 & _T_155; // @[NBuffers.scala 34:150:@40356.4]
  assign _T_162 = _T_161 & anyEnabled; // @[NBuffers.scala 34:154:@40357.4]
  assign _T_164 = _T_162 == 1'h0; // @[package.scala 100:49:@40358.4]
  assign io_statesInW_0 = NBufCtr_io_output_count[3:0]; // @[NBuffers.scala 44:21:@40374.4]
  assign io_statesInW_1 = NBufCtr_1_io_output_count[3:0]; // @[NBuffers.scala 44:21:@40385.4]
  assign io_statesInR_6 = statesInR_6_io_output_count[3:0]; // @[NBuffers.scala 54:21:@40462.4]
  assign sEn_latch_0_clock = clock; // @[:@40037.4]
  assign sEn_latch_0_reset = reset; // @[:@40038.4]
  assign sEn_latch_0_io_input_set = io_sEn_0 & _T_33; // @[NBuffers.scala 26:31:@40081.4]
  assign sEn_latch_0_io_input_reset = RetimeWrapper_io_out; // @[NBuffers.scala 27:33:@40089.4]
  assign sEn_latch_0_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[NBuffers.scala 28:38:@40097.4]
  assign sEn_latch_1_clock = clock; // @[:@40040.4]
  assign sEn_latch_1_reset = reset; // @[:@40041.4]
  assign sEn_latch_1_io_input_set = io_sEn_1 & _T_48; // @[NBuffers.scala 26:31:@40117.4]
  assign sEn_latch_1_io_input_reset = RetimeWrapper_4_io_out; // @[NBuffers.scala 27:33:@40125.4]
  assign sEn_latch_1_io_input_asyn_reset = RetimeWrapper_5_io_out; // @[NBuffers.scala 28:38:@40133.4]
  assign sEn_latch_2_clock = clock; // @[:@40043.4]
  assign sEn_latch_2_reset = reset; // @[:@40044.4]
  assign sEn_latch_2_io_input_set = io_sEn_2 & _T_63; // @[NBuffers.scala 26:31:@40153.4]
  assign sEn_latch_2_io_input_reset = RetimeWrapper_8_io_out; // @[NBuffers.scala 27:33:@40161.4]
  assign sEn_latch_2_io_input_asyn_reset = RetimeWrapper_9_io_out; // @[NBuffers.scala 28:38:@40169.4]
  assign sEn_latch_3_clock = clock; // @[:@40046.4]
  assign sEn_latch_3_reset = reset; // @[:@40047.4]
  assign sEn_latch_3_io_input_set = io_sEn_3 & _T_78; // @[NBuffers.scala 26:31:@40189.4]
  assign sEn_latch_3_io_input_reset = RetimeWrapper_12_io_out; // @[NBuffers.scala 27:33:@40197.4]
  assign sEn_latch_3_io_input_asyn_reset = RetimeWrapper_13_io_out; // @[NBuffers.scala 28:38:@40205.4]
  assign sEn_latch_4_clock = clock; // @[:@40049.4]
  assign sEn_latch_4_reset = reset; // @[:@40050.4]
  assign sEn_latch_4_io_input_set = io_sEn_4 & _T_93; // @[NBuffers.scala 26:31:@40225.4]
  assign sEn_latch_4_io_input_reset = RetimeWrapper_16_io_out; // @[NBuffers.scala 27:33:@40233.4]
  assign sEn_latch_4_io_input_asyn_reset = RetimeWrapper_17_io_out; // @[NBuffers.scala 28:38:@40241.4]
  assign sEn_latch_5_clock = clock; // @[:@40052.4]
  assign sEn_latch_5_reset = reset; // @[:@40053.4]
  assign sEn_latch_5_io_input_set = io_sEn_5 & _T_108; // @[NBuffers.scala 26:31:@40261.4]
  assign sEn_latch_5_io_input_reset = RetimeWrapper_20_io_out; // @[NBuffers.scala 27:33:@40269.4]
  assign sEn_latch_5_io_input_asyn_reset = RetimeWrapper_21_io_out; // @[NBuffers.scala 28:38:@40277.4]
  assign sEn_latch_6_clock = clock; // @[:@40055.4]
  assign sEn_latch_6_reset = reset; // @[:@40056.4]
  assign sEn_latch_6_io_input_set = io_sEn_6 & _T_123; // @[NBuffers.scala 26:31:@40297.4]
  assign sEn_latch_6_io_input_reset = RetimeWrapper_24_io_out; // @[NBuffers.scala 27:33:@40305.4]
  assign sEn_latch_6_io_input_asyn_reset = RetimeWrapper_25_io_out; // @[NBuffers.scala 28:38:@40313.4]
  assign sDone_latch_0_clock = clock; // @[:@40058.4]
  assign sDone_latch_0_reset = reset; // @[:@40059.4]
  assign sDone_latch_0_io_input_set = io_sDone_0; // @[NBuffers.scala 29:33:@40098.4]
  assign sDone_latch_0_io_input_reset = RetimeWrapper_2_io_out; // @[NBuffers.scala 30:35:@40106.4]
  assign sDone_latch_0_io_input_asyn_reset = RetimeWrapper_3_io_out; // @[NBuffers.scala 31:40:@40114.4]
  assign sDone_latch_1_clock = clock; // @[:@40061.4]
  assign sDone_latch_1_reset = reset; // @[:@40062.4]
  assign sDone_latch_1_io_input_set = io_sDone_1; // @[NBuffers.scala 29:33:@40134.4]
  assign sDone_latch_1_io_input_reset = RetimeWrapper_6_io_out; // @[NBuffers.scala 30:35:@40142.4]
  assign sDone_latch_1_io_input_asyn_reset = RetimeWrapper_7_io_out; // @[NBuffers.scala 31:40:@40150.4]
  assign sDone_latch_2_clock = clock; // @[:@40064.4]
  assign sDone_latch_2_reset = reset; // @[:@40065.4]
  assign sDone_latch_2_io_input_set = io_sDone_2; // @[NBuffers.scala 29:33:@40170.4]
  assign sDone_latch_2_io_input_reset = RetimeWrapper_10_io_out; // @[NBuffers.scala 30:35:@40178.4]
  assign sDone_latch_2_io_input_asyn_reset = RetimeWrapper_11_io_out; // @[NBuffers.scala 31:40:@40186.4]
  assign sDone_latch_3_clock = clock; // @[:@40067.4]
  assign sDone_latch_3_reset = reset; // @[:@40068.4]
  assign sDone_latch_3_io_input_set = io_sDone_3; // @[NBuffers.scala 29:33:@40206.4]
  assign sDone_latch_3_io_input_reset = RetimeWrapper_14_io_out; // @[NBuffers.scala 30:35:@40214.4]
  assign sDone_latch_3_io_input_asyn_reset = RetimeWrapper_15_io_out; // @[NBuffers.scala 31:40:@40222.4]
  assign sDone_latch_4_clock = clock; // @[:@40070.4]
  assign sDone_latch_4_reset = reset; // @[:@40071.4]
  assign sDone_latch_4_io_input_set = io_sDone_4; // @[NBuffers.scala 29:33:@40242.4]
  assign sDone_latch_4_io_input_reset = RetimeWrapper_18_io_out; // @[NBuffers.scala 30:35:@40250.4]
  assign sDone_latch_4_io_input_asyn_reset = RetimeWrapper_19_io_out; // @[NBuffers.scala 31:40:@40258.4]
  assign sDone_latch_5_clock = clock; // @[:@40073.4]
  assign sDone_latch_5_reset = reset; // @[:@40074.4]
  assign sDone_latch_5_io_input_set = io_sDone_5; // @[NBuffers.scala 29:33:@40278.4]
  assign sDone_latch_5_io_input_reset = RetimeWrapper_22_io_out; // @[NBuffers.scala 30:35:@40286.4]
  assign sDone_latch_5_io_input_asyn_reset = RetimeWrapper_23_io_out; // @[NBuffers.scala 31:40:@40294.4]
  assign sDone_latch_6_clock = clock; // @[:@40076.4]
  assign sDone_latch_6_reset = reset; // @[:@40077.4]
  assign sDone_latch_6_io_input_set = io_sDone_6; // @[NBuffers.scala 29:33:@40314.4]
  assign sDone_latch_6_io_input_reset = RetimeWrapper_26_io_out; // @[NBuffers.scala 30:35:@40322.4]
  assign sDone_latch_6_io_input_asyn_reset = RetimeWrapper_27_io_out; // @[NBuffers.scala 31:40:@40330.4]
  assign RetimeWrapper_clock = clock; // @[:@40083.4]
  assign RetimeWrapper_reset = reset; // @[:@40084.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@40086.4]
  assign RetimeWrapper_io_in = _T_162 & _T_167; // @[package.scala 94:16:@40085.4]
  assign RetimeWrapper_1_clock = clock; // @[:@40091.4]
  assign RetimeWrapper_1_reset = reset; // @[:@40092.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@40094.4]
  assign RetimeWrapper_1_io_in = reset; // @[package.scala 94:16:@40093.4]
  assign RetimeWrapper_2_clock = clock; // @[:@40100.4]
  assign RetimeWrapper_2_reset = reset; // @[:@40101.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@40103.4]
  assign RetimeWrapper_2_io_in = _T_162 & _T_167; // @[package.scala 94:16:@40102.4]
  assign RetimeWrapper_3_clock = clock; // @[:@40108.4]
  assign RetimeWrapper_3_reset = reset; // @[:@40109.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@40111.4]
  assign RetimeWrapper_3_io_in = reset; // @[package.scala 94:16:@40110.4]
  assign RetimeWrapper_4_clock = clock; // @[:@40119.4]
  assign RetimeWrapper_4_reset = reset; // @[:@40120.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@40122.4]
  assign RetimeWrapper_4_io_in = _T_162 & _T_167; // @[package.scala 94:16:@40121.4]
  assign RetimeWrapper_5_clock = clock; // @[:@40127.4]
  assign RetimeWrapper_5_reset = reset; // @[:@40128.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@40130.4]
  assign RetimeWrapper_5_io_in = reset; // @[package.scala 94:16:@40129.4]
  assign RetimeWrapper_6_clock = clock; // @[:@40136.4]
  assign RetimeWrapper_6_reset = reset; // @[:@40137.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@40139.4]
  assign RetimeWrapper_6_io_in = _T_162 & _T_167; // @[package.scala 94:16:@40138.4]
  assign RetimeWrapper_7_clock = clock; // @[:@40144.4]
  assign RetimeWrapper_7_reset = reset; // @[:@40145.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@40147.4]
  assign RetimeWrapper_7_io_in = reset; // @[package.scala 94:16:@40146.4]
  assign RetimeWrapper_8_clock = clock; // @[:@40155.4]
  assign RetimeWrapper_8_reset = reset; // @[:@40156.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@40158.4]
  assign RetimeWrapper_8_io_in = _T_162 & _T_167; // @[package.scala 94:16:@40157.4]
  assign RetimeWrapper_9_clock = clock; // @[:@40163.4]
  assign RetimeWrapper_9_reset = reset; // @[:@40164.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@40166.4]
  assign RetimeWrapper_9_io_in = reset; // @[package.scala 94:16:@40165.4]
  assign RetimeWrapper_10_clock = clock; // @[:@40172.4]
  assign RetimeWrapper_10_reset = reset; // @[:@40173.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@40175.4]
  assign RetimeWrapper_10_io_in = _T_162 & _T_167; // @[package.scala 94:16:@40174.4]
  assign RetimeWrapper_11_clock = clock; // @[:@40180.4]
  assign RetimeWrapper_11_reset = reset; // @[:@40181.4]
  assign RetimeWrapper_11_io_flow = 1'h1; // @[package.scala 95:18:@40183.4]
  assign RetimeWrapper_11_io_in = reset; // @[package.scala 94:16:@40182.4]
  assign RetimeWrapper_12_clock = clock; // @[:@40191.4]
  assign RetimeWrapper_12_reset = reset; // @[:@40192.4]
  assign RetimeWrapper_12_io_flow = 1'h1; // @[package.scala 95:18:@40194.4]
  assign RetimeWrapper_12_io_in = _T_162 & _T_167; // @[package.scala 94:16:@40193.4]
  assign RetimeWrapper_13_clock = clock; // @[:@40199.4]
  assign RetimeWrapper_13_reset = reset; // @[:@40200.4]
  assign RetimeWrapper_13_io_flow = 1'h1; // @[package.scala 95:18:@40202.4]
  assign RetimeWrapper_13_io_in = reset; // @[package.scala 94:16:@40201.4]
  assign RetimeWrapper_14_clock = clock; // @[:@40208.4]
  assign RetimeWrapper_14_reset = reset; // @[:@40209.4]
  assign RetimeWrapper_14_io_flow = 1'h1; // @[package.scala 95:18:@40211.4]
  assign RetimeWrapper_14_io_in = _T_162 & _T_167; // @[package.scala 94:16:@40210.4]
  assign RetimeWrapper_15_clock = clock; // @[:@40216.4]
  assign RetimeWrapper_15_reset = reset; // @[:@40217.4]
  assign RetimeWrapper_15_io_flow = 1'h1; // @[package.scala 95:18:@40219.4]
  assign RetimeWrapper_15_io_in = reset; // @[package.scala 94:16:@40218.4]
  assign RetimeWrapper_16_clock = clock; // @[:@40227.4]
  assign RetimeWrapper_16_reset = reset; // @[:@40228.4]
  assign RetimeWrapper_16_io_flow = 1'h1; // @[package.scala 95:18:@40230.4]
  assign RetimeWrapper_16_io_in = _T_162 & _T_167; // @[package.scala 94:16:@40229.4]
  assign RetimeWrapper_17_clock = clock; // @[:@40235.4]
  assign RetimeWrapper_17_reset = reset; // @[:@40236.4]
  assign RetimeWrapper_17_io_flow = 1'h1; // @[package.scala 95:18:@40238.4]
  assign RetimeWrapper_17_io_in = reset; // @[package.scala 94:16:@40237.4]
  assign RetimeWrapper_18_clock = clock; // @[:@40244.4]
  assign RetimeWrapper_18_reset = reset; // @[:@40245.4]
  assign RetimeWrapper_18_io_flow = 1'h1; // @[package.scala 95:18:@40247.4]
  assign RetimeWrapper_18_io_in = _T_162 & _T_167; // @[package.scala 94:16:@40246.4]
  assign RetimeWrapper_19_clock = clock; // @[:@40252.4]
  assign RetimeWrapper_19_reset = reset; // @[:@40253.4]
  assign RetimeWrapper_19_io_flow = 1'h1; // @[package.scala 95:18:@40255.4]
  assign RetimeWrapper_19_io_in = reset; // @[package.scala 94:16:@40254.4]
  assign RetimeWrapper_20_clock = clock; // @[:@40263.4]
  assign RetimeWrapper_20_reset = reset; // @[:@40264.4]
  assign RetimeWrapper_20_io_flow = 1'h1; // @[package.scala 95:18:@40266.4]
  assign RetimeWrapper_20_io_in = _T_162 & _T_167; // @[package.scala 94:16:@40265.4]
  assign RetimeWrapper_21_clock = clock; // @[:@40271.4]
  assign RetimeWrapper_21_reset = reset; // @[:@40272.4]
  assign RetimeWrapper_21_io_flow = 1'h1; // @[package.scala 95:18:@40274.4]
  assign RetimeWrapper_21_io_in = reset; // @[package.scala 94:16:@40273.4]
  assign RetimeWrapper_22_clock = clock; // @[:@40280.4]
  assign RetimeWrapper_22_reset = reset; // @[:@40281.4]
  assign RetimeWrapper_22_io_flow = 1'h1; // @[package.scala 95:18:@40283.4]
  assign RetimeWrapper_22_io_in = _T_162 & _T_167; // @[package.scala 94:16:@40282.4]
  assign RetimeWrapper_23_clock = clock; // @[:@40288.4]
  assign RetimeWrapper_23_reset = reset; // @[:@40289.4]
  assign RetimeWrapper_23_io_flow = 1'h1; // @[package.scala 95:18:@40291.4]
  assign RetimeWrapper_23_io_in = reset; // @[package.scala 94:16:@40290.4]
  assign RetimeWrapper_24_clock = clock; // @[:@40299.4]
  assign RetimeWrapper_24_reset = reset; // @[:@40300.4]
  assign RetimeWrapper_24_io_flow = 1'h1; // @[package.scala 95:18:@40302.4]
  assign RetimeWrapper_24_io_in = _T_162 & _T_167; // @[package.scala 94:16:@40301.4]
  assign RetimeWrapper_25_clock = clock; // @[:@40307.4]
  assign RetimeWrapper_25_reset = reset; // @[:@40308.4]
  assign RetimeWrapper_25_io_flow = 1'h1; // @[package.scala 95:18:@40310.4]
  assign RetimeWrapper_25_io_in = reset; // @[package.scala 94:16:@40309.4]
  assign RetimeWrapper_26_clock = clock; // @[:@40316.4]
  assign RetimeWrapper_26_reset = reset; // @[:@40317.4]
  assign RetimeWrapper_26_io_flow = 1'h1; // @[package.scala 95:18:@40319.4]
  assign RetimeWrapper_26_io_in = _T_162 & _T_167; // @[package.scala 94:16:@40318.4]
  assign RetimeWrapper_27_clock = clock; // @[:@40324.4]
  assign RetimeWrapper_27_reset = reset; // @[:@40325.4]
  assign RetimeWrapper_27_io_flow = 1'h1; // @[package.scala 95:18:@40327.4]
  assign RetimeWrapper_27_io_in = reset; // @[package.scala 94:16:@40326.4]
  assign NBufCtr_clock = clock; // @[:@40365.4]
  assign NBufCtr_reset = reset; // @[:@40366.4]
  assign NBufCtr_io_input_countUp = 1'h0; // @[NBuffers.scala 43:24:@40373.4]
  assign NBufCtr_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 42:23:@40372.4]
  assign NBufCtr_1_clock = clock; // @[:@40376.4]
  assign NBufCtr_1_reset = reset; // @[:@40377.4]
  assign NBufCtr_1_io_input_countUp = 1'h0; // @[NBuffers.scala 43:24:@40384.4]
  assign NBufCtr_1_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 42:23:@40383.4]
  assign statesInR_0_clock = clock; // @[:@40387.4]
  assign statesInR_0_reset = reset; // @[:@40388.4]
  assign statesInR_0_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@40395.4]
  assign statesInR_0_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@40394.4]
  assign statesInR_1_clock = clock; // @[:@40398.4]
  assign statesInR_1_reset = reset; // @[:@40399.4]
  assign statesInR_1_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@40406.4]
  assign statesInR_1_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@40405.4]
  assign statesInR_2_clock = clock; // @[:@40409.4]
  assign statesInR_2_reset = reset; // @[:@40410.4]
  assign statesInR_2_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@40417.4]
  assign statesInR_2_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@40416.4]
  assign statesInR_3_clock = clock; // @[:@40420.4]
  assign statesInR_3_reset = reset; // @[:@40421.4]
  assign statesInR_3_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@40428.4]
  assign statesInR_3_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@40427.4]
  assign statesInR_4_clock = clock; // @[:@40431.4]
  assign statesInR_4_reset = reset; // @[:@40432.4]
  assign statesInR_4_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@40439.4]
  assign statesInR_4_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@40438.4]
  assign statesInR_5_clock = clock; // @[:@40442.4]
  assign statesInR_5_reset = reset; // @[:@40443.4]
  assign statesInR_5_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@40450.4]
  assign statesInR_5_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@40449.4]
  assign statesInR_6_clock = clock; // @[:@40453.4]
  assign statesInR_6_reset = reset; // @[:@40454.4]
  assign statesInR_6_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@40461.4]
  assign statesInR_6_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@40460.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_167 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_167 <= 1'h0;
    end else begin
      _T_167 <= _T_164;
    end
  end
endmodule
module x558_tmp_4( // @[:@41983.2]
  input         clock, // @[:@41984.4]
  input         reset, // @[:@41985.4]
  input  [1:0]  io_rPort_0_ofs_0, // @[:@41986.4]
  input         io_rPort_0_en_0, // @[:@41986.4]
  output [31:0] io_rPort_0_output_0, // @[:@41986.4]
  input  [1:0]  io_wPort_1_ofs_0, // @[:@41986.4]
  input  [31:0] io_wPort_1_data_0, // @[:@41986.4]
  input         io_wPort_1_en_0, // @[:@41986.4]
  input  [1:0]  io_wPort_0_ofs_0, // @[:@41986.4]
  input  [31:0] io_wPort_0_data_0, // @[:@41986.4]
  input         io_wPort_0_en_0, // @[:@41986.4]
  input         io_sEn_0, // @[:@41986.4]
  input         io_sEn_1, // @[:@41986.4]
  input         io_sEn_2, // @[:@41986.4]
  input         io_sEn_3, // @[:@41986.4]
  input         io_sEn_4, // @[:@41986.4]
  input         io_sEn_5, // @[:@41986.4]
  input         io_sEn_6, // @[:@41986.4]
  input         io_sDone_0, // @[:@41986.4]
  input         io_sDone_1, // @[:@41986.4]
  input         io_sDone_2, // @[:@41986.4]
  input         io_sDone_3, // @[:@41986.4]
  input         io_sDone_4, // @[:@41986.4]
  input         io_sDone_5, // @[:@41986.4]
  input         io_sDone_6 // @[:@41986.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@41996.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@41996.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@41996.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@41996.4]
  wire  ctrl_io_sEn_2; // @[NBuffers.scala 83:20:@41996.4]
  wire  ctrl_io_sEn_3; // @[NBuffers.scala 83:20:@41996.4]
  wire  ctrl_io_sEn_4; // @[NBuffers.scala 83:20:@41996.4]
  wire  ctrl_io_sEn_5; // @[NBuffers.scala 83:20:@41996.4]
  wire  ctrl_io_sEn_6; // @[NBuffers.scala 83:20:@41996.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@41996.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@41996.4]
  wire  ctrl_io_sDone_2; // @[NBuffers.scala 83:20:@41996.4]
  wire  ctrl_io_sDone_3; // @[NBuffers.scala 83:20:@41996.4]
  wire  ctrl_io_sDone_4; // @[NBuffers.scala 83:20:@41996.4]
  wire  ctrl_io_sDone_5; // @[NBuffers.scala 83:20:@41996.4]
  wire  ctrl_io_sDone_6; // @[NBuffers.scala 83:20:@41996.4]
  wire [3:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@41996.4]
  wire [3:0] ctrl_io_statesInW_1; // @[NBuffers.scala 83:20:@41996.4]
  wire [3:0] ctrl_io_statesInR_6; // @[NBuffers.scala 83:20:@41996.4]
  wire  SRAM_clock; // @[NBuffers.scala 94:23:@42013.4]
  wire  SRAM_reset; // @[NBuffers.scala 94:23:@42013.4]
  wire [1:0] SRAM_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@42013.4]
  wire  SRAM_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@42013.4]
  wire  SRAM_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@42013.4]
  wire [31:0] SRAM_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@42013.4]
  wire [1:0] SRAM_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@42013.4]
  wire [31:0] SRAM_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@42013.4]
  wire  SRAM_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@42013.4]
  wire [1:0] SRAM_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@42013.4]
  wire [31:0] SRAM_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@42013.4]
  wire  SRAM_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@42013.4]
  wire  SRAM_1_clock; // @[NBuffers.scala 94:23:@42036.4]
  wire  SRAM_1_reset; // @[NBuffers.scala 94:23:@42036.4]
  wire [1:0] SRAM_1_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@42036.4]
  wire  SRAM_1_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@42036.4]
  wire  SRAM_1_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@42036.4]
  wire [31:0] SRAM_1_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@42036.4]
  wire [1:0] SRAM_1_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@42036.4]
  wire [31:0] SRAM_1_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@42036.4]
  wire  SRAM_1_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@42036.4]
  wire [1:0] SRAM_1_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@42036.4]
  wire [31:0] SRAM_1_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@42036.4]
  wire  SRAM_1_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@42036.4]
  wire  SRAM_2_clock; // @[NBuffers.scala 94:23:@42059.4]
  wire  SRAM_2_reset; // @[NBuffers.scala 94:23:@42059.4]
  wire [1:0] SRAM_2_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@42059.4]
  wire  SRAM_2_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@42059.4]
  wire  SRAM_2_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@42059.4]
  wire [31:0] SRAM_2_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@42059.4]
  wire [1:0] SRAM_2_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@42059.4]
  wire [31:0] SRAM_2_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@42059.4]
  wire  SRAM_2_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@42059.4]
  wire [1:0] SRAM_2_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@42059.4]
  wire [31:0] SRAM_2_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@42059.4]
  wire  SRAM_2_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@42059.4]
  wire  SRAM_3_clock; // @[NBuffers.scala 94:23:@42082.4]
  wire  SRAM_3_reset; // @[NBuffers.scala 94:23:@42082.4]
  wire [1:0] SRAM_3_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@42082.4]
  wire  SRAM_3_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@42082.4]
  wire  SRAM_3_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@42082.4]
  wire [31:0] SRAM_3_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@42082.4]
  wire [1:0] SRAM_3_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@42082.4]
  wire [31:0] SRAM_3_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@42082.4]
  wire  SRAM_3_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@42082.4]
  wire [1:0] SRAM_3_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@42082.4]
  wire [31:0] SRAM_3_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@42082.4]
  wire  SRAM_3_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@42082.4]
  wire  SRAM_4_clock; // @[NBuffers.scala 94:23:@42105.4]
  wire  SRAM_4_reset; // @[NBuffers.scala 94:23:@42105.4]
  wire [1:0] SRAM_4_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@42105.4]
  wire  SRAM_4_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@42105.4]
  wire  SRAM_4_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@42105.4]
  wire [31:0] SRAM_4_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@42105.4]
  wire [1:0] SRAM_4_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@42105.4]
  wire [31:0] SRAM_4_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@42105.4]
  wire  SRAM_4_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@42105.4]
  wire [1:0] SRAM_4_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@42105.4]
  wire [31:0] SRAM_4_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@42105.4]
  wire  SRAM_4_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@42105.4]
  wire  SRAM_5_clock; // @[NBuffers.scala 94:23:@42128.4]
  wire  SRAM_5_reset; // @[NBuffers.scala 94:23:@42128.4]
  wire [1:0] SRAM_5_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@42128.4]
  wire  SRAM_5_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@42128.4]
  wire  SRAM_5_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@42128.4]
  wire [31:0] SRAM_5_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@42128.4]
  wire [1:0] SRAM_5_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@42128.4]
  wire [31:0] SRAM_5_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@42128.4]
  wire  SRAM_5_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@42128.4]
  wire [1:0] SRAM_5_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@42128.4]
  wire [31:0] SRAM_5_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@42128.4]
  wire  SRAM_5_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@42128.4]
  wire  SRAM_6_clock; // @[NBuffers.scala 94:23:@42151.4]
  wire  SRAM_6_reset; // @[NBuffers.scala 94:23:@42151.4]
  wire [1:0] SRAM_6_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@42151.4]
  wire  SRAM_6_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@42151.4]
  wire  SRAM_6_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@42151.4]
  wire [31:0] SRAM_6_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@42151.4]
  wire [1:0] SRAM_6_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@42151.4]
  wire [31:0] SRAM_6_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@42151.4]
  wire  SRAM_6_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@42151.4]
  wire [1:0] SRAM_6_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@42151.4]
  wire [31:0] SRAM_6_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@42151.4]
  wire  SRAM_6_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@42151.4]
  wire  _T_148; // @[NBuffers.scala 104:105:@42174.4]
  wire  _T_152; // @[NBuffers.scala 104:105:@42184.4]
  wire  _T_156; // @[NBuffers.scala 108:92:@42194.4]
  wire  _T_159; // @[NBuffers.scala 104:105:@42200.4]
  wire  _T_163; // @[NBuffers.scala 104:105:@42210.4]
  wire  _T_167; // @[NBuffers.scala 108:92:@42220.4]
  wire  _T_170; // @[NBuffers.scala 104:105:@42226.4]
  wire  _T_174; // @[NBuffers.scala 104:105:@42236.4]
  wire  _T_178; // @[NBuffers.scala 108:92:@42246.4]
  wire  _T_181; // @[NBuffers.scala 104:105:@42252.4]
  wire  _T_185; // @[NBuffers.scala 104:105:@42262.4]
  wire  _T_189; // @[NBuffers.scala 108:92:@42272.4]
  wire  _T_192; // @[NBuffers.scala 104:105:@42278.4]
  wire  _T_196; // @[NBuffers.scala 104:105:@42288.4]
  wire  _T_200; // @[NBuffers.scala 108:92:@42298.4]
  wire  _T_203; // @[NBuffers.scala 104:105:@42304.4]
  wire  _T_207; // @[NBuffers.scala 104:105:@42314.4]
  wire  _T_211; // @[NBuffers.scala 108:92:@42324.4]
  wire  _T_214; // @[NBuffers.scala 104:105:@42330.4]
  wire  _T_218; // @[NBuffers.scala 104:105:@42340.4]
  wire  _T_222; // @[NBuffers.scala 108:92:@42350.4]
  wire [31:0] _T_240; // @[Mux.scala 19:72:@42363.4]
  wire [31:0] _T_242; // @[Mux.scala 19:72:@42364.4]
  wire [31:0] _T_244; // @[Mux.scala 19:72:@42365.4]
  wire [31:0] _T_246; // @[Mux.scala 19:72:@42366.4]
  wire [31:0] _T_248; // @[Mux.scala 19:72:@42367.4]
  wire [31:0] _T_250; // @[Mux.scala 19:72:@42368.4]
  wire [31:0] _T_252; // @[Mux.scala 19:72:@42369.4]
  wire [31:0] _T_253; // @[Mux.scala 19:72:@42370.4]
  wire [31:0] _T_254; // @[Mux.scala 19:72:@42371.4]
  wire [31:0] _T_255; // @[Mux.scala 19:72:@42372.4]
  wire [31:0] _T_256; // @[Mux.scala 19:72:@42373.4]
  wire [31:0] _T_257; // @[Mux.scala 19:72:@42374.4]
  NBufController_9 ctrl ( // @[NBuffers.scala 83:20:@41996.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sEn_2(ctrl_io_sEn_2),
    .io_sEn_3(ctrl_io_sEn_3),
    .io_sEn_4(ctrl_io_sEn_4),
    .io_sEn_5(ctrl_io_sEn_5),
    .io_sEn_6(ctrl_io_sEn_6),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_sDone_2(ctrl_io_sDone_2),
    .io_sDone_3(ctrl_io_sDone_3),
    .io_sDone_4(ctrl_io_sDone_4),
    .io_sDone_5(ctrl_io_sDone_5),
    .io_sDone_6(ctrl_io_sDone_6),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInW_1(ctrl_io_statesInW_1),
    .io_statesInR_6(ctrl_io_statesInR_6)
  );
  SRAM_10 SRAM ( // @[NBuffers.scala 94:23:@42013.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_rPort_0_ofs_0(SRAM_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_1 ( // @[NBuffers.scala 94:23:@42036.4]
    .clock(SRAM_1_clock),
    .reset(SRAM_1_reset),
    .io_rPort_0_ofs_0(SRAM_1_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_1_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_1_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_1_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_1_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_1_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_1_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_1_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_1_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_2 ( // @[NBuffers.scala 94:23:@42059.4]
    .clock(SRAM_2_clock),
    .reset(SRAM_2_reset),
    .io_rPort_0_ofs_0(SRAM_2_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_2_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_2_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_2_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_2_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_2_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_2_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_2_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_2_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_2_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_3 ( // @[NBuffers.scala 94:23:@42082.4]
    .clock(SRAM_3_clock),
    .reset(SRAM_3_reset),
    .io_rPort_0_ofs_0(SRAM_3_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_3_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_3_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_3_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_3_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_3_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_3_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_3_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_3_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_3_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_4 ( // @[NBuffers.scala 94:23:@42105.4]
    .clock(SRAM_4_clock),
    .reset(SRAM_4_reset),
    .io_rPort_0_ofs_0(SRAM_4_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_4_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_4_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_4_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_4_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_4_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_4_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_4_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_4_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_4_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_5 ( // @[NBuffers.scala 94:23:@42128.4]
    .clock(SRAM_5_clock),
    .reset(SRAM_5_reset),
    .io_rPort_0_ofs_0(SRAM_5_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_5_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_5_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_5_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_5_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_5_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_5_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_5_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_5_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_5_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_6 ( // @[NBuffers.scala 94:23:@42151.4]
    .clock(SRAM_6_clock),
    .reset(SRAM_6_reset),
    .io_rPort_0_ofs_0(SRAM_6_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_6_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_6_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_6_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_6_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_6_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_6_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_6_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_6_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_6_io_wPort_0_en_0)
  );
  assign _T_148 = ctrl_io_statesInW_0 == 4'h0; // @[NBuffers.scala 104:105:@42174.4]
  assign _T_152 = ctrl_io_statesInW_1 == 4'h0; // @[NBuffers.scala 104:105:@42184.4]
  assign _T_156 = ctrl_io_statesInR_6 == 4'h0; // @[NBuffers.scala 108:92:@42194.4]
  assign _T_159 = ctrl_io_statesInW_0 == 4'h1; // @[NBuffers.scala 104:105:@42200.4]
  assign _T_163 = ctrl_io_statesInW_1 == 4'h1; // @[NBuffers.scala 104:105:@42210.4]
  assign _T_167 = ctrl_io_statesInR_6 == 4'h1; // @[NBuffers.scala 108:92:@42220.4]
  assign _T_170 = ctrl_io_statesInW_0 == 4'h2; // @[NBuffers.scala 104:105:@42226.4]
  assign _T_174 = ctrl_io_statesInW_1 == 4'h2; // @[NBuffers.scala 104:105:@42236.4]
  assign _T_178 = ctrl_io_statesInR_6 == 4'h2; // @[NBuffers.scala 108:92:@42246.4]
  assign _T_181 = ctrl_io_statesInW_0 == 4'h3; // @[NBuffers.scala 104:105:@42252.4]
  assign _T_185 = ctrl_io_statesInW_1 == 4'h3; // @[NBuffers.scala 104:105:@42262.4]
  assign _T_189 = ctrl_io_statesInR_6 == 4'h3; // @[NBuffers.scala 108:92:@42272.4]
  assign _T_192 = ctrl_io_statesInW_0 == 4'h4; // @[NBuffers.scala 104:105:@42278.4]
  assign _T_196 = ctrl_io_statesInW_1 == 4'h4; // @[NBuffers.scala 104:105:@42288.4]
  assign _T_200 = ctrl_io_statesInR_6 == 4'h4; // @[NBuffers.scala 108:92:@42298.4]
  assign _T_203 = ctrl_io_statesInW_0 == 4'h5; // @[NBuffers.scala 104:105:@42304.4]
  assign _T_207 = ctrl_io_statesInW_1 == 4'h5; // @[NBuffers.scala 104:105:@42314.4]
  assign _T_211 = ctrl_io_statesInR_6 == 4'h5; // @[NBuffers.scala 108:92:@42324.4]
  assign _T_214 = ctrl_io_statesInW_0 == 4'h6; // @[NBuffers.scala 104:105:@42330.4]
  assign _T_218 = ctrl_io_statesInW_1 == 4'h6; // @[NBuffers.scala 104:105:@42340.4]
  assign _T_222 = ctrl_io_statesInR_6 == 4'h6; // @[NBuffers.scala 108:92:@42350.4]
  assign _T_240 = _T_156 ? SRAM_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@42363.4]
  assign _T_242 = _T_167 ? SRAM_1_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@42364.4]
  assign _T_244 = _T_178 ? SRAM_2_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@42365.4]
  assign _T_246 = _T_189 ? SRAM_3_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@42366.4]
  assign _T_248 = _T_200 ? SRAM_4_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@42367.4]
  assign _T_250 = _T_211 ? SRAM_5_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@42368.4]
  assign _T_252 = _T_222 ? SRAM_6_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@42369.4]
  assign _T_253 = _T_240 | _T_242; // @[Mux.scala 19:72:@42370.4]
  assign _T_254 = _T_253 | _T_244; // @[Mux.scala 19:72:@42371.4]
  assign _T_255 = _T_254 | _T_246; // @[Mux.scala 19:72:@42372.4]
  assign _T_256 = _T_255 | _T_248; // @[Mux.scala 19:72:@42373.4]
  assign _T_257 = _T_256 | _T_250; // @[Mux.scala 19:72:@42374.4]
  assign io_rPort_0_output_0 = _T_257 | _T_252; // @[NBuffers.scala 115:66:@42378.4]
  assign ctrl_clock = clock; // @[:@41997.4]
  assign ctrl_reset = reset; // @[:@41998.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@41999.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@42001.4]
  assign ctrl_io_sEn_2 = io_sEn_2; // @[NBuffers.scala 85:20:@42003.4]
  assign ctrl_io_sEn_3 = io_sEn_3; // @[NBuffers.scala 85:20:@42005.4]
  assign ctrl_io_sEn_4 = io_sEn_4; // @[NBuffers.scala 85:20:@42007.4]
  assign ctrl_io_sEn_5 = io_sEn_5; // @[NBuffers.scala 85:20:@42009.4]
  assign ctrl_io_sEn_6 = io_sEn_6; // @[NBuffers.scala 85:20:@42011.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@42000.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@42002.4]
  assign ctrl_io_sDone_2 = io_sDone_2; // @[NBuffers.scala 86:22:@42004.4]
  assign ctrl_io_sDone_3 = io_sDone_3; // @[NBuffers.scala 86:22:@42006.4]
  assign ctrl_io_sDone_4 = io_sDone_4; // @[NBuffers.scala 86:22:@42008.4]
  assign ctrl_io_sDone_5 = io_sDone_5; // @[NBuffers.scala 86:22:@42010.4]
  assign ctrl_io_sDone_6 = io_sDone_6; // @[NBuffers.scala 86:22:@42012.4]
  assign SRAM_clock = clock; // @[:@42014.4]
  assign SRAM_reset = reset; // @[:@42015.4]
  assign SRAM_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@42196.4]
  assign SRAM_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_156; // @[MemPrimitives.scala 43:33:@42198.4]
  assign SRAM_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@42199.4]
  assign SRAM_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@42186.4]
  assign SRAM_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@42187.4]
  assign SRAM_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_152; // @[MemPrimitives.scala 37:29:@42193.4]
  assign SRAM_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@42176.4]
  assign SRAM_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@42177.4]
  assign SRAM_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_148; // @[MemPrimitives.scala 37:29:@42183.4]
  assign SRAM_1_clock = clock; // @[:@42037.4]
  assign SRAM_1_reset = reset; // @[:@42038.4]
  assign SRAM_1_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@42222.4]
  assign SRAM_1_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_167; // @[MemPrimitives.scala 43:33:@42224.4]
  assign SRAM_1_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@42225.4]
  assign SRAM_1_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@42212.4]
  assign SRAM_1_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@42213.4]
  assign SRAM_1_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_163; // @[MemPrimitives.scala 37:29:@42219.4]
  assign SRAM_1_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@42202.4]
  assign SRAM_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@42203.4]
  assign SRAM_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_159; // @[MemPrimitives.scala 37:29:@42209.4]
  assign SRAM_2_clock = clock; // @[:@42060.4]
  assign SRAM_2_reset = reset; // @[:@42061.4]
  assign SRAM_2_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@42248.4]
  assign SRAM_2_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_178; // @[MemPrimitives.scala 43:33:@42250.4]
  assign SRAM_2_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@42251.4]
  assign SRAM_2_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@42238.4]
  assign SRAM_2_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@42239.4]
  assign SRAM_2_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_174; // @[MemPrimitives.scala 37:29:@42245.4]
  assign SRAM_2_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@42228.4]
  assign SRAM_2_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@42229.4]
  assign SRAM_2_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_170; // @[MemPrimitives.scala 37:29:@42235.4]
  assign SRAM_3_clock = clock; // @[:@42083.4]
  assign SRAM_3_reset = reset; // @[:@42084.4]
  assign SRAM_3_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@42274.4]
  assign SRAM_3_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_189; // @[MemPrimitives.scala 43:33:@42276.4]
  assign SRAM_3_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@42277.4]
  assign SRAM_3_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@42264.4]
  assign SRAM_3_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@42265.4]
  assign SRAM_3_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_185; // @[MemPrimitives.scala 37:29:@42271.4]
  assign SRAM_3_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@42254.4]
  assign SRAM_3_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@42255.4]
  assign SRAM_3_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_181; // @[MemPrimitives.scala 37:29:@42261.4]
  assign SRAM_4_clock = clock; // @[:@42106.4]
  assign SRAM_4_reset = reset; // @[:@42107.4]
  assign SRAM_4_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@42300.4]
  assign SRAM_4_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_200; // @[MemPrimitives.scala 43:33:@42302.4]
  assign SRAM_4_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@42303.4]
  assign SRAM_4_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@42290.4]
  assign SRAM_4_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@42291.4]
  assign SRAM_4_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_196; // @[MemPrimitives.scala 37:29:@42297.4]
  assign SRAM_4_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@42280.4]
  assign SRAM_4_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@42281.4]
  assign SRAM_4_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_192; // @[MemPrimitives.scala 37:29:@42287.4]
  assign SRAM_5_clock = clock; // @[:@42129.4]
  assign SRAM_5_reset = reset; // @[:@42130.4]
  assign SRAM_5_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@42326.4]
  assign SRAM_5_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_211; // @[MemPrimitives.scala 43:33:@42328.4]
  assign SRAM_5_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@42329.4]
  assign SRAM_5_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@42316.4]
  assign SRAM_5_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@42317.4]
  assign SRAM_5_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_207; // @[MemPrimitives.scala 37:29:@42323.4]
  assign SRAM_5_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@42306.4]
  assign SRAM_5_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@42307.4]
  assign SRAM_5_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_203; // @[MemPrimitives.scala 37:29:@42313.4]
  assign SRAM_6_clock = clock; // @[:@42152.4]
  assign SRAM_6_reset = reset; // @[:@42153.4]
  assign SRAM_6_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@42352.4]
  assign SRAM_6_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_222; // @[MemPrimitives.scala 43:33:@42354.4]
  assign SRAM_6_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@42355.4]
  assign SRAM_6_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@42342.4]
  assign SRAM_6_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@42343.4]
  assign SRAM_6_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_218; // @[MemPrimitives.scala 37:29:@42349.4]
  assign SRAM_6_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@42332.4]
  assign SRAM_6_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@42333.4]
  assign SRAM_6_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_214; // @[MemPrimitives.scala 37:29:@42339.4]
endmodule
module RetimeWrapper_452( // @[:@42581.2]
  input   clock, // @[:@42582.4]
  input   reset, // @[:@42583.4]
  input   io_flow, // @[:@42584.4]
  input   io_in, // @[:@42584.4]
  output  io_out // @[:@42584.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@42586.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@42586.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@42586.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@42586.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@42586.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@42586.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@42586.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@42599.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@42598.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@42597.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@42596.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@42595.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@42593.4]
endmodule
module x579_inr_Foreach_sm( // @[:@42729.2]
  input   clock, // @[:@42730.4]
  input   reset, // @[:@42731.4]
  input   io_enable, // @[:@42732.4]
  output  io_done, // @[:@42732.4]
  input   io_ctrDone, // @[:@42732.4]
  output  io_datapathEn, // @[:@42732.4]
  output  io_ctrInc, // @[:@42732.4]
  output  io_ctrRst, // @[:@42732.4]
  input   io_parentAck, // @[:@42732.4]
  input   io_backpressure, // @[:@42732.4]
  input   io_break // @[:@42732.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@42734.4]
  wire  active_reset; // @[Controllers.scala 261:22:@42734.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@42734.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@42734.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@42734.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@42734.4]
  wire  done_clock; // @[Controllers.scala 262:20:@42737.4]
  wire  done_reset; // @[Controllers.scala 262:20:@42737.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@42737.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@42737.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@42737.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@42737.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@42771.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@42771.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@42771.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@42771.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@42771.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@42793.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@42793.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@42793.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@42793.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@42793.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@42805.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@42805.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@42805.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@42805.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@42805.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@42813.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@42813.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@42813.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@42813.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@42813.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@42829.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@42829.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@42829.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@42829.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@42829.4]
  wire  _T_80; // @[Controllers.scala 264:48:@42742.4]
  wire  _T_81; // @[Controllers.scala 264:46:@42743.4]
  wire  _T_82; // @[Controllers.scala 264:62:@42744.4]
  wire  _T_100; // @[package.scala 100:49:@42762.4]
  reg  _T_103; // @[package.scala 48:56:@42763.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@42776.4 package.scala 96:25:@42777.4]
  wire  _T_110; // @[package.scala 100:49:@42778.4]
  reg  _T_113; // @[package.scala 48:56:@42779.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@42781.4]
  wire  _T_118; // @[Controllers.scala 283:41:@42786.4]
  wire  _T_124; // @[package.scala 96:25:@42798.4 package.scala 96:25:@42799.4]
  wire  _T_126; // @[package.scala 100:49:@42800.4]
  reg  _T_129; // @[package.scala 48:56:@42801.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@42825.4]
  reg  _T_153; // @[package.scala 48:56:@42826.4]
  reg [31:0] _RAND_3;
  SRFF active ( // @[Controllers.scala 261:22:@42734.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@42737.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_452 RetimeWrapper ( // @[package.scala 93:22:@42771.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_452 RetimeWrapper_1 ( // @[package.scala 93:22:@42793.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@42805.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@42813.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_4 ( // @[package.scala 93:22:@42829.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@42742.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@42743.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@42744.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@42762.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@42776.4 package.scala 96:25:@42777.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@42778.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@42781.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@42786.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@42798.4 package.scala 96:25:@42799.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@42800.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@42825.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@42804.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@42789.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@42792.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@42784.4]
  assign active_clock = clock; // @[:@42735.4]
  assign active_reset = reset; // @[:@42736.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@42747.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@42751.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@42752.4]
  assign done_clock = clock; // @[:@42738.4]
  assign done_reset = reset; // @[:@42739.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@42767.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@42760.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@42761.4]
  assign RetimeWrapper_clock = clock; // @[:@42772.4]
  assign RetimeWrapper_reset = reset; // @[:@42773.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@42775.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@42774.4]
  assign RetimeWrapper_1_clock = clock; // @[:@42794.4]
  assign RetimeWrapper_1_reset = reset; // @[:@42795.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@42797.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@42796.4]
  assign RetimeWrapper_2_clock = clock; // @[:@42806.4]
  assign RetimeWrapper_2_reset = reset; // @[:@42807.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@42809.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@42808.4]
  assign RetimeWrapper_3_clock = clock; // @[:@42814.4]
  assign RetimeWrapper_3_reset = reset; // @[:@42815.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@42817.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@42816.4]
  assign RetimeWrapper_4_clock = clock; // @[:@42830.4]
  assign RetimeWrapper_4_reset = reset; // @[:@42831.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@42833.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@42832.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox_38( // @[:@44087.2]
  input  [31:0] io_a, // @[:@44090.4]
  output [32:0] io_b // @[:@44090.4]
);
  wire [21:0] tmp_frac; // @[SimBlackBoxes.scala 56:25:@44098.4]
  wire  _T_19; // @[implicits.scala 70:16:@44100.4]
  wire [9:0] _T_20; // @[SimBlackBoxes.scala 88:77:@44102.4]
  wire [10:0] new_dec; // @[Cat.scala 30:58:@44103.4]
  assign tmp_frac = io_a[21:0]; // @[SimBlackBoxes.scala 56:25:@44098.4]
  assign _T_19 = io_a[31]; // @[implicits.scala 70:16:@44100.4]
  assign _T_20 = io_a[31:22]; // @[SimBlackBoxes.scala 88:77:@44102.4]
  assign new_dec = {_T_19,_T_20}; // @[Cat.scala 30:58:@44103.4]
  assign io_b = {new_dec,tmp_frac}; // @[SimBlackBoxes.scala 98:40:@44106.4]
endmodule
module __37( // @[:@44108.2]
  input  [31:0] io_b, // @[:@44111.4]
  output [32:0] io_result // @[:@44111.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@44116.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@44116.4]
  SimBlackBoxesfix2fixBox_38 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@44116.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 717:17:@44129.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@44124.4]
endmodule
module fix2fixBox_12( // @[:@44207.2]
  input         clock, // @[:@44208.4]
  input         reset, // @[:@44209.4]
  input  [32:0] io_a, // @[:@44210.4]
  input         io_flow, // @[:@44210.4]
  output [31:0] io_b // @[:@44210.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@44224.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@44224.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@44224.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@44224.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@44224.4]
  wire [21:0] tmp_frac; // @[Converter.scala 52:23:@44218.4]
  wire [9:0] new_dec; // @[Converter.scala 63:26:@44221.4]
  RetimeWrapper_32 RetimeWrapper ( // @[package.scala 93:22:@44224.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign tmp_frac = io_a[21:0]; // @[Converter.scala 52:23:@44218.4]
  assign new_dec = io_a[31:22]; // @[Converter.scala 63:26:@44221.4]
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 94:38:@44231.4]
  assign RetimeWrapper_clock = clock; // @[:@44225.4]
  assign RetimeWrapper_reset = reset; // @[:@44226.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@44228.4]
  assign RetimeWrapper_io_in = {new_dec,tmp_frac}; // @[package.scala 94:16:@44227.4]
endmodule
module x573_sub( // @[:@44233.2]
  input         clock, // @[:@44234.4]
  input         reset, // @[:@44235.4]
  input  [31:0] io_a, // @[:@44236.4]
  input  [31:0] io_b, // @[:@44236.4]
  output [31:0] io_result // @[:@44236.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@44244.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@44244.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@44251.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@44251.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@44270.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@44270.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@44270.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@44270.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@44270.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@44249.4 Math.scala 724:14:@44250.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@44256.4 Math.scala 724:14:@44257.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@44258.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@44259.4]
  __37 _ ( // @[Math.scala 720:24:@44244.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __37 __1 ( // @[Math.scala 720:24:@44251.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_12 fix2fixBox ( // @[Math.scala 182:30:@44270.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@44249.4 Math.scala 724:14:@44250.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@44256.4 Math.scala 724:14:@44257.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@44258.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@44259.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@44278.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@44247.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@44254.4]
  assign fix2fixBox_clock = clock; // @[:@44271.4]
  assign fix2fixBox_reset = reset; // @[:@44272.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@44273.4]
  assign fix2fixBox_io_flow = 1'h1; // @[Math.scala 186:26:@44276.4]
endmodule
module RetimeWrapper_475( // @[:@44292.2]
  input         clock, // @[:@44293.4]
  input         reset, // @[:@44294.4]
  input  [31:0] io_in, // @[:@44295.4]
  output [31:0] io_out // @[:@44295.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@44297.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@44297.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@44297.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@44297.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@44297.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@44297.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@44297.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@44310.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@44309.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@44308.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@44307.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@44306.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@44304.4]
endmodule
module x579_inr_Foreach_kernelx579_inr_Foreach_concrete1( // @[:@44728.2]
  input         clock, // @[:@44729.4]
  input         reset, // @[:@44730.4]
  output [1:0]  io_in_x555_tmp_1_wPort_0_ofs_0, // @[:@44731.4]
  output [31:0] io_in_x555_tmp_1_wPort_0_data_0, // @[:@44731.4]
  output        io_in_x555_tmp_1_wPort_0_en_0, // @[:@44731.4]
  output        io_in_x555_tmp_1_sEn_0, // @[:@44731.4]
  output        io_in_x555_tmp_1_sDone_0, // @[:@44731.4]
  input  [31:0] io_in_b550_number, // @[:@44731.4]
  output [8:0]  io_in_x472_A_sram_1_rPort_0_ofs_0, // @[:@44731.4]
  output        io_in_x472_A_sram_1_rPort_0_en_0, // @[:@44731.4]
  input  [31:0] io_in_x472_A_sram_1_rPort_0_output_0, // @[:@44731.4]
  input  [31:0] io_in_b542_number, // @[:@44731.4]
  output [8:0]  io_in_x471_A_sram_0_rPort_0_ofs_0, // @[:@44731.4]
  output        io_in_x471_A_sram_0_rPort_0_en_0, // @[:@44731.4]
  input  [31:0] io_in_x471_A_sram_0_rPort_0_output_0, // @[:@44731.4]
  output [1:0]  io_in_x554_tmp_0_wPort_0_ofs_0, // @[:@44731.4]
  output [31:0] io_in_x554_tmp_0_wPort_0_data_0, // @[:@44731.4]
  output        io_in_x554_tmp_0_wPort_0_en_0, // @[:@44731.4]
  output        io_in_x554_tmp_0_sEn_0, // @[:@44731.4]
  output        io_in_x554_tmp_0_sDone_0, // @[:@44731.4]
  output [1:0]  io_in_x558_tmp_4_wPort_0_ofs_0, // @[:@44731.4]
  output [31:0] io_in_x558_tmp_4_wPort_0_data_0, // @[:@44731.4]
  output        io_in_x558_tmp_4_wPort_0_en_0, // @[:@44731.4]
  output        io_in_x558_tmp_4_sEn_0, // @[:@44731.4]
  output        io_in_x558_tmp_4_sDone_0, // @[:@44731.4]
  input         io_in_b552, // @[:@44731.4]
  output [1:0]  io_in_x557_tmp_3_wPort_0_ofs_0, // @[:@44731.4]
  output [31:0] io_in_x557_tmp_3_wPort_0_data_0, // @[:@44731.4]
  output        io_in_x557_tmp_3_wPort_0_en_0, // @[:@44731.4]
  output        io_in_x557_tmp_3_sEn_0, // @[:@44731.4]
  output        io_in_x557_tmp_3_sDone_0, // @[:@44731.4]
  output [1:0]  io_in_x556_tmp_2_wPort_0_ofs_0, // @[:@44731.4]
  output [31:0] io_in_x556_tmp_2_wPort_0_data_0, // @[:@44731.4]
  output        io_in_x556_tmp_2_wPort_0_en_0, // @[:@44731.4]
  output        io_in_x556_tmp_2_sEn_0, // @[:@44731.4]
  output        io_in_x556_tmp_2_sDone_0, // @[:@44731.4]
  input         io_in_b543, // @[:@44731.4]
  output [63:0] io_in_instrctrs_8_cycs, // @[:@44731.4]
  output [63:0] io_in_instrctrs_8_iters, // @[:@44731.4]
  input         io_sigsIn_done, // @[:@44731.4]
  input         io_sigsIn_datapathEn, // @[:@44731.4]
  input         io_sigsIn_baseEn, // @[:@44731.4]
  input         io_sigsIn_break, // @[:@44731.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@44731.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@44731.4]
  input         io_rr // @[:@44731.4]
);
  wire  cycles_x579_inr_Foreach_clock; // @[sm_x579_inr_Foreach.scala 101:43:@45080.4]
  wire  cycles_x579_inr_Foreach_reset; // @[sm_x579_inr_Foreach.scala 101:43:@45080.4]
  wire  cycles_x579_inr_Foreach_io_enable; // @[sm_x579_inr_Foreach.scala 101:43:@45080.4]
  wire [63:0] cycles_x579_inr_Foreach_io_count; // @[sm_x579_inr_Foreach.scala 101:43:@45080.4]
  wire  iters_x579_inr_Foreach_clock; // @[sm_x579_inr_Foreach.scala 102:42:@45083.4]
  wire  iters_x579_inr_Foreach_reset; // @[sm_x579_inr_Foreach.scala 102:42:@45083.4]
  wire  iters_x579_inr_Foreach_io_enable; // @[sm_x579_inr_Foreach.scala 102:42:@45083.4]
  wire [63:0] iters_x579_inr_Foreach_io_count; // @[sm_x579_inr_Foreach.scala 102:42:@45083.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@45100.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@45100.4]
  wire  x745_sum_1_clock; // @[Math.scala 150:24:@45115.4]
  wire  x745_sum_1_reset; // @[Math.scala 150:24:@45115.4]
  wire [31:0] x745_sum_1_io_a; // @[Math.scala 150:24:@45115.4]
  wire [31:0] x745_sum_1_io_b; // @[Math.scala 150:24:@45115.4]
  wire  x745_sum_1_io_flow; // @[Math.scala 150:24:@45115.4]
  wire [31:0] x745_sum_1_io_result; // @[Math.scala 150:24:@45115.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@45126.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@45126.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@45126.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@45126.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@45126.4]
  wire  x565_sum_1_clock; // @[Math.scala 150:24:@45135.4]
  wire  x565_sum_1_reset; // @[Math.scala 150:24:@45135.4]
  wire [31:0] x565_sum_1_io_a; // @[Math.scala 150:24:@45135.4]
  wire [31:0] x565_sum_1_io_b; // @[Math.scala 150:24:@45135.4]
  wire  x565_sum_1_io_flow; // @[Math.scala 150:24:@45135.4]
  wire [31:0] x565_sum_1_io_result; // @[Math.scala 150:24:@45135.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@45146.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@45146.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@45146.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@45146.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@45146.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@45156.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@45156.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@45156.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@45156.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@45156.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@45166.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@45166.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@45166.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@45166.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@45166.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@45178.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@45178.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@45178.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@45178.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@45178.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@45190.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@45190.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@45190.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@45190.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@45190.4]
  wire  x747_sum_1_clock; // @[Math.scala 150:24:@45216.4]
  wire  x747_sum_1_reset; // @[Math.scala 150:24:@45216.4]
  wire [31:0] x747_sum_1_io_a; // @[Math.scala 150:24:@45216.4]
  wire [31:0] x747_sum_1_io_b; // @[Math.scala 150:24:@45216.4]
  wire  x747_sum_1_io_flow; // @[Math.scala 150:24:@45216.4]
  wire [31:0] x747_sum_1_io_result; // @[Math.scala 150:24:@45216.4]
  wire  x570_sum_1_clock; // @[Math.scala 150:24:@45226.4]
  wire  x570_sum_1_reset; // @[Math.scala 150:24:@45226.4]
  wire [31:0] x570_sum_1_io_a; // @[Math.scala 150:24:@45226.4]
  wire [31:0] x570_sum_1_io_b; // @[Math.scala 150:24:@45226.4]
  wire  x570_sum_1_io_flow; // @[Math.scala 150:24:@45226.4]
  wire [31:0] x570_sum_1_io_result; // @[Math.scala 150:24:@45226.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@45239.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@45239.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@45239.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@45239.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@45239.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@45251.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@45251.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@45251.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@45251.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@45251.4]
  wire  x573_sub_1_clock; // @[Math.scala 191:24:@45272.4]
  wire  x573_sub_1_reset; // @[Math.scala 191:24:@45272.4]
  wire [31:0] x573_sub_1_io_a; // @[Math.scala 191:24:@45272.4]
  wire [31:0] x573_sub_1_io_b; // @[Math.scala 191:24:@45272.4]
  wire [31:0] x573_sub_1_io_result; // @[Math.scala 191:24:@45272.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@45283.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@45283.4]
  wire [31:0] RetimeWrapper_8_io_in; // @[package.scala 93:22:@45283.4]
  wire [31:0] RetimeWrapper_8_io_out; // @[package.scala 93:22:@45283.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@45293.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@45293.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@45293.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@45293.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@45293.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@45303.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@45303.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@45303.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@45303.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@45303.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@45313.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@45313.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@45313.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@45313.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@45313.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@45327.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@45327.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@45327.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@45327.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@45327.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@45353.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@45353.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@45353.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@45353.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@45353.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@45379.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@45379.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@45379.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@45379.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@45379.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@45405.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@45405.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@45405.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@45405.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@45405.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@45431.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@45431.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@45431.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@45431.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@45431.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@45452.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@45452.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@45452.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@45452.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@45452.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@45463.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@45463.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@45463.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@45463.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@45463.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@45474.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@45474.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@45474.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@45474.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@45474.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@45485.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@45485.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@45485.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@45485.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@45485.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@45496.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@45496.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@45496.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@45496.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@45496.4]
  wire  _T_1814; // @[package.scala 100:49:@45087.4]
  reg  _T_1817; // @[package.scala 48:56:@45088.4]
  reg [31:0] _RAND_0;
  wire [32:0] _GEN_0; // @[Math.scala 461:32:@45111.4]
  wire [32:0] _T_1831; // @[Math.scala 461:32:@45111.4]
  wire  _T_1873; // @[package.scala 96:25:@45183.4 package.scala 96:25:@45184.4]
  wire  _T_1875; // @[implicits.scala 56:10:@45185.4]
  wire  _T_1876; // @[sm_x579_inr_Foreach.scala 126:114:@45186.4]
  wire  _T_1877; // @[sm_x579_inr_Foreach.scala 126:111:@45187.4]
  wire  _T_1882; // @[package.scala 96:25:@45195.4 package.scala 96:25:@45196.4]
  wire  _T_1884; // @[implicits.scala 56:10:@45197.4]
  wire  _T_1885; // @[sm_x579_inr_Foreach.scala 126:131:@45198.4]
  wire  x772_b562_D2; // @[package.scala 96:25:@45171.4 package.scala 96:25:@45172.4]
  wire  _T_1886; // @[sm_x579_inr_Foreach.scala 126:228:@45199.4]
  wire  x771_b552_D2; // @[package.scala 96:25:@45161.4 package.scala 96:25:@45162.4]
  wire  _T_1887; // @[sm_x579_inr_Foreach.scala 126:236:@45200.4]
  wire  x770_b543_D2; // @[package.scala 96:25:@45151.4 package.scala 96:25:@45152.4]
  wire [32:0] _GEN_1; // @[Math.scala 461:32:@45212.4]
  wire [32:0] _T_1893; // @[Math.scala 461:32:@45212.4]
  wire  _T_1915; // @[package.scala 96:25:@45244.4 package.scala 96:25:@45245.4]
  wire  _T_1917; // @[implicits.scala 56:10:@45246.4]
  wire  _T_1919; // @[sm_x579_inr_Foreach.scala 141:111:@45248.4]
  wire  _T_1924; // @[package.scala 96:25:@45256.4 package.scala 96:25:@45257.4]
  wire  _T_1926; // @[implicits.scala 56:10:@45258.4]
  wire  _T_1927; // @[sm_x579_inr_Foreach.scala 141:131:@45259.4]
  wire  _T_1928; // @[sm_x579_inr_Foreach.scala 141:228:@45260.4]
  wire  _T_1929; // @[sm_x579_inr_Foreach.scala 141:236:@45261.4]
  wire  _T_1966; // @[package.scala 96:25:@45332.4 package.scala 96:25:@45333.4]
  wire  _T_1968; // @[implicits.scala 56:10:@45334.4]
  wire  _T_1969; // @[sm_x579_inr_Foreach.scala 160:115:@45335.4]
  wire  _T_1971; // @[sm_x579_inr_Foreach.scala 160:212:@45337.4]
  wire  x774_b562_D5; // @[package.scala 96:25:@45298.4 package.scala 96:25:@45299.4]
  wire  _T_1973; // @[sm_x579_inr_Foreach.scala 160:257:@45339.4]
  wire  x775_b552_D5; // @[package.scala 96:25:@45308.4 package.scala 96:25:@45309.4]
  wire  _T_1974; // @[sm_x579_inr_Foreach.scala 160:265:@45340.4]
  wire  x776_b543_D5; // @[package.scala 96:25:@45318.4 package.scala 96:25:@45319.4]
  wire  _T_1986; // @[package.scala 96:25:@45358.4 package.scala 96:25:@45359.4]
  wire  _T_1988; // @[implicits.scala 56:10:@45360.4]
  wire  _T_1989; // @[sm_x579_inr_Foreach.scala 165:115:@45361.4]
  wire  _T_1991; // @[sm_x579_inr_Foreach.scala 165:212:@45363.4]
  wire  _T_1993; // @[sm_x579_inr_Foreach.scala 165:257:@45365.4]
  wire  _T_1994; // @[sm_x579_inr_Foreach.scala 165:265:@45366.4]
  wire  _T_2006; // @[package.scala 96:25:@45384.4 package.scala 96:25:@45385.4]
  wire  _T_2008; // @[implicits.scala 56:10:@45386.4]
  wire  _T_2009; // @[sm_x579_inr_Foreach.scala 170:115:@45387.4]
  wire  _T_2011; // @[sm_x579_inr_Foreach.scala 170:212:@45389.4]
  wire  _T_2013; // @[sm_x579_inr_Foreach.scala 170:257:@45391.4]
  wire  _T_2014; // @[sm_x579_inr_Foreach.scala 170:265:@45392.4]
  wire  _T_2026; // @[package.scala 96:25:@45410.4 package.scala 96:25:@45411.4]
  wire  _T_2028; // @[implicits.scala 56:10:@45412.4]
  wire  _T_2029; // @[sm_x579_inr_Foreach.scala 175:115:@45413.4]
  wire  _T_2031; // @[sm_x579_inr_Foreach.scala 175:212:@45415.4]
  wire  _T_2033; // @[sm_x579_inr_Foreach.scala 175:257:@45417.4]
  wire  _T_2034; // @[sm_x579_inr_Foreach.scala 175:265:@45418.4]
  wire  _T_2046; // @[package.scala 96:25:@45436.4 package.scala 96:25:@45437.4]
  wire  _T_2048; // @[implicits.scala 56:10:@45438.4]
  wire  _T_2049; // @[sm_x579_inr_Foreach.scala 180:115:@45439.4]
  wire  _T_2051; // @[sm_x579_inr_Foreach.scala 180:212:@45441.4]
  wire  _T_2053; // @[sm_x579_inr_Foreach.scala 180:257:@45443.4]
  wire  _T_2054; // @[sm_x579_inr_Foreach.scala 180:265:@45444.4]
  wire  _T_2059; // @[package.scala 96:25:@45457.4 package.scala 96:25:@45458.4]
  wire  _T_2065; // @[package.scala 96:25:@45468.4 package.scala 96:25:@45469.4]
  wire  _T_2071; // @[package.scala 96:25:@45479.4 package.scala 96:25:@45480.4]
  wire  _T_2077; // @[package.scala 96:25:@45490.4 package.scala 96:25:@45491.4]
  wire  _T_2083; // @[package.scala 96:25:@45501.4 package.scala 96:25:@45502.4]
  wire [31:0] x565_sum_number; // @[Math.scala 154:22:@45141.4 Math.scala 155:14:@45142.4]
  wire [31:0] x570_sum_number; // @[Math.scala 154:22:@45232.4 Math.scala 155:14:@45233.4]
  wire [31:0] x773_b561_D5_number; // @[package.scala 96:25:@45288.4 package.scala 96:25:@45289.4]
  InstrumentationCounter cycles_x579_inr_Foreach ( // @[sm_x579_inr_Foreach.scala 101:43:@45080.4]
    .clock(cycles_x579_inr_Foreach_clock),
    .reset(cycles_x579_inr_Foreach_reset),
    .io_enable(cycles_x579_inr_Foreach_io_enable),
    .io_count(cycles_x579_inr_Foreach_io_count)
  );
  InstrumentationCounter iters_x579_inr_Foreach ( // @[sm_x579_inr_Foreach.scala 102:42:@45083.4]
    .clock(iters_x579_inr_Foreach_clock),
    .reset(iters_x579_inr_Foreach_reset),
    .io_enable(iters_x579_inr_Foreach_io_enable),
    .io_count(iters_x579_inr_Foreach_io_count)
  );
  _ _ ( // @[Math.scala 720:24:@45100.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x739_sum x745_sum_1 ( // @[Math.scala 150:24:@45115.4]
    .clock(x745_sum_1_clock),
    .reset(x745_sum_1_reset),
    .io_a(x745_sum_1_io_a),
    .io_b(x745_sum_1_io_b),
    .io_flow(x745_sum_1_io_flow),
    .io_result(x745_sum_1_io_result)
  );
  RetimeWrapper_32 RetimeWrapper ( // @[package.scala 93:22:@45126.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x739_sum x565_sum_1 ( // @[Math.scala 150:24:@45135.4]
    .clock(x565_sum_1_clock),
    .reset(x565_sum_1_reset),
    .io_a(x565_sum_1_io_a),
    .io_b(x565_sum_1_io_b),
    .io_flow(x565_sum_1_io_flow),
    .io_result(x565_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@45146.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@45156.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@45166.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@45178.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@45190.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  x739_sum x747_sum_1 ( // @[Math.scala 150:24:@45216.4]
    .clock(x747_sum_1_clock),
    .reset(x747_sum_1_reset),
    .io_a(x747_sum_1_io_a),
    .io_b(x747_sum_1_io_b),
    .io_flow(x747_sum_1_io_flow),
    .io_result(x747_sum_1_io_result)
  );
  x739_sum x570_sum_1 ( // @[Math.scala 150:24:@45226.4]
    .clock(x570_sum_1_clock),
    .reset(x570_sum_1_reset),
    .io_a(x570_sum_1_io_a),
    .io_b(x570_sum_1_io_b),
    .io_flow(x570_sum_1_io_flow),
    .io_result(x570_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@45239.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@45251.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  x573_sub x573_sub_1 ( // @[Math.scala 191:24:@45272.4]
    .clock(x573_sub_1_clock),
    .reset(x573_sub_1_reset),
    .io_a(x573_sub_1_io_a),
    .io_b(x573_sub_1_io_b),
    .io_result(x573_sub_1_io_result)
  );
  RetimeWrapper_475 RetimeWrapper_8 ( // @[package.scala 93:22:@45283.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_9 ( // @[package.scala 93:22:@45293.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_10 ( // @[package.scala 93:22:@45303.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_11 ( // @[package.scala 93:22:@45313.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_12 ( // @[package.scala 93:22:@45327.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_13 ( // @[package.scala 93:22:@45353.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_14 ( // @[package.scala 93:22:@45379.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_15 ( // @[package.scala 93:22:@45405.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_16 ( // @[package.scala 93:22:@45431.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper RetimeWrapper_17 ( // @[package.scala 93:22:@45452.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 ( // @[package.scala 93:22:@45463.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper RetimeWrapper_19 ( // @[package.scala 93:22:@45474.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper RetimeWrapper_20 ( // @[package.scala 93:22:@45485.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper RetimeWrapper_21 ( // @[package.scala 93:22:@45496.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  assign _T_1814 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@45087.4]
  assign _GEN_0 = {{1'd0}, io_in_b542_number}; // @[Math.scala 461:32:@45111.4]
  assign _T_1831 = _GEN_0 << 1; // @[Math.scala 461:32:@45111.4]
  assign _T_1873 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@45183.4 package.scala 96:25:@45184.4]
  assign _T_1875 = io_rr ? _T_1873 : 1'h0; // @[implicits.scala 56:10:@45185.4]
  assign _T_1876 = ~ io_sigsIn_break; // @[sm_x579_inr_Foreach.scala 126:114:@45186.4]
  assign _T_1877 = _T_1875 & _T_1876; // @[sm_x579_inr_Foreach.scala 126:111:@45187.4]
  assign _T_1882 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@45195.4 package.scala 96:25:@45196.4]
  assign _T_1884 = io_rr ? _T_1882 : 1'h0; // @[implicits.scala 56:10:@45197.4]
  assign _T_1885 = _T_1877 & _T_1884; // @[sm_x579_inr_Foreach.scala 126:131:@45198.4]
  assign x772_b562_D2 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@45171.4 package.scala 96:25:@45172.4]
  assign _T_1886 = _T_1885 & x772_b562_D2; // @[sm_x579_inr_Foreach.scala 126:228:@45199.4]
  assign x771_b552_D2 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@45161.4 package.scala 96:25:@45162.4]
  assign _T_1887 = _T_1886 & x771_b552_D2; // @[sm_x579_inr_Foreach.scala 126:236:@45200.4]
  assign x770_b543_D2 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@45151.4 package.scala 96:25:@45152.4]
  assign _GEN_1 = {{1'd0}, io_in_b550_number}; // @[Math.scala 461:32:@45212.4]
  assign _T_1893 = _GEN_1 << 1; // @[Math.scala 461:32:@45212.4]
  assign _T_1915 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@45244.4 package.scala 96:25:@45245.4]
  assign _T_1917 = io_rr ? _T_1915 : 1'h0; // @[implicits.scala 56:10:@45246.4]
  assign _T_1919 = _T_1917 & _T_1876; // @[sm_x579_inr_Foreach.scala 141:111:@45248.4]
  assign _T_1924 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@45256.4 package.scala 96:25:@45257.4]
  assign _T_1926 = io_rr ? _T_1924 : 1'h0; // @[implicits.scala 56:10:@45258.4]
  assign _T_1927 = _T_1919 & _T_1926; // @[sm_x579_inr_Foreach.scala 141:131:@45259.4]
  assign _T_1928 = _T_1927 & x772_b562_D2; // @[sm_x579_inr_Foreach.scala 141:228:@45260.4]
  assign _T_1929 = _T_1928 & x771_b552_D2; // @[sm_x579_inr_Foreach.scala 141:236:@45261.4]
  assign _T_1966 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@45332.4 package.scala 96:25:@45333.4]
  assign _T_1968 = io_rr ? _T_1966 : 1'h0; // @[implicits.scala 56:10:@45334.4]
  assign _T_1969 = _T_1876 & _T_1968; // @[sm_x579_inr_Foreach.scala 160:115:@45335.4]
  assign _T_1971 = _T_1969 & _T_1876; // @[sm_x579_inr_Foreach.scala 160:212:@45337.4]
  assign x774_b562_D5 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@45298.4 package.scala 96:25:@45299.4]
  assign _T_1973 = _T_1971 & x774_b562_D5; // @[sm_x579_inr_Foreach.scala 160:257:@45339.4]
  assign x775_b552_D5 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@45308.4 package.scala 96:25:@45309.4]
  assign _T_1974 = _T_1973 & x775_b552_D5; // @[sm_x579_inr_Foreach.scala 160:265:@45340.4]
  assign x776_b543_D5 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@45318.4 package.scala 96:25:@45319.4]
  assign _T_1986 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@45358.4 package.scala 96:25:@45359.4]
  assign _T_1988 = io_rr ? _T_1986 : 1'h0; // @[implicits.scala 56:10:@45360.4]
  assign _T_1989 = _T_1876 & _T_1988; // @[sm_x579_inr_Foreach.scala 165:115:@45361.4]
  assign _T_1991 = _T_1989 & _T_1876; // @[sm_x579_inr_Foreach.scala 165:212:@45363.4]
  assign _T_1993 = _T_1991 & x774_b562_D5; // @[sm_x579_inr_Foreach.scala 165:257:@45365.4]
  assign _T_1994 = _T_1993 & x775_b552_D5; // @[sm_x579_inr_Foreach.scala 165:265:@45366.4]
  assign _T_2006 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@45384.4 package.scala 96:25:@45385.4]
  assign _T_2008 = io_rr ? _T_2006 : 1'h0; // @[implicits.scala 56:10:@45386.4]
  assign _T_2009 = _T_1876 & _T_2008; // @[sm_x579_inr_Foreach.scala 170:115:@45387.4]
  assign _T_2011 = _T_2009 & _T_1876; // @[sm_x579_inr_Foreach.scala 170:212:@45389.4]
  assign _T_2013 = _T_2011 & x774_b562_D5; // @[sm_x579_inr_Foreach.scala 170:257:@45391.4]
  assign _T_2014 = _T_2013 & x775_b552_D5; // @[sm_x579_inr_Foreach.scala 170:265:@45392.4]
  assign _T_2026 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@45410.4 package.scala 96:25:@45411.4]
  assign _T_2028 = io_rr ? _T_2026 : 1'h0; // @[implicits.scala 56:10:@45412.4]
  assign _T_2029 = _T_1876 & _T_2028; // @[sm_x579_inr_Foreach.scala 175:115:@45413.4]
  assign _T_2031 = _T_2029 & _T_1876; // @[sm_x579_inr_Foreach.scala 175:212:@45415.4]
  assign _T_2033 = _T_2031 & x774_b562_D5; // @[sm_x579_inr_Foreach.scala 175:257:@45417.4]
  assign _T_2034 = _T_2033 & x775_b552_D5; // @[sm_x579_inr_Foreach.scala 175:265:@45418.4]
  assign _T_2046 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@45436.4 package.scala 96:25:@45437.4]
  assign _T_2048 = io_rr ? _T_2046 : 1'h0; // @[implicits.scala 56:10:@45438.4]
  assign _T_2049 = _T_1876 & _T_2048; // @[sm_x579_inr_Foreach.scala 180:115:@45439.4]
  assign _T_2051 = _T_2049 & _T_1876; // @[sm_x579_inr_Foreach.scala 180:212:@45441.4]
  assign _T_2053 = _T_2051 & x774_b562_D5; // @[sm_x579_inr_Foreach.scala 180:257:@45443.4]
  assign _T_2054 = _T_2053 & x775_b552_D5; // @[sm_x579_inr_Foreach.scala 180:265:@45444.4]
  assign _T_2059 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@45457.4 package.scala 96:25:@45458.4]
  assign _T_2065 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@45468.4 package.scala 96:25:@45469.4]
  assign _T_2071 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@45479.4 package.scala 96:25:@45480.4]
  assign _T_2077 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@45490.4 package.scala 96:25:@45491.4]
  assign _T_2083 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@45501.4 package.scala 96:25:@45502.4]
  assign x565_sum_number = x565_sum_1_io_result; // @[Math.scala 154:22:@45141.4 Math.scala 155:14:@45142.4]
  assign x570_sum_number = x570_sum_1_io_result; // @[Math.scala 154:22:@45232.4 Math.scala 155:14:@45233.4]
  assign x773_b561_D5_number = RetimeWrapper_8_io_out; // @[package.scala 96:25:@45288.4 package.scala 96:25:@45289.4]
  assign io_in_x555_tmp_1_wPort_0_ofs_0 = x773_b561_D5_number[1:0]; // @[MemInterfaceType.scala 89:54:@45343.4]
  assign io_in_x555_tmp_1_wPort_0_data_0 = x573_sub_1_io_result; // @[MemInterfaceType.scala 90:56:@45344.4]
  assign io_in_x555_tmp_1_wPort_0_en_0 = _T_1974 & x776_b543_D5; // @[MemInterfaceType.scala 93:57:@45346.4]
  assign io_in_x555_tmp_1_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@45471.4]
  assign io_in_x555_tmp_1_sDone_0 = io_rr ? _T_2065 : 1'h0; // @[MemInterfaceType.scala 197:17:@45472.4]
  assign io_in_x472_A_sram_1_rPort_0_ofs_0 = x570_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@45265.4]
  assign io_in_x472_A_sram_1_rPort_0_en_0 = _T_1929 & x770_b543_D2; // @[MemInterfaceType.scala 110:79:@45267.4]
  assign io_in_x471_A_sram_0_rPort_0_ofs_0 = x565_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@45204.4]
  assign io_in_x471_A_sram_0_rPort_0_en_0 = _T_1887 & x770_b543_D2; // @[MemInterfaceType.scala 110:79:@45206.4]
  assign io_in_x554_tmp_0_wPort_0_ofs_0 = x773_b561_D5_number[1:0]; // @[MemInterfaceType.scala 89:54:@45369.4]
  assign io_in_x554_tmp_0_wPort_0_data_0 = x573_sub_1_io_result; // @[MemInterfaceType.scala 90:56:@45370.4]
  assign io_in_x554_tmp_0_wPort_0_en_0 = _T_1994 & x776_b543_D5; // @[MemInterfaceType.scala 93:57:@45372.4]
  assign io_in_x554_tmp_0_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@45460.4]
  assign io_in_x554_tmp_0_sDone_0 = io_rr ? _T_2059 : 1'h0; // @[MemInterfaceType.scala 197:17:@45461.4]
  assign io_in_x558_tmp_4_wPort_0_ofs_0 = x773_b561_D5_number[1:0]; // @[MemInterfaceType.scala 89:54:@45395.4]
  assign io_in_x558_tmp_4_wPort_0_data_0 = x573_sub_1_io_result; // @[MemInterfaceType.scala 90:56:@45396.4]
  assign io_in_x558_tmp_4_wPort_0_en_0 = _T_2014 & x776_b543_D5; // @[MemInterfaceType.scala 93:57:@45398.4]
  assign io_in_x558_tmp_4_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@45504.4]
  assign io_in_x558_tmp_4_sDone_0 = io_rr ? _T_2083 : 1'h0; // @[MemInterfaceType.scala 197:17:@45505.4]
  assign io_in_x557_tmp_3_wPort_0_ofs_0 = x773_b561_D5_number[1:0]; // @[MemInterfaceType.scala 89:54:@45421.4]
  assign io_in_x557_tmp_3_wPort_0_data_0 = x573_sub_1_io_result; // @[MemInterfaceType.scala 90:56:@45422.4]
  assign io_in_x557_tmp_3_wPort_0_en_0 = _T_2034 & x776_b543_D5; // @[MemInterfaceType.scala 93:57:@45424.4]
  assign io_in_x557_tmp_3_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@45493.4]
  assign io_in_x557_tmp_3_sDone_0 = io_rr ? _T_2077 : 1'h0; // @[MemInterfaceType.scala 197:17:@45494.4]
  assign io_in_x556_tmp_2_wPort_0_ofs_0 = x773_b561_D5_number[1:0]; // @[MemInterfaceType.scala 89:54:@45447.4]
  assign io_in_x556_tmp_2_wPort_0_data_0 = x573_sub_1_io_result; // @[MemInterfaceType.scala 90:56:@45448.4]
  assign io_in_x556_tmp_2_wPort_0_en_0 = _T_2054 & x776_b543_D5; // @[MemInterfaceType.scala 93:57:@45450.4]
  assign io_in_x556_tmp_2_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@45482.4]
  assign io_in_x556_tmp_2_sDone_0 = io_rr ? _T_2071 : 1'h0; // @[MemInterfaceType.scala 197:17:@45483.4]
  assign io_in_instrctrs_8_cycs = cycles_x579_inr_Foreach_io_count; // @[Ledger.scala 293:21:@45092.4]
  assign io_in_instrctrs_8_iters = iters_x579_inr_Foreach_io_count; // @[Ledger.scala 294:22:@45093.4]
  assign cycles_x579_inr_Foreach_clock = clock; // @[:@45081.4]
  assign cycles_x579_inr_Foreach_reset = reset; // @[:@45082.4]
  assign cycles_x579_inr_Foreach_io_enable = io_sigsIn_baseEn; // @[sm_x579_inr_Foreach.scala 103:41:@45086.4]
  assign iters_x579_inr_Foreach_clock = clock; // @[:@45084.4]
  assign iters_x579_inr_Foreach_reset = reset; // @[:@45085.4]
  assign iters_x579_inr_Foreach_io_enable = io_sigsIn_done & _T_1817; // @[sm_x579_inr_Foreach.scala 104:40:@45091.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@45103.4]
  assign x745_sum_1_clock = clock; // @[:@45116.4]
  assign x745_sum_1_reset = reset; // @[:@45117.4]
  assign x745_sum_1_io_a = _T_1831[31:0]; // @[Math.scala 151:17:@45118.4]
  assign x745_sum_1_io_b = io_in_b542_number; // @[Math.scala 152:17:@45119.4]
  assign x745_sum_1_io_flow = 1'h1; // @[Math.scala 153:20:@45120.4]
  assign RetimeWrapper_clock = clock; // @[:@45127.4]
  assign RetimeWrapper_reset = reset; // @[:@45128.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@45130.4]
  assign RetimeWrapper_io_in = __io_result; // @[package.scala 94:16:@45129.4]
  assign x565_sum_1_clock = clock; // @[:@45136.4]
  assign x565_sum_1_reset = reset; // @[:@45137.4]
  assign x565_sum_1_io_a = x745_sum_1_io_result; // @[Math.scala 151:17:@45138.4]
  assign x565_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@45139.4]
  assign x565_sum_1_io_flow = 1'h1; // @[Math.scala 153:20:@45140.4]
  assign RetimeWrapper_1_clock = clock; // @[:@45147.4]
  assign RetimeWrapper_1_reset = reset; // @[:@45148.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@45150.4]
  assign RetimeWrapper_1_io_in = io_in_b543; // @[package.scala 94:16:@45149.4]
  assign RetimeWrapper_2_clock = clock; // @[:@45157.4]
  assign RetimeWrapper_2_reset = reset; // @[:@45158.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@45160.4]
  assign RetimeWrapper_2_io_in = io_in_b552; // @[package.scala 94:16:@45159.4]
  assign RetimeWrapper_3_clock = clock; // @[:@45167.4]
  assign RetimeWrapper_3_reset = reset; // @[:@45168.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@45170.4]
  assign RetimeWrapper_3_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@45169.4]
  assign RetimeWrapper_4_clock = clock; // @[:@45179.4]
  assign RetimeWrapper_4_reset = reset; // @[:@45180.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@45182.4]
  assign RetimeWrapper_4_io_in = 1'h1; // @[package.scala 94:16:@45181.4]
  assign RetimeWrapper_5_clock = clock; // @[:@45191.4]
  assign RetimeWrapper_5_reset = reset; // @[:@45192.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@45194.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45193.4]
  assign x747_sum_1_clock = clock; // @[:@45217.4]
  assign x747_sum_1_reset = reset; // @[:@45218.4]
  assign x747_sum_1_io_a = _T_1893[31:0]; // @[Math.scala 151:17:@45219.4]
  assign x747_sum_1_io_b = io_in_b550_number; // @[Math.scala 152:17:@45220.4]
  assign x747_sum_1_io_flow = 1'h1; // @[Math.scala 153:20:@45221.4]
  assign x570_sum_1_clock = clock; // @[:@45227.4]
  assign x570_sum_1_reset = reset; // @[:@45228.4]
  assign x570_sum_1_io_a = x747_sum_1_io_result; // @[Math.scala 151:17:@45229.4]
  assign x570_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@45230.4]
  assign x570_sum_1_io_flow = 1'h1; // @[Math.scala 153:20:@45231.4]
  assign RetimeWrapper_6_clock = clock; // @[:@45240.4]
  assign RetimeWrapper_6_reset = reset; // @[:@45241.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@45243.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@45242.4]
  assign RetimeWrapper_7_clock = clock; // @[:@45252.4]
  assign RetimeWrapper_7_reset = reset; // @[:@45253.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@45255.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45254.4]
  assign x573_sub_1_clock = clock; // @[:@45273.4]
  assign x573_sub_1_reset = reset; // @[:@45274.4]
  assign x573_sub_1_io_a = io_in_x471_A_sram_0_rPort_0_output_0; // @[Math.scala 192:17:@45275.4]
  assign x573_sub_1_io_b = io_in_x472_A_sram_1_rPort_0_output_0; // @[Math.scala 193:17:@45276.4]
  assign RetimeWrapper_8_clock = clock; // @[:@45284.4]
  assign RetimeWrapper_8_reset = reset; // @[:@45285.4]
  assign RetimeWrapper_8_io_in = __io_result; // @[package.scala 94:16:@45286.4]
  assign RetimeWrapper_9_clock = clock; // @[:@45294.4]
  assign RetimeWrapper_9_reset = reset; // @[:@45295.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@45297.4]
  assign RetimeWrapper_9_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@45296.4]
  assign RetimeWrapper_10_clock = clock; // @[:@45304.4]
  assign RetimeWrapper_10_reset = reset; // @[:@45305.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@45307.4]
  assign RetimeWrapper_10_io_in = io_in_b552; // @[package.scala 94:16:@45306.4]
  assign RetimeWrapper_11_clock = clock; // @[:@45314.4]
  assign RetimeWrapper_11_reset = reset; // @[:@45315.4]
  assign RetimeWrapper_11_io_flow = 1'h1; // @[package.scala 95:18:@45317.4]
  assign RetimeWrapper_11_io_in = io_in_b543; // @[package.scala 94:16:@45316.4]
  assign RetimeWrapper_12_clock = clock; // @[:@45328.4]
  assign RetimeWrapper_12_reset = reset; // @[:@45329.4]
  assign RetimeWrapper_12_io_flow = 1'h1; // @[package.scala 95:18:@45331.4]
  assign RetimeWrapper_12_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45330.4]
  assign RetimeWrapper_13_clock = clock; // @[:@45354.4]
  assign RetimeWrapper_13_reset = reset; // @[:@45355.4]
  assign RetimeWrapper_13_io_flow = 1'h1; // @[package.scala 95:18:@45357.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45356.4]
  assign RetimeWrapper_14_clock = clock; // @[:@45380.4]
  assign RetimeWrapper_14_reset = reset; // @[:@45381.4]
  assign RetimeWrapper_14_io_flow = 1'h1; // @[package.scala 95:18:@45383.4]
  assign RetimeWrapper_14_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45382.4]
  assign RetimeWrapper_15_clock = clock; // @[:@45406.4]
  assign RetimeWrapper_15_reset = reset; // @[:@45407.4]
  assign RetimeWrapper_15_io_flow = 1'h1; // @[package.scala 95:18:@45409.4]
  assign RetimeWrapper_15_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45408.4]
  assign RetimeWrapper_16_clock = clock; // @[:@45432.4]
  assign RetimeWrapper_16_reset = reset; // @[:@45433.4]
  assign RetimeWrapper_16_io_flow = 1'h1; // @[package.scala 95:18:@45435.4]
  assign RetimeWrapper_16_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@45434.4]
  assign RetimeWrapper_17_clock = clock; // @[:@45453.4]
  assign RetimeWrapper_17_reset = reset; // @[:@45454.4]
  assign RetimeWrapper_17_io_flow = 1'h1; // @[package.scala 95:18:@45456.4]
  assign RetimeWrapper_17_io_in = io_sigsIn_done; // @[package.scala 94:16:@45455.4]
  assign RetimeWrapper_18_clock = clock; // @[:@45464.4]
  assign RetimeWrapper_18_reset = reset; // @[:@45465.4]
  assign RetimeWrapper_18_io_flow = 1'h1; // @[package.scala 95:18:@45467.4]
  assign RetimeWrapper_18_io_in = io_sigsIn_done; // @[package.scala 94:16:@45466.4]
  assign RetimeWrapper_19_clock = clock; // @[:@45475.4]
  assign RetimeWrapper_19_reset = reset; // @[:@45476.4]
  assign RetimeWrapper_19_io_flow = 1'h1; // @[package.scala 95:18:@45478.4]
  assign RetimeWrapper_19_io_in = io_sigsIn_done; // @[package.scala 94:16:@45477.4]
  assign RetimeWrapper_20_clock = clock; // @[:@45486.4]
  assign RetimeWrapper_20_reset = reset; // @[:@45487.4]
  assign RetimeWrapper_20_io_flow = 1'h1; // @[package.scala 95:18:@45489.4]
  assign RetimeWrapper_20_io_in = io_sigsIn_done; // @[package.scala 94:16:@45488.4]
  assign RetimeWrapper_21_clock = clock; // @[:@45497.4]
  assign RetimeWrapper_21_reset = reset; // @[:@45498.4]
  assign RetimeWrapper_21_io_flow = 1'h1; // @[package.scala 95:18:@45500.4]
  assign RetimeWrapper_21_io_in = io_sigsIn_done; // @[package.scala 94:16:@45499.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1817 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1817 <= 1'h0;
    end else begin
      _T_1817 <= _T_1814;
    end
  end
endmodule
module RetimeWrapper_501( // @[:@45981.2]
  input         clock, // @[:@45982.4]
  input         reset, // @[:@45983.4]
  input         io_flow, // @[:@45984.4]
  input  [31:0] io_in, // @[:@45984.4]
  output [31:0] io_out // @[:@45984.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@45986.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@45986.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@45986.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@45986.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@45986.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@45986.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@45986.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@45999.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@45998.4]
  assign sr_init = 32'h2; // @[RetimeShiftRegister.scala 19:16:@45997.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@45996.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@45995.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@45993.4]
endmodule
module NBufCtr_66( // @[:@46001.2]
  input         clock, // @[:@46002.4]
  input         reset, // @[:@46003.4]
  input         io_input_enable, // @[:@46004.4]
  output [31:0] io_output_count // @[:@46004.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@46041.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@46041.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@46041.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@46041.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@46041.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@46046.4 package.scala 96:25:@46047.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@46007.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@46008.4]
  wire  _T_21; // @[Counter.scala 49:55:@46009.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@46010.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@46011.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@46012.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@46013.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@46014.4]
  wire  _T_33; // @[Counter.scala 51:52:@46018.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@46019.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@46020.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@46021.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@46022.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@46023.4]
  RetimeWrapper_501 RetimeWrapper ( // @[package.scala 93:22:@46041.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@46046.4 package.scala 96:25:@46047.4]
  assign _T_18 = {{1'd0}, _T_66}; // @[Counter.scala 49:32:@46007.4]
  assign _T_19 = _T_18[31:0]; // @[Counter.scala 49:32:@46008.4]
  assign _T_21 = _T_19 >= 32'h3; // @[Counter.scala 49:55:@46009.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@46010.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh3); // @[Counter.scala 49:91:@46011.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh3); // @[Counter.scala 49:91:@46012.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@46013.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@46014.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@46018.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@46019.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@46020.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@46021.4]
  assign _T_39 = _T_33 ? 32'h2 : _T_38; // @[Counter.scala 51:47:@46022.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@46023.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@46049.4]
  assign RetimeWrapper_clock = clock; // @[:@46042.4]
  assign RetimeWrapper_reset = reset; // @[:@46043.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@46045.4]
  assign RetimeWrapper_io_in = reset ? 32'h2 : _T_40; // @[package.scala 94:16:@46044.4]
endmodule
module NBufCtr_68( // @[:@46165.2]
  input         clock, // @[:@46166.4]
  input         reset, // @[:@46167.4]
  input         io_input_enable, // @[:@46168.4]
  output [31:0] io_output_count // @[:@46168.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@46205.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@46205.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@46205.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@46205.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@46205.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@46210.4 package.scala 96:25:@46211.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@46171.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@46172.4]
  wire  _T_21; // @[Counter.scala 49:55:@46173.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@46174.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@46175.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@46176.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@46177.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@46178.4]
  wire  _T_33; // @[Counter.scala 51:52:@46182.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@46183.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@46184.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@46185.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@46186.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@46187.4]
  RetimeWrapper_501 RetimeWrapper ( // @[package.scala 93:22:@46205.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@46210.4 package.scala 96:25:@46211.4]
  assign _T_18 = _T_66 + 32'h1; // @[Counter.scala 49:32:@46171.4]
  assign _T_19 = _T_66 + 32'h1; // @[Counter.scala 49:32:@46172.4]
  assign _T_21 = _T_19 >= 32'h3; // @[Counter.scala 49:55:@46173.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@46174.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh2); // @[Counter.scala 49:91:@46175.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh2); // @[Counter.scala 49:91:@46176.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@46177.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@46178.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@46182.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@46183.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@46184.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@46185.4]
  assign _T_39 = _T_33 ? 32'h2 : _T_38; // @[Counter.scala 51:47:@46186.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@46187.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@46213.4]
  assign RetimeWrapper_clock = clock; // @[:@46206.4]
  assign RetimeWrapper_reset = reset; // @[:@46207.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@46209.4]
  assign RetimeWrapper_io_in = reset ? 32'h2 : _T_40; // @[package.scala 94:16:@46208.4]
endmodule
module NBufCtr_69( // @[:@46247.2]
  input         clock, // @[:@46248.4]
  input         reset, // @[:@46249.4]
  input         io_input_enable, // @[:@46250.4]
  output [31:0] io_output_count // @[:@46250.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@46287.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@46287.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@46287.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@46287.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@46287.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@46292.4 package.scala 96:25:@46293.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@46253.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@46254.4]
  wire  _T_21; // @[Counter.scala 49:55:@46255.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@46256.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@46257.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@46258.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@46259.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@46260.4]
  wire  _T_33; // @[Counter.scala 51:52:@46264.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@46265.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@46266.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@46267.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@46268.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@46269.4]
  RetimeWrapper_501 RetimeWrapper ( // @[package.scala 93:22:@46287.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@46292.4 package.scala 96:25:@46293.4]
  assign _T_18 = _T_66 + 32'h2; // @[Counter.scala 49:32:@46253.4]
  assign _T_19 = _T_66 + 32'h2; // @[Counter.scala 49:32:@46254.4]
  assign _T_21 = _T_19 >= 32'h3; // @[Counter.scala 49:55:@46255.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@46256.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 49:91:@46257.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 49:91:@46258.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@46259.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@46260.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@46264.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@46265.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@46266.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@46267.4]
  assign _T_39 = _T_33 ? 32'h2 : _T_38; // @[Counter.scala 51:47:@46268.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@46269.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@46295.4]
  assign RetimeWrapper_clock = clock; // @[:@46288.4]
  assign RetimeWrapper_reset = reset; // @[:@46289.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@46291.4]
  assign RetimeWrapper_io_in = reset ? 32'h2 : _T_40; // @[package.scala 94:16:@46290.4]
endmodule
module NBufController_10( // @[:@46297.2]
  input        clock, // @[:@46298.4]
  input        reset, // @[:@46299.4]
  input        io_sEn_0, // @[:@46300.4]
  input        io_sEn_1, // @[:@46300.4]
  input        io_sEn_2, // @[:@46300.4]
  input        io_sDone_0, // @[:@46300.4]
  input        io_sDone_1, // @[:@46300.4]
  input        io_sDone_2, // @[:@46300.4]
  output [2:0] io_statesInW_0, // @[:@46300.4]
  output [2:0] io_statesInR_1, // @[:@46300.4]
  output [2:0] io_statesInR_2 // @[:@46300.4]
);
  wire  sEn_latch_0_clock; // @[NBuffers.scala 21:52:@46302.4]
  wire  sEn_latch_0_reset; // @[NBuffers.scala 21:52:@46302.4]
  wire  sEn_latch_0_io_input_set; // @[NBuffers.scala 21:52:@46302.4]
  wire  sEn_latch_0_io_input_reset; // @[NBuffers.scala 21:52:@46302.4]
  wire  sEn_latch_0_io_input_asyn_reset; // @[NBuffers.scala 21:52:@46302.4]
  wire  sEn_latch_0_io_output; // @[NBuffers.scala 21:52:@46302.4]
  wire  sEn_latch_1_clock; // @[NBuffers.scala 21:52:@46305.4]
  wire  sEn_latch_1_reset; // @[NBuffers.scala 21:52:@46305.4]
  wire  sEn_latch_1_io_input_set; // @[NBuffers.scala 21:52:@46305.4]
  wire  sEn_latch_1_io_input_reset; // @[NBuffers.scala 21:52:@46305.4]
  wire  sEn_latch_1_io_input_asyn_reset; // @[NBuffers.scala 21:52:@46305.4]
  wire  sEn_latch_1_io_output; // @[NBuffers.scala 21:52:@46305.4]
  wire  sEn_latch_2_clock; // @[NBuffers.scala 21:52:@46308.4]
  wire  sEn_latch_2_reset; // @[NBuffers.scala 21:52:@46308.4]
  wire  sEn_latch_2_io_input_set; // @[NBuffers.scala 21:52:@46308.4]
  wire  sEn_latch_2_io_input_reset; // @[NBuffers.scala 21:52:@46308.4]
  wire  sEn_latch_2_io_input_asyn_reset; // @[NBuffers.scala 21:52:@46308.4]
  wire  sEn_latch_2_io_output; // @[NBuffers.scala 21:52:@46308.4]
  wire  sDone_latch_0_clock; // @[NBuffers.scala 22:54:@46311.4]
  wire  sDone_latch_0_reset; // @[NBuffers.scala 22:54:@46311.4]
  wire  sDone_latch_0_io_input_set; // @[NBuffers.scala 22:54:@46311.4]
  wire  sDone_latch_0_io_input_reset; // @[NBuffers.scala 22:54:@46311.4]
  wire  sDone_latch_0_io_input_asyn_reset; // @[NBuffers.scala 22:54:@46311.4]
  wire  sDone_latch_0_io_output; // @[NBuffers.scala 22:54:@46311.4]
  wire  sDone_latch_1_clock; // @[NBuffers.scala 22:54:@46314.4]
  wire  sDone_latch_1_reset; // @[NBuffers.scala 22:54:@46314.4]
  wire  sDone_latch_1_io_input_set; // @[NBuffers.scala 22:54:@46314.4]
  wire  sDone_latch_1_io_input_reset; // @[NBuffers.scala 22:54:@46314.4]
  wire  sDone_latch_1_io_input_asyn_reset; // @[NBuffers.scala 22:54:@46314.4]
  wire  sDone_latch_1_io_output; // @[NBuffers.scala 22:54:@46314.4]
  wire  sDone_latch_2_clock; // @[NBuffers.scala 22:54:@46317.4]
  wire  sDone_latch_2_reset; // @[NBuffers.scala 22:54:@46317.4]
  wire  sDone_latch_2_io_input_set; // @[NBuffers.scala 22:54:@46317.4]
  wire  sDone_latch_2_io_input_reset; // @[NBuffers.scala 22:54:@46317.4]
  wire  sDone_latch_2_io_input_asyn_reset; // @[NBuffers.scala 22:54:@46317.4]
  wire  sDone_latch_2_io_output; // @[NBuffers.scala 22:54:@46317.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@46324.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@46324.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@46324.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@46324.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@46324.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@46332.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@46332.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@46332.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@46332.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@46332.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@46341.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@46341.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@46341.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@46341.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@46341.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@46349.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@46349.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@46349.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@46349.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@46349.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@46360.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@46360.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@46360.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@46360.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@46360.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@46368.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@46368.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@46368.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@46368.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@46368.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@46377.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@46377.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@46377.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@46377.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@46377.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@46385.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@46385.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@46385.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@46385.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@46385.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@46396.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@46396.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@46396.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@46396.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@46396.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@46404.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@46404.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@46404.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@46404.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@46404.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@46413.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@46413.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@46413.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@46413.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@46413.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@46421.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@46421.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@46421.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@46421.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@46421.4]
  wire  NBufCtr_clock; // @[NBuffers.scala 40:19:@46446.4]
  wire  NBufCtr_reset; // @[NBuffers.scala 40:19:@46446.4]
  wire  NBufCtr_io_input_enable; // @[NBuffers.scala 40:19:@46446.4]
  wire [31:0] NBufCtr_io_output_count; // @[NBuffers.scala 40:19:@46446.4]
  wire  statesInR_0_clock; // @[NBuffers.scala 50:19:@46457.4]
  wire  statesInR_0_reset; // @[NBuffers.scala 50:19:@46457.4]
  wire  statesInR_0_io_input_enable; // @[NBuffers.scala 50:19:@46457.4]
  wire [31:0] statesInR_0_io_output_count; // @[NBuffers.scala 50:19:@46457.4]
  wire  statesInR_1_clock; // @[NBuffers.scala 50:19:@46468.4]
  wire  statesInR_1_reset; // @[NBuffers.scala 50:19:@46468.4]
  wire  statesInR_1_io_input_enable; // @[NBuffers.scala 50:19:@46468.4]
  wire [31:0] statesInR_1_io_output_count; // @[NBuffers.scala 50:19:@46468.4]
  wire  statesInR_2_clock; // @[NBuffers.scala 50:19:@46479.4]
  wire  statesInR_2_reset; // @[NBuffers.scala 50:19:@46479.4]
  wire  statesInR_2_io_input_enable; // @[NBuffers.scala 50:19:@46479.4]
  wire [31:0] statesInR_2_io_output_count; // @[NBuffers.scala 50:19:@46479.4]
  wire  _T_33; // @[NBuffers.scala 26:46:@46321.4]
  wire  _T_48; // @[NBuffers.scala 26:46:@46357.4]
  wire  _T_63; // @[NBuffers.scala 26:46:@46393.4]
  wire  _T_77; // @[NBuffers.scala 33:64:@46429.4]
  wire  anyEnabled; // @[NBuffers.scala 33:64:@46430.4]
  wire  _T_78; // @[NBuffers.scala 34:124:@46431.4]
  wire  _T_79; // @[NBuffers.scala 34:104:@46432.4]
  wire  _T_80; // @[NBuffers.scala 34:124:@46433.4]
  wire  _T_81; // @[NBuffers.scala 34:104:@46434.4]
  wire  _T_82; // @[NBuffers.scala 34:124:@46435.4]
  wire  _T_83; // @[NBuffers.scala 34:104:@46436.4]
  wire  _T_84; // @[NBuffers.scala 34:150:@46437.4]
  wire  _T_85; // @[NBuffers.scala 34:150:@46438.4]
  wire  _T_86; // @[NBuffers.scala 34:154:@46439.4]
  wire  _T_88; // @[package.scala 100:49:@46440.4]
  reg  _T_91; // @[package.scala 48:56:@46441.4]
  reg [31:0] _RAND_0;
  SRFF sEn_latch_0 ( // @[NBuffers.scala 21:52:@46302.4]
    .clock(sEn_latch_0_clock),
    .reset(sEn_latch_0_reset),
    .io_input_set(sEn_latch_0_io_input_set),
    .io_input_reset(sEn_latch_0_io_input_reset),
    .io_input_asyn_reset(sEn_latch_0_io_input_asyn_reset),
    .io_output(sEn_latch_0_io_output)
  );
  SRFF sEn_latch_1 ( // @[NBuffers.scala 21:52:@46305.4]
    .clock(sEn_latch_1_clock),
    .reset(sEn_latch_1_reset),
    .io_input_set(sEn_latch_1_io_input_set),
    .io_input_reset(sEn_latch_1_io_input_reset),
    .io_input_asyn_reset(sEn_latch_1_io_input_asyn_reset),
    .io_output(sEn_latch_1_io_output)
  );
  SRFF sEn_latch_2 ( // @[NBuffers.scala 21:52:@46308.4]
    .clock(sEn_latch_2_clock),
    .reset(sEn_latch_2_reset),
    .io_input_set(sEn_latch_2_io_input_set),
    .io_input_reset(sEn_latch_2_io_input_reset),
    .io_input_asyn_reset(sEn_latch_2_io_input_asyn_reset),
    .io_output(sEn_latch_2_io_output)
  );
  SRFF sDone_latch_0 ( // @[NBuffers.scala 22:54:@46311.4]
    .clock(sDone_latch_0_clock),
    .reset(sDone_latch_0_reset),
    .io_input_set(sDone_latch_0_io_input_set),
    .io_input_reset(sDone_latch_0_io_input_reset),
    .io_input_asyn_reset(sDone_latch_0_io_input_asyn_reset),
    .io_output(sDone_latch_0_io_output)
  );
  SRFF sDone_latch_1 ( // @[NBuffers.scala 22:54:@46314.4]
    .clock(sDone_latch_1_clock),
    .reset(sDone_latch_1_reset),
    .io_input_set(sDone_latch_1_io_input_set),
    .io_input_reset(sDone_latch_1_io_input_reset),
    .io_input_asyn_reset(sDone_latch_1_io_input_asyn_reset),
    .io_output(sDone_latch_1_io_output)
  );
  SRFF sDone_latch_2 ( // @[NBuffers.scala 22:54:@46317.4]
    .clock(sDone_latch_2_clock),
    .reset(sDone_latch_2_reset),
    .io_input_set(sDone_latch_2_io_input_set),
    .io_input_reset(sDone_latch_2_io_input_reset),
    .io_input_asyn_reset(sDone_latch_2_io_input_asyn_reset),
    .io_output(sDone_latch_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@46324.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@46332.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@46341.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@46349.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@46360.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@46368.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@46377.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@46385.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@46396.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@46404.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@46413.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 ( // @[package.scala 93:22:@46421.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  NBufCtr_66 NBufCtr ( // @[NBuffers.scala 40:19:@46446.4]
    .clock(NBufCtr_clock),
    .reset(NBufCtr_reset),
    .io_input_enable(NBufCtr_io_input_enable),
    .io_output_count(NBufCtr_io_output_count)
  );
  NBufCtr_66 statesInR_0 ( // @[NBuffers.scala 50:19:@46457.4]
    .clock(statesInR_0_clock),
    .reset(statesInR_0_reset),
    .io_input_enable(statesInR_0_io_input_enable),
    .io_output_count(statesInR_0_io_output_count)
  );
  NBufCtr_68 statesInR_1 ( // @[NBuffers.scala 50:19:@46468.4]
    .clock(statesInR_1_clock),
    .reset(statesInR_1_reset),
    .io_input_enable(statesInR_1_io_input_enable),
    .io_output_count(statesInR_1_io_output_count)
  );
  NBufCtr_69 statesInR_2 ( // @[NBuffers.scala 50:19:@46479.4]
    .clock(statesInR_2_clock),
    .reset(statesInR_2_reset),
    .io_input_enable(statesInR_2_io_input_enable),
    .io_output_count(statesInR_2_io_output_count)
  );
  assign _T_33 = io_sDone_0 == 1'h0; // @[NBuffers.scala 26:46:@46321.4]
  assign _T_48 = io_sDone_1 == 1'h0; // @[NBuffers.scala 26:46:@46357.4]
  assign _T_63 = io_sDone_2 == 1'h0; // @[NBuffers.scala 26:46:@46393.4]
  assign _T_77 = sEn_latch_0_io_output | sEn_latch_1_io_output; // @[NBuffers.scala 33:64:@46429.4]
  assign anyEnabled = _T_77 | sEn_latch_2_io_output; // @[NBuffers.scala 33:64:@46430.4]
  assign _T_78 = sDone_latch_0_io_output | io_sDone_0; // @[NBuffers.scala 34:124:@46431.4]
  assign _T_79 = sEn_latch_0_io_output == _T_78; // @[NBuffers.scala 34:104:@46432.4]
  assign _T_80 = sDone_latch_1_io_output | io_sDone_1; // @[NBuffers.scala 34:124:@46433.4]
  assign _T_81 = sEn_latch_1_io_output == _T_80; // @[NBuffers.scala 34:104:@46434.4]
  assign _T_82 = sDone_latch_2_io_output | io_sDone_2; // @[NBuffers.scala 34:124:@46435.4]
  assign _T_83 = sEn_latch_2_io_output == _T_82; // @[NBuffers.scala 34:104:@46436.4]
  assign _T_84 = _T_79 & _T_81; // @[NBuffers.scala 34:150:@46437.4]
  assign _T_85 = _T_84 & _T_83; // @[NBuffers.scala 34:150:@46438.4]
  assign _T_86 = _T_85 & anyEnabled; // @[NBuffers.scala 34:154:@46439.4]
  assign _T_88 = _T_86 == 1'h0; // @[package.scala 100:49:@46440.4]
  assign io_statesInW_0 = NBufCtr_io_output_count[2:0]; // @[NBuffers.scala 44:21:@46456.4]
  assign io_statesInR_1 = statesInR_1_io_output_count[2:0]; // @[NBuffers.scala 54:21:@46478.4]
  assign io_statesInR_2 = statesInR_2_io_output_count[2:0]; // @[NBuffers.scala 54:21:@46489.4]
  assign sEn_latch_0_clock = clock; // @[:@46303.4]
  assign sEn_latch_0_reset = reset; // @[:@46304.4]
  assign sEn_latch_0_io_input_set = io_sEn_0 & _T_33; // @[NBuffers.scala 26:31:@46323.4]
  assign sEn_latch_0_io_input_reset = RetimeWrapper_io_out; // @[NBuffers.scala 27:33:@46331.4]
  assign sEn_latch_0_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[NBuffers.scala 28:38:@46339.4]
  assign sEn_latch_1_clock = clock; // @[:@46306.4]
  assign sEn_latch_1_reset = reset; // @[:@46307.4]
  assign sEn_latch_1_io_input_set = io_sEn_1 & _T_48; // @[NBuffers.scala 26:31:@46359.4]
  assign sEn_latch_1_io_input_reset = RetimeWrapper_4_io_out; // @[NBuffers.scala 27:33:@46367.4]
  assign sEn_latch_1_io_input_asyn_reset = RetimeWrapper_5_io_out; // @[NBuffers.scala 28:38:@46375.4]
  assign sEn_latch_2_clock = clock; // @[:@46309.4]
  assign sEn_latch_2_reset = reset; // @[:@46310.4]
  assign sEn_latch_2_io_input_set = io_sEn_2 & _T_63; // @[NBuffers.scala 26:31:@46395.4]
  assign sEn_latch_2_io_input_reset = RetimeWrapper_8_io_out; // @[NBuffers.scala 27:33:@46403.4]
  assign sEn_latch_2_io_input_asyn_reset = RetimeWrapper_9_io_out; // @[NBuffers.scala 28:38:@46411.4]
  assign sDone_latch_0_clock = clock; // @[:@46312.4]
  assign sDone_latch_0_reset = reset; // @[:@46313.4]
  assign sDone_latch_0_io_input_set = io_sDone_0; // @[NBuffers.scala 29:33:@46340.4]
  assign sDone_latch_0_io_input_reset = RetimeWrapper_2_io_out; // @[NBuffers.scala 30:35:@46348.4]
  assign sDone_latch_0_io_input_asyn_reset = RetimeWrapper_3_io_out; // @[NBuffers.scala 31:40:@46356.4]
  assign sDone_latch_1_clock = clock; // @[:@46315.4]
  assign sDone_latch_1_reset = reset; // @[:@46316.4]
  assign sDone_latch_1_io_input_set = io_sDone_1; // @[NBuffers.scala 29:33:@46376.4]
  assign sDone_latch_1_io_input_reset = RetimeWrapper_6_io_out; // @[NBuffers.scala 30:35:@46384.4]
  assign sDone_latch_1_io_input_asyn_reset = RetimeWrapper_7_io_out; // @[NBuffers.scala 31:40:@46392.4]
  assign sDone_latch_2_clock = clock; // @[:@46318.4]
  assign sDone_latch_2_reset = reset; // @[:@46319.4]
  assign sDone_latch_2_io_input_set = io_sDone_2; // @[NBuffers.scala 29:33:@46412.4]
  assign sDone_latch_2_io_input_reset = RetimeWrapper_10_io_out; // @[NBuffers.scala 30:35:@46420.4]
  assign sDone_latch_2_io_input_asyn_reset = RetimeWrapper_11_io_out; // @[NBuffers.scala 31:40:@46428.4]
  assign RetimeWrapper_clock = clock; // @[:@46325.4]
  assign RetimeWrapper_reset = reset; // @[:@46326.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@46328.4]
  assign RetimeWrapper_io_in = _T_86 & _T_91; // @[package.scala 94:16:@46327.4]
  assign RetimeWrapper_1_clock = clock; // @[:@46333.4]
  assign RetimeWrapper_1_reset = reset; // @[:@46334.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@46336.4]
  assign RetimeWrapper_1_io_in = reset; // @[package.scala 94:16:@46335.4]
  assign RetimeWrapper_2_clock = clock; // @[:@46342.4]
  assign RetimeWrapper_2_reset = reset; // @[:@46343.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@46345.4]
  assign RetimeWrapper_2_io_in = _T_86 & _T_91; // @[package.scala 94:16:@46344.4]
  assign RetimeWrapper_3_clock = clock; // @[:@46350.4]
  assign RetimeWrapper_3_reset = reset; // @[:@46351.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@46353.4]
  assign RetimeWrapper_3_io_in = reset; // @[package.scala 94:16:@46352.4]
  assign RetimeWrapper_4_clock = clock; // @[:@46361.4]
  assign RetimeWrapper_4_reset = reset; // @[:@46362.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@46364.4]
  assign RetimeWrapper_4_io_in = _T_86 & _T_91; // @[package.scala 94:16:@46363.4]
  assign RetimeWrapper_5_clock = clock; // @[:@46369.4]
  assign RetimeWrapper_5_reset = reset; // @[:@46370.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@46372.4]
  assign RetimeWrapper_5_io_in = reset; // @[package.scala 94:16:@46371.4]
  assign RetimeWrapper_6_clock = clock; // @[:@46378.4]
  assign RetimeWrapper_6_reset = reset; // @[:@46379.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@46381.4]
  assign RetimeWrapper_6_io_in = _T_86 & _T_91; // @[package.scala 94:16:@46380.4]
  assign RetimeWrapper_7_clock = clock; // @[:@46386.4]
  assign RetimeWrapper_7_reset = reset; // @[:@46387.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@46389.4]
  assign RetimeWrapper_7_io_in = reset; // @[package.scala 94:16:@46388.4]
  assign RetimeWrapper_8_clock = clock; // @[:@46397.4]
  assign RetimeWrapper_8_reset = reset; // @[:@46398.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@46400.4]
  assign RetimeWrapper_8_io_in = _T_86 & _T_91; // @[package.scala 94:16:@46399.4]
  assign RetimeWrapper_9_clock = clock; // @[:@46405.4]
  assign RetimeWrapper_9_reset = reset; // @[:@46406.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@46408.4]
  assign RetimeWrapper_9_io_in = reset; // @[package.scala 94:16:@46407.4]
  assign RetimeWrapper_10_clock = clock; // @[:@46414.4]
  assign RetimeWrapper_10_reset = reset; // @[:@46415.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@46417.4]
  assign RetimeWrapper_10_io_in = _T_86 & _T_91; // @[package.scala 94:16:@46416.4]
  assign RetimeWrapper_11_clock = clock; // @[:@46422.4]
  assign RetimeWrapper_11_reset = reset; // @[:@46423.4]
  assign RetimeWrapper_11_io_flow = 1'h1; // @[package.scala 95:18:@46425.4]
  assign RetimeWrapper_11_io_in = reset; // @[package.scala 94:16:@46424.4]
  assign NBufCtr_clock = clock; // @[:@46447.4]
  assign NBufCtr_reset = reset; // @[:@46448.4]
  assign NBufCtr_io_input_enable = _T_86 & _T_91; // @[NBuffers.scala 42:23:@46454.4]
  assign statesInR_0_clock = clock; // @[:@46458.4]
  assign statesInR_0_reset = reset; // @[:@46459.4]
  assign statesInR_0_io_input_enable = _T_86 & _T_91; // @[NBuffers.scala 52:23:@46465.4]
  assign statesInR_1_clock = clock; // @[:@46469.4]
  assign statesInR_1_reset = reset; // @[:@46470.4]
  assign statesInR_1_io_input_enable = _T_86 & _T_91; // @[NBuffers.scala 52:23:@46476.4]
  assign statesInR_2_clock = clock; // @[:@46480.4]
  assign statesInR_2_reset = reset; // @[:@46481.4]
  assign statesInR_2_io_input_enable = _T_86 & _T_91; // @[NBuffers.scala 52:23:@46487.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_91 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_91 <= 1'h0;
    end else begin
      _T_91 <= _T_88;
    end
  end
endmodule
module Mem1D_39( // @[:@46555.2]
  input         clock, // @[:@46556.4]
  input         reset, // @[:@46557.4]
  input         io_r_ofs_0, // @[:@46558.4]
  input         io_r_backpressure, // @[:@46558.4]
  input         io_w_ofs_0, // @[:@46558.4]
  input  [31:0] io_w_data_0, // @[:@46558.4]
  input         io_w_en_0, // @[:@46558.4]
  output [31:0] io_output // @[:@46558.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@46568.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@46568.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@46568.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@46568.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@46568.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@46577.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@46577.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@46577.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@46577.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@46577.4]
  reg [31:0] _T_127; // @[MemPrimitives.scala 746:26:@46562.4]
  reg [31:0] _RAND_0;
  wire  _T_130; // @[MemPrimitives.scala 747:61:@46564.4]
  wire  _T_131; // @[MemPrimitives.scala 747:44:@46565.4]
  wire [31:0] _T_132; // @[MemPrimitives.scala 747:19:@46566.4]
  wire  _T_135; // @[package.scala 96:25:@46573.4 package.scala 96:25:@46574.4]
  wire  _T_137; // @[Mux.scala 46:19:@46575.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@46568.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_32 RetimeWrapper_1 ( // @[package.scala 93:22:@46577.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_130 = io_w_ofs_0 == 1'h0; // @[MemPrimitives.scala 747:61:@46564.4]
  assign _T_131 = io_w_en_0 & _T_130; // @[MemPrimitives.scala 747:44:@46565.4]
  assign _T_132 = _T_131 ? io_w_data_0 : _T_127; // @[MemPrimitives.scala 747:19:@46566.4]
  assign _T_135 = RetimeWrapper_io_out; // @[package.scala 96:25:@46573.4 package.scala 96:25:@46574.4]
  assign _T_137 = 1'h0 == _T_135; // @[Mux.scala 46:19:@46575.4]
  assign io_output = RetimeWrapper_1_io_out; // @[MemPrimitives.scala 751:17:@46584.4]
  assign RetimeWrapper_clock = clock; // @[:@46569.4]
  assign RetimeWrapper_reset = reset; // @[:@46570.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@46572.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@46571.4]
  assign RetimeWrapper_1_clock = clock; // @[:@46578.4]
  assign RetimeWrapper_1_reset = reset; // @[:@46579.4]
  assign RetimeWrapper_1_io_flow = io_r_backpressure; // @[package.scala 95:18:@46581.4]
  assign RetimeWrapper_1_io_in = _T_137 ? _T_127 : 32'h0; // @[package.scala 94:16:@46580.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_127 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_127 <= 32'h0;
    end else begin
      if (_T_131) begin
        _T_127 <= io_w_data_0;
      end
    end
  end
endmodule
module StickySelects_38( // @[:@46586.2]
  input   clock, // @[:@46587.4]
  input   reset, // @[:@46588.4]
  input   io_ins_0, // @[:@46589.4]
  input   io_ins_1, // @[:@46589.4]
  output  io_outs_0, // @[:@46589.4]
  output  io_outs_1 // @[:@46589.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@46591.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@46592.4]
  reg [31:0] _RAND_1;
  wire  _T_23; // @[StickySelects.scala 49:53:@46593.4]
  wire  _T_24; // @[StickySelects.scala 49:21:@46594.4]
  wire  _T_25; // @[StickySelects.scala 49:53:@46596.4]
  wire  _T_26; // @[StickySelects.scala 49:21:@46597.4]
  assign _T_23 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@46593.4]
  assign _T_24 = io_ins_1 ? io_ins_0 : _T_23; // @[StickySelects.scala 49:21:@46594.4]
  assign _T_25 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@46596.4]
  assign _T_26 = io_ins_0 ? io_ins_1 : _T_25; // @[StickySelects.scala 49:21:@46597.4]
  assign io_outs_0 = io_ins_1 ? io_ins_0 : _T_23; // @[StickySelects.scala 53:57:@46599.4]
  assign io_outs_1 = io_ins_0 ? io_ins_1 : _T_25; // @[StickySelects.scala 53:57:@46600.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (io_ins_1) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_23;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (io_ins_0) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_25;
      end
    end
  end
endmodule
module SRAM_71( // @[:@46666.2]
  input         clock, // @[:@46667.4]
  input         reset, // @[:@46668.4]
  input         io_rPort_1_en_0, // @[:@46669.4]
  output [31:0] io_rPort_1_output_0, // @[:@46669.4]
  input         io_rPort_0_en_0, // @[:@46669.4]
  output [31:0] io_rPort_0_output_0, // @[:@46669.4]
  input  [31:0] io_wPort_0_data_0, // @[:@46669.4]
  input         io_wPort_0_en_0 // @[:@46669.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@46689.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@46689.4]
  wire  Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@46689.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@46689.4]
  wire  Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@46689.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@46689.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@46689.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@46689.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@46716.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@46716.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@46716.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@46716.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@46716.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@46716.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@46735.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@46735.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@46735.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@46735.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@46735.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@46744.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@46744.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@46744.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@46744.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@46744.4]
  wire [33:0] _T_96; // @[Cat.scala 30:58:@46707.4]
  wire  _T_104; // @[MemPrimitives.scala 126:35:@46721.4]
  wire  _T_105; // @[MemPrimitives.scala 126:35:@46722.4]
  wire [2:0] _T_107; // @[Cat.scala 30:58:@46724.4]
  wire [2:0] _T_109; // @[Cat.scala 30:58:@46726.4]
  wire [2:0] _T_110; // @[Mux.scala 31:69:@46727.4]
  Mem1D_39 Mem1D ( // @[MemPrimitives.scala 64:21:@46689.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  StickySelects_38 StickySelects ( // @[MemPrimitives.scala 124:33:@46716.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@46735.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@46744.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_96 = {io_wPort_0_en_0,io_wPort_0_data_0,1'h0}; // @[Cat.scala 30:58:@46707.4]
  assign _T_104 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@46721.4]
  assign _T_105 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@46722.4]
  assign _T_107 = {_T_104,1'h1,1'h0}; // @[Cat.scala 30:58:@46724.4]
  assign _T_109 = {_T_105,1'h1,1'h0}; // @[Cat.scala 30:58:@46726.4]
  assign _T_110 = _T_104 ? _T_107 : _T_109; // @[Mux.scala 31:69:@46727.4]
  assign io_rPort_1_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@46751.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@46742.4]
  assign Mem1D_clock = clock; // @[:@46690.4]
  assign Mem1D_reset = reset; // @[:@46691.4]
  assign Mem1D_io_r_ofs_0 = _T_110[0]; // @[MemPrimitives.scala 131:28:@46731.4]
  assign Mem1D_io_r_backpressure = _T_110[1]; // @[MemPrimitives.scala 132:32:@46732.4]
  assign Mem1D_io_w_ofs_0 = _T_96[0]; // @[MemPrimitives.scala 94:28:@46711.4]
  assign Mem1D_io_w_data_0 = _T_96[32:1]; // @[MemPrimitives.scala 95:29:@46712.4]
  assign Mem1D_io_w_en_0 = _T_96[33]; // @[MemPrimitives.scala 96:27:@46713.4]
  assign StickySelects_clock = clock; // @[:@46717.4]
  assign StickySelects_reset = reset; // @[:@46718.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@46719.4]
  assign StickySelects_io_ins_1 = io_rPort_1_en_0; // @[MemPrimitives.scala 125:64:@46720.4]
  assign RetimeWrapper_clock = clock; // @[:@46736.4]
  assign RetimeWrapper_reset = reset; // @[:@46737.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@46739.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@46738.4]
  assign RetimeWrapper_1_clock = clock; // @[:@46745.4]
  assign RetimeWrapper_1_reset = reset; // @[:@46746.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@46748.4]
  assign RetimeWrapper_1_io_in = io_rPort_1_en_0; // @[package.scala 94:16:@46747.4]
endmodule
module x580_r_0( // @[:@47277.2]
  input         clock, // @[:@47278.4]
  input         reset, // @[:@47279.4]
  input         io_rPort_1_en_0, // @[:@47280.4]
  output [31:0] io_rPort_1_output_0, // @[:@47280.4]
  input         io_rPort_0_en_0, // @[:@47280.4]
  output [31:0] io_rPort_0_output_0, // @[:@47280.4]
  input  [31:0] io_wPort_0_data_0, // @[:@47280.4]
  input         io_wPort_0_en_0, // @[:@47280.4]
  input         io_sEn_0, // @[:@47280.4]
  input         io_sEn_1, // @[:@47280.4]
  input         io_sEn_2, // @[:@47280.4]
  input         io_sDone_0, // @[:@47280.4]
  input         io_sDone_1, // @[:@47280.4]
  input         io_sDone_2 // @[:@47280.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@47290.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@47290.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@47290.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@47290.4]
  wire  ctrl_io_sEn_2; // @[NBuffers.scala 83:20:@47290.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@47290.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@47290.4]
  wire  ctrl_io_sDone_2; // @[NBuffers.scala 83:20:@47290.4]
  wire [2:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@47290.4]
  wire [2:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@47290.4]
  wire [2:0] ctrl_io_statesInR_2; // @[NBuffers.scala 83:20:@47290.4]
  wire  SRAM_clock; // @[NBuffers.scala 94:23:@47299.4]
  wire  SRAM_reset; // @[NBuffers.scala 94:23:@47299.4]
  wire  SRAM_io_rPort_1_en_0; // @[NBuffers.scala 94:23:@47299.4]
  wire [31:0] SRAM_io_rPort_1_output_0; // @[NBuffers.scala 94:23:@47299.4]
  wire  SRAM_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@47299.4]
  wire [31:0] SRAM_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@47299.4]
  wire [31:0] SRAM_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@47299.4]
  wire  SRAM_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@47299.4]
  wire  SRAM_1_clock; // @[NBuffers.scala 94:23:@47320.4]
  wire  SRAM_1_reset; // @[NBuffers.scala 94:23:@47320.4]
  wire  SRAM_1_io_rPort_1_en_0; // @[NBuffers.scala 94:23:@47320.4]
  wire [31:0] SRAM_1_io_rPort_1_output_0; // @[NBuffers.scala 94:23:@47320.4]
  wire  SRAM_1_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@47320.4]
  wire [31:0] SRAM_1_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@47320.4]
  wire [31:0] SRAM_1_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@47320.4]
  wire  SRAM_1_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@47320.4]
  wire  SRAM_2_clock; // @[NBuffers.scala 94:23:@47341.4]
  wire  SRAM_2_reset; // @[NBuffers.scala 94:23:@47341.4]
  wire  SRAM_2_io_rPort_1_en_0; // @[NBuffers.scala 94:23:@47341.4]
  wire [31:0] SRAM_2_io_rPort_1_output_0; // @[NBuffers.scala 94:23:@47341.4]
  wire  SRAM_2_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@47341.4]
  wire [31:0] SRAM_2_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@47341.4]
  wire [31:0] SRAM_2_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@47341.4]
  wire  SRAM_2_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@47341.4]
  wire  _T_140; // @[NBuffers.scala 104:105:@47362.4]
  wire  _T_144; // @[NBuffers.scala 108:92:@47372.4]
  wire  _T_147; // @[NBuffers.scala 108:92:@47378.4]
  wire  _T_150; // @[NBuffers.scala 104:105:@47384.4]
  wire  _T_154; // @[NBuffers.scala 108:92:@47394.4]
  wire  _T_157; // @[NBuffers.scala 108:92:@47400.4]
  wire  _T_160; // @[NBuffers.scala 104:105:@47406.4]
  wire  _T_164; // @[NBuffers.scala 108:92:@47416.4]
  wire  _T_167; // @[NBuffers.scala 108:92:@47422.4]
  wire [31:0] _T_177; // @[Mux.scala 19:72:@47431.4]
  wire [31:0] _T_179; // @[Mux.scala 19:72:@47432.4]
  wire [31:0] _T_181; // @[Mux.scala 19:72:@47433.4]
  wire [31:0] _T_182; // @[Mux.scala 19:72:@47434.4]
  wire [31:0] _T_194; // @[Mux.scala 19:72:@47442.4]
  wire [31:0] _T_196; // @[Mux.scala 19:72:@47443.4]
  wire [31:0] _T_198; // @[Mux.scala 19:72:@47444.4]
  wire [31:0] _T_199; // @[Mux.scala 19:72:@47445.4]
  NBufController_10 ctrl ( // @[NBuffers.scala 83:20:@47290.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sEn_2(ctrl_io_sEn_2),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_sDone_2(ctrl_io_sDone_2),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1),
    .io_statesInR_2(ctrl_io_statesInR_2)
  );
  SRAM_71 SRAM ( // @[NBuffers.scala 94:23:@47299.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_rPort_1_en_0(SRAM_io_rPort_1_en_0),
    .io_rPort_1_output_0(SRAM_io_rPort_1_output_0),
    .io_rPort_0_en_0(SRAM_io_rPort_0_en_0),
    .io_rPort_0_output_0(SRAM_io_rPort_0_output_0),
    .io_wPort_0_data_0(SRAM_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_io_wPort_0_en_0)
  );
  SRAM_71 SRAM_1 ( // @[NBuffers.scala 94:23:@47320.4]
    .clock(SRAM_1_clock),
    .reset(SRAM_1_reset),
    .io_rPort_1_en_0(SRAM_1_io_rPort_1_en_0),
    .io_rPort_1_output_0(SRAM_1_io_rPort_1_output_0),
    .io_rPort_0_en_0(SRAM_1_io_rPort_0_en_0),
    .io_rPort_0_output_0(SRAM_1_io_rPort_0_output_0),
    .io_wPort_0_data_0(SRAM_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_1_io_wPort_0_en_0)
  );
  SRAM_71 SRAM_2 ( // @[NBuffers.scala 94:23:@47341.4]
    .clock(SRAM_2_clock),
    .reset(SRAM_2_reset),
    .io_rPort_1_en_0(SRAM_2_io_rPort_1_en_0),
    .io_rPort_1_output_0(SRAM_2_io_rPort_1_output_0),
    .io_rPort_0_en_0(SRAM_2_io_rPort_0_en_0),
    .io_rPort_0_output_0(SRAM_2_io_rPort_0_output_0),
    .io_wPort_0_data_0(SRAM_2_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_2_io_wPort_0_en_0)
  );
  assign _T_140 = ctrl_io_statesInW_0 == 3'h0; // @[NBuffers.scala 104:105:@47362.4]
  assign _T_144 = ctrl_io_statesInR_1 == 3'h0; // @[NBuffers.scala 108:92:@47372.4]
  assign _T_147 = ctrl_io_statesInR_2 == 3'h0; // @[NBuffers.scala 108:92:@47378.4]
  assign _T_150 = ctrl_io_statesInW_0 == 3'h1; // @[NBuffers.scala 104:105:@47384.4]
  assign _T_154 = ctrl_io_statesInR_1 == 3'h1; // @[NBuffers.scala 108:92:@47394.4]
  assign _T_157 = ctrl_io_statesInR_2 == 3'h1; // @[NBuffers.scala 108:92:@47400.4]
  assign _T_160 = ctrl_io_statesInW_0 == 3'h2; // @[NBuffers.scala 104:105:@47406.4]
  assign _T_164 = ctrl_io_statesInR_1 == 3'h2; // @[NBuffers.scala 108:92:@47416.4]
  assign _T_167 = ctrl_io_statesInR_2 == 3'h2; // @[NBuffers.scala 108:92:@47422.4]
  assign _T_177 = _T_144 ? SRAM_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@47431.4]
  assign _T_179 = _T_154 ? SRAM_1_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@47432.4]
  assign _T_181 = _T_164 ? SRAM_2_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@47433.4]
  assign _T_182 = _T_177 | _T_179; // @[Mux.scala 19:72:@47434.4]
  assign _T_194 = _T_147 ? SRAM_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@47442.4]
  assign _T_196 = _T_157 ? SRAM_1_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@47443.4]
  assign _T_198 = _T_167 ? SRAM_2_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@47444.4]
  assign _T_199 = _T_194 | _T_196; // @[Mux.scala 19:72:@47445.4]
  assign io_rPort_1_output_0 = _T_199 | _T_198; // @[NBuffers.scala 115:66:@47449.4]
  assign io_rPort_0_output_0 = _T_182 | _T_181; // @[NBuffers.scala 115:66:@47438.4]
  assign ctrl_clock = clock; // @[:@47291.4]
  assign ctrl_reset = reset; // @[:@47292.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@47293.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@47295.4]
  assign ctrl_io_sEn_2 = io_sEn_2; // @[NBuffers.scala 85:20:@47297.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@47294.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@47296.4]
  assign ctrl_io_sDone_2 = io_sDone_2; // @[NBuffers.scala 86:22:@47298.4]
  assign SRAM_clock = clock; // @[:@47300.4]
  assign SRAM_reset = reset; // @[:@47301.4]
  assign SRAM_io_rPort_1_en_0 = io_rPort_1_en_0 & _T_147; // @[MemPrimitives.scala 43:33:@47382.4]
  assign SRAM_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_144; // @[MemPrimitives.scala 43:33:@47376.4]
  assign SRAM_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@47365.4]
  assign SRAM_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_140; // @[MemPrimitives.scala 37:29:@47371.4]
  assign SRAM_1_clock = clock; // @[:@47321.4]
  assign SRAM_1_reset = reset; // @[:@47322.4]
  assign SRAM_1_io_rPort_1_en_0 = io_rPort_1_en_0 & _T_157; // @[MemPrimitives.scala 43:33:@47404.4]
  assign SRAM_1_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_154; // @[MemPrimitives.scala 43:33:@47398.4]
  assign SRAM_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@47387.4]
  assign SRAM_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_150; // @[MemPrimitives.scala 37:29:@47393.4]
  assign SRAM_2_clock = clock; // @[:@47342.4]
  assign SRAM_2_reset = reset; // @[:@47343.4]
  assign SRAM_2_io_rPort_1_en_0 = io_rPort_1_en_0 & _T_167; // @[MemPrimitives.scala 43:33:@47426.4]
  assign SRAM_2_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_164; // @[MemPrimitives.scala 43:33:@47420.4]
  assign SRAM_2_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@47409.4]
  assign SRAM_2_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_160; // @[MemPrimitives.scala 37:29:@47415.4]
endmodule
module RetimeWrapper_517( // @[:@47489.2]
  input   clock, // @[:@47490.4]
  input   reset, // @[:@47491.4]
  input   io_in, // @[:@47492.4]
  output  io_out // @[:@47492.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@47494.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@47494.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@47494.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@47494.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@47494.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@47494.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@47494.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@47507.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@47506.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@47505.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@47504.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@47503.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@47501.4]
endmodule
module RetimeWrapper_521( // @[:@47617.2]
  input   clock, // @[:@47618.4]
  input   reset, // @[:@47619.4]
  input   io_flow, // @[:@47620.4]
  input   io_in, // @[:@47620.4]
  output  io_out // @[:@47620.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@47622.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@47622.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@47622.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@47622.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@47622.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@47622.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@47622.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@47635.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@47634.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@47633.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@47632.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@47631.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@47629.4]
endmodule
module x593_inr_UnitPipe_sm( // @[:@47637.2]
  input   clock, // @[:@47638.4]
  input   reset, // @[:@47639.4]
  input   io_enable, // @[:@47640.4]
  output  io_done, // @[:@47640.4]
  input   io_ctrDone, // @[:@47640.4]
  output  io_datapathEn, // @[:@47640.4]
  output  io_ctrInc, // @[:@47640.4]
  input   io_parentAck, // @[:@47640.4]
  input   io_backpressure, // @[:@47640.4]
  input   io_break // @[:@47640.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@47642.4]
  wire  active_reset; // @[Controllers.scala 261:22:@47642.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@47642.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@47642.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@47642.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@47642.4]
  wire  done_clock; // @[Controllers.scala 262:20:@47645.4]
  wire  done_reset; // @[Controllers.scala 262:20:@47645.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@47645.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@47645.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@47645.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@47645.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@47679.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@47679.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@47679.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@47679.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@47701.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@47701.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@47701.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@47701.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@47713.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@47713.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@47713.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@47713.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@47713.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@47721.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@47721.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@47721.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@47721.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@47721.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@47737.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@47737.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@47737.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@47737.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@47737.4]
  wire  _T_80; // @[Controllers.scala 264:48:@47650.4]
  wire  _T_81; // @[Controllers.scala 264:46:@47651.4]
  wire  _T_82; // @[Controllers.scala 264:62:@47652.4]
  wire  _T_100; // @[package.scala 100:49:@47670.4]
  reg  _T_103; // @[package.scala 48:56:@47671.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@47694.4]
  wire  _T_124; // @[package.scala 96:25:@47706.4 package.scala 96:25:@47707.4]
  wire  _T_126; // @[package.scala 100:49:@47708.4]
  reg  _T_129; // @[package.scala 48:56:@47709.4]
  reg [31:0] _RAND_1;
  wire  _T_150; // @[package.scala 100:49:@47733.4]
  reg  _T_153; // @[package.scala 48:56:@47734.4]
  reg [31:0] _RAND_2;
  SRFF active ( // @[Controllers.scala 261:22:@47642.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@47645.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_517 RetimeWrapper ( // @[package.scala 93:22:@47679.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_517 RetimeWrapper_1 ( // @[package.scala 93:22:@47701.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@47713.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@47721.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_521 RetimeWrapper_4 ( // @[package.scala 93:22:@47737.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@47650.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@47651.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@47652.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@47670.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@47694.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@47706.4 package.scala 96:25:@47707.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@47708.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@47733.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@47712.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@47697.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@47700.4]
  assign active_clock = clock; // @[:@47643.4]
  assign active_reset = reset; // @[:@47644.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@47655.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@47659.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@47660.4]
  assign done_clock = clock; // @[:@47646.4]
  assign done_reset = reset; // @[:@47647.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@47675.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@47668.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@47669.4]
  assign RetimeWrapper_clock = clock; // @[:@47680.4]
  assign RetimeWrapper_reset = reset; // @[:@47681.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@47682.4]
  assign RetimeWrapper_1_clock = clock; // @[:@47702.4]
  assign RetimeWrapper_1_reset = reset; // @[:@47703.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@47704.4]
  assign RetimeWrapper_2_clock = clock; // @[:@47714.4]
  assign RetimeWrapper_2_reset = reset; // @[:@47715.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@47717.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@47716.4]
  assign RetimeWrapper_3_clock = clock; // @[:@47722.4]
  assign RetimeWrapper_3_reset = reset; // @[:@47723.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@47725.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@47724.4]
  assign RetimeWrapper_4_clock = clock; // @[:@47738.4]
  assign RetimeWrapper_4_reset = reset; // @[:@47739.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@47741.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@47740.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_153 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module RetimeWrapper_526( // @[:@47922.2]
  input          clock, // @[:@47923.4]
  input          reset, // @[:@47924.4]
  input          io_flow, // @[:@47925.4]
  input  [107:0] io_in, // @[:@47925.4]
  output [107:0] io_out // @[:@47925.4]
);
  wire [107:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@47927.4]
  wire [107:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@47927.4]
  wire [107:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@47927.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@47927.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@47927.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@47927.4]
  RetimeShiftRegister #(.WIDTH(108), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@47927.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@47940.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@47939.4]
  assign sr_init = 108'h0; // @[RetimeShiftRegister.scala 19:16:@47938.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@47937.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@47936.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@47934.4]
endmodule
module fix2fixBox_13( // @[:@48006.2]
  input  [53:0] io_a, // @[:@48009.4]
  output [31:0] io_b // @[:@48009.4]
);
  wire [21:0] tmp_frac; // @[Converter.scala 38:42:@48017.4]
  wire [9:0] new_dec; // @[Converter.scala 88:34:@48020.4]
  assign tmp_frac = io_a[43:22]; // @[Converter.scala 38:42:@48017.4]
  assign new_dec = io_a[53:44]; // @[Converter.scala 88:34:@48020.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@48023.4]
endmodule
module x586_mul( // @[:@48025.2]
  input         clock, // @[:@48026.4]
  input         reset, // @[:@48027.4]
  input  [31:0] io_a, // @[:@48028.4]
  input  [31:0] io_b, // @[:@48028.4]
  input         io_flow, // @[:@48028.4]
  output [31:0] io_result // @[:@48028.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@48044.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@48044.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@48044.4]
  wire [107:0] RetimeWrapper_io_in; // @[package.scala 93:22:@48044.4]
  wire [107:0] RetimeWrapper_io_out; // @[package.scala 93:22:@48044.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@48056.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@48056.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@48056.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@48056.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@48056.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@48067.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@48067.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@48067.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@48067.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@48067.4]
  wire [53:0] fix2fixBox_io_a; // @[Math.scala 253:30:@48074.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@48074.4]
  wire  _T_16; // @[FixedPoint.scala 50:25:@48035.4]
  wire [21:0] _T_20; // @[Bitwise.scala 72:12:@48037.4]
  wire [53:0] _T_21; // @[Cat.scala 30:58:@48038.4]
  wire  _T_22; // @[FixedPoint.scala 50:25:@48039.4]
  wire [21:0] _T_26; // @[Bitwise.scala 72:12:@48041.4]
  wire [53:0] _T_27; // @[Cat.scala 30:58:@48042.4]
  wire  _T_34; // @[Math.scala 251:56:@48055.4]
  wire [107:0] _T_30; // @[package.scala 96:25:@48049.4 package.scala 96:25:@48050.4]
  RetimeWrapper_526 RetimeWrapper ( // @[package.scala 93:22:@48044.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_452 RetimeWrapper_1 ( // @[package.scala 93:22:@48056.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_452 RetimeWrapper_2 ( // @[package.scala 93:22:@48067.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  fix2fixBox_13 fix2fixBox ( // @[Math.scala 253:30:@48074.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_16 = io_a[31]; // @[FixedPoint.scala 50:25:@48035.4]
  assign _T_20 = _T_16 ? 22'h3fffff : 22'h0; // @[Bitwise.scala 72:12:@48037.4]
  assign _T_21 = {_T_20,io_a}; // @[Cat.scala 30:58:@48038.4]
  assign _T_22 = io_b[31]; // @[FixedPoint.scala 50:25:@48039.4]
  assign _T_26 = _T_22 ? 22'h3fffff : 22'h0; // @[Bitwise.scala 72:12:@48041.4]
  assign _T_27 = {_T_26,io_b}; // @[Cat.scala 30:58:@48042.4]
  assign _T_34 = _T_16 ^ _T_22; // @[Math.scala 251:56:@48055.4]
  assign _T_30 = RetimeWrapper_io_out; // @[package.scala 96:25:@48049.4 package.scala 96:25:@48050.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@48082.4]
  assign RetimeWrapper_clock = clock; // @[:@48045.4]
  assign RetimeWrapper_reset = reset; // @[:@48046.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@48048.4]
  assign RetimeWrapper_io_in = _T_21 * _T_27; // @[package.scala 94:16:@48047.4]
  assign RetimeWrapper_1_clock = clock; // @[:@48057.4]
  assign RetimeWrapper_1_reset = reset; // @[:@48058.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@48060.4]
  assign RetimeWrapper_1_io_in = _T_16 ^ _T_22; // @[package.scala 94:16:@48059.4]
  assign RetimeWrapper_2_clock = clock; // @[:@48068.4]
  assign RetimeWrapper_2_reset = reset; // @[:@48069.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@48071.4]
  assign RetimeWrapper_2_io_in = _T_34 == 1'h0; // @[package.scala 94:16:@48070.4]
  assign fix2fixBox_io_a = _T_30[53:0]; // @[Math.scala 254:23:@48077.4]
endmodule
module RetimeWrapper_529( // @[:@48096.2]
  input         clock, // @[:@48097.4]
  input         reset, // @[:@48098.4]
  input         io_flow, // @[:@48099.4]
  input  [31:0] io_in, // @[:@48099.4]
  output [31:0] io_out // @[:@48099.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@48101.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@48101.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@48101.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@48101.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@48101.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@48101.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@48101.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@48114.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@48113.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@48112.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@48111.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@48110.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@48108.4]
endmodule
module fix2fixBox_15( // @[:@48410.2]
  input  [32:0] io_a, // @[:@48413.4]
  output [31:0] io_b // @[:@48413.4]
);
  wire [21:0] tmp_frac; // @[Converter.scala 52:23:@48421.4]
  wire [9:0] new_dec; // @[Converter.scala 63:26:@48424.4]
  assign tmp_frac = io_a[21:0]; // @[Converter.scala 52:23:@48421.4]
  assign new_dec = io_a[31:22]; // @[Converter.scala 63:26:@48424.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@48427.4]
endmodule
module add( // @[:@48429.2]
  input  [31:0] io_a, // @[:@48432.4]
  input  [31:0] io_b, // @[:@48432.4]
  output [31:0] io_result // @[:@48432.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@48440.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@48440.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@48447.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@48447.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@48465.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@48465.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@48445.4 Math.scala 724:14:@48446.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@48452.4 Math.scala 724:14:@48453.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@48454.4]
  __37 _ ( // @[Math.scala 720:24:@48440.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __37 __1 ( // @[Math.scala 720:24:@48447.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_15 fix2fixBox ( // @[Math.scala 141:30:@48465.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@48445.4 Math.scala 724:14:@48446.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@48452.4 Math.scala 724:14:@48453.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@48454.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@48473.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@48443.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@48450.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@48468.4]
endmodule
module x748( // @[:@48475.2]
  input         clock, // @[:@48476.4]
  input         reset, // @[:@48477.4]
  input  [31:0] io_m0, // @[:@48478.4]
  input  [31:0] io_m1, // @[:@48478.4]
  input  [31:0] io_add, // @[:@48478.4]
  output [31:0] io_result // @[:@48478.4]
);
  wire  fmamul_x748_clock; // @[Math.scala 262:24:@48486.4]
  wire  fmamul_x748_reset; // @[Math.scala 262:24:@48486.4]
  wire [31:0] fmamul_x748_io_a; // @[Math.scala 262:24:@48486.4]
  wire [31:0] fmamul_x748_io_b; // @[Math.scala 262:24:@48486.4]
  wire  fmamul_x748_io_flow; // @[Math.scala 262:24:@48486.4]
  wire [31:0] fmamul_x748_io_result; // @[Math.scala 262:24:@48486.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@48494.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@48494.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@48494.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@48494.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@48494.4]
  wire [31:0] add_1_io_a; // @[Math.scala 150:24:@48504.4]
  wire [31:0] add_1_io_b; // @[Math.scala 150:24:@48504.4]
  wire [31:0] add_1_io_result; // @[Math.scala 150:24:@48504.4]
  x586_mul fmamul_x748 ( // @[Math.scala 262:24:@48486.4]
    .clock(fmamul_x748_clock),
    .reset(fmamul_x748_reset),
    .io_a(fmamul_x748_io_a),
    .io_b(fmamul_x748_io_b),
    .io_flow(fmamul_x748_io_flow),
    .io_result(fmamul_x748_io_result)
  );
  RetimeWrapper_529 RetimeWrapper ( // @[package.scala 93:22:@48494.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  add add_1 ( // @[Math.scala 150:24:@48504.4]
    .io_a(add_1_io_a),
    .io_b(add_1_io_b),
    .io_result(add_1_io_result)
  );
  assign io_result = add_1_io_result; // @[Math.scala 857:17:@48512.4]
  assign fmamul_x748_clock = clock; // @[:@48487.4]
  assign fmamul_x748_reset = reset; // @[:@48488.4]
  assign fmamul_x748_io_a = io_m0; // @[Math.scala 263:17:@48489.4]
  assign fmamul_x748_io_b = io_m1; // @[Math.scala 264:17:@48490.4]
  assign fmamul_x748_io_flow = 1'h1; // @[Math.scala 265:20:@48491.4]
  assign RetimeWrapper_clock = clock; // @[:@48495.4]
  assign RetimeWrapper_reset = reset; // @[:@48496.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@48498.4]
  assign RetimeWrapper_io_in = io_add; // @[package.scala 94:16:@48497.4]
  assign add_1_io_a = fmamul_x748_io_result; // @[Math.scala 151:17:@48507.4]
  assign add_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@48508.4]
endmodule
module SimBlackBoxesfix2fixBox_42( // @[:@48514.2]
  input  [31:0] io_a, // @[:@48517.4]
  output [31:0] io_b // @[:@48517.4]
);
  wire [21:0] tmp_frac; // @[SimBlackBoxes.scala 56:25:@48525.4]
  wire [9:0] new_dec; // @[SimBlackBoxes.scala 92:36:@48528.4]
  assign tmp_frac = io_a[21:0]; // @[SimBlackBoxes.scala 56:25:@48525.4]
  assign new_dec = io_a[31:22]; // @[SimBlackBoxes.scala 92:36:@48528.4]
  assign io_b = {new_dec,tmp_frac}; // @[SimBlackBoxes.scala 98:40:@48531.4]
endmodule
module cast_x748( // @[:@48533.2]
  input  [31:0] io_b, // @[:@48536.4]
  output [31:0] io_result // @[:@48536.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@48541.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@48541.4]
  SimBlackBoxesfix2fixBox_42 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@48541.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 717:17:@48554.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@48549.4]
endmodule
module RetimeWrapper_534( // @[:@48568.2]
  input         clock, // @[:@48569.4]
  input         reset, // @[:@48570.4]
  input  [31:0] io_in, // @[:@48571.4]
  output [31:0] io_out // @[:@48571.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@48573.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@48573.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@48573.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@48573.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@48573.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@48573.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(12)) sr ( // @[RetimeShiftRegister.scala 15:20:@48573.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@48586.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@48585.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@48584.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@48583.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@48582.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@48580.4]
endmodule
module x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1( // @[:@49252.2]
  input         clock, // @[:@49253.4]
  input         reset, // @[:@49254.4]
  output        io_in_x555_tmp_1_rPort_0_en_0, // @[:@49255.4]
  input  [31:0] io_in_x555_tmp_1_rPort_0_output_0, // @[:@49255.4]
  output        io_in_x555_tmp_1_sEn_1, // @[:@49255.4]
  output        io_in_x555_tmp_1_sDone_1, // @[:@49255.4]
  output        io_in_x554_tmp_0_rPort_0_en_0, // @[:@49255.4]
  input  [31:0] io_in_x554_tmp_0_rPort_0_output_0, // @[:@49255.4]
  output        io_in_x554_tmp_0_sEn_1, // @[:@49255.4]
  output        io_in_x554_tmp_0_sDone_1, // @[:@49255.4]
  output        io_in_x558_tmp_4_sEn_1, // @[:@49255.4]
  output        io_in_x558_tmp_4_sDone_1, // @[:@49255.4]
  output        io_in_x557_tmp_3_sEn_1, // @[:@49255.4]
  output        io_in_x557_tmp_3_sDone_1, // @[:@49255.4]
  output [31:0] io_in_x580_r_0_wPort_0_data_0, // @[:@49255.4]
  output        io_in_x580_r_0_wPort_0_en_0, // @[:@49255.4]
  output        io_in_x580_r_0_sEn_0, // @[:@49255.4]
  output        io_in_x580_r_0_sDone_0, // @[:@49255.4]
  output        io_in_x556_tmp_2_rPort_0_en_0, // @[:@49255.4]
  input  [31:0] io_in_x556_tmp_2_rPort_0_output_0, // @[:@49255.4]
  output        io_in_x556_tmp_2_sEn_1, // @[:@49255.4]
  output        io_in_x556_tmp_2_sDone_1, // @[:@49255.4]
  output [63:0] io_in_instrctrs_9_cycs, // @[:@49255.4]
  output [63:0] io_in_instrctrs_9_iters, // @[:@49255.4]
  input         io_sigsIn_done, // @[:@49255.4]
  input         io_sigsIn_datapathEn, // @[:@49255.4]
  input         io_sigsIn_baseEn, // @[:@49255.4]
  input         io_sigsIn_break, // @[:@49255.4]
  input         io_rr // @[:@49255.4]
);
  wire  cycles_x593_inr_UnitPipe_clock; // @[sm_x593_inr_UnitPipe.scala 87:44:@49613.4]
  wire  cycles_x593_inr_UnitPipe_reset; // @[sm_x593_inr_UnitPipe.scala 87:44:@49613.4]
  wire  cycles_x593_inr_UnitPipe_io_enable; // @[sm_x593_inr_UnitPipe.scala 87:44:@49613.4]
  wire [63:0] cycles_x593_inr_UnitPipe_io_count; // @[sm_x593_inr_UnitPipe.scala 87:44:@49613.4]
  wire  iters_x593_inr_UnitPipe_clock; // @[sm_x593_inr_UnitPipe.scala 88:43:@49616.4]
  wire  iters_x593_inr_UnitPipe_reset; // @[sm_x593_inr_UnitPipe.scala 88:43:@49616.4]
  wire  iters_x593_inr_UnitPipe_io_enable; // @[sm_x593_inr_UnitPipe.scala 88:43:@49616.4]
  wire [63:0] iters_x593_inr_UnitPipe_io_count; // @[sm_x593_inr_UnitPipe.scala 88:43:@49616.4]
  wire  x586_mul_1_clock; // @[Math.scala 262:24:@49674.4]
  wire  x586_mul_1_reset; // @[Math.scala 262:24:@49674.4]
  wire [31:0] x586_mul_1_io_a; // @[Math.scala 262:24:@49674.4]
  wire [31:0] x586_mul_1_io_b; // @[Math.scala 262:24:@49674.4]
  wire  x586_mul_1_io_flow; // @[Math.scala 262:24:@49674.4]
  wire [31:0] x586_mul_1_io_result; // @[Math.scala 262:24:@49674.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@49685.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@49685.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@49685.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@49685.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@49685.4]
  wire  x748_1_clock; // @[Math.scala 860:24:@49694.4]
  wire  x748_1_reset; // @[Math.scala 860:24:@49694.4]
  wire [31:0] x748_1_io_m0; // @[Math.scala 860:24:@49694.4]
  wire [31:0] x748_1_io_m1; // @[Math.scala 860:24:@49694.4]
  wire [31:0] x748_1_io_add; // @[Math.scala 860:24:@49694.4]
  wire [31:0] x748_1_io_result; // @[Math.scala 860:24:@49694.4]
  wire [31:0] cast_x748_io_b; // @[Math.scala 720:24:@49703.4]
  wire [31:0] cast_x748_io_result; // @[Math.scala 720:24:@49703.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@49735.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@49735.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@49735.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@49735.4]
  wire  x749_1_clock; // @[Math.scala 860:24:@49744.4]
  wire  x749_1_reset; // @[Math.scala 860:24:@49744.4]
  wire [31:0] x749_1_io_m0; // @[Math.scala 860:24:@49744.4]
  wire [31:0] x749_1_io_m1; // @[Math.scala 860:24:@49744.4]
  wire [31:0] x749_1_io_add; // @[Math.scala 860:24:@49744.4]
  wire [31:0] x749_1_io_result; // @[Math.scala 860:24:@49744.4]
  wire [31:0] cast_x749_io_b; // @[Math.scala 720:24:@49753.4]
  wire [31:0] cast_x749_io_result; // @[Math.scala 720:24:@49753.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@49769.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@49769.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@49769.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@49769.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@49769.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@49788.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@49788.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@49788.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@49788.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@49788.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@49799.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@49799.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@49799.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@49799.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@49799.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@49810.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@49810.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@49810.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@49810.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@49810.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@49821.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@49821.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@49821.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@49821.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@49821.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@49832.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@49832.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@49832.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@49832.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@49832.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@49843.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@49843.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@49843.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@49843.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@49843.4]
  wire  _T_1828; // @[package.scala 100:49:@49620.4]
  reg  _T_1831; // @[package.scala 48:56:@49621.4]
  reg [31:0] _RAND_0;
  wire  _T_1853; // @[sm_x593_inr_UnitPipe.scala 96:114:@49636.4]
  wire  _T_1854; // @[sm_x593_inr_UnitPipe.scala 96:111:@49637.4]
  wire  _T_1859; // @[implicits.scala 56:10:@49640.4]
  wire  _T_1964; // @[package.scala 96:25:@49774.4 package.scala 96:25:@49775.4]
  wire  _T_1966; // @[implicits.scala 56:10:@49776.4]
  wire  _T_1967; // @[sm_x593_inr_UnitPipe.scala 133:113:@49777.4]
  wire  _T_1976; // @[package.scala 96:25:@49793.4 package.scala 96:25:@49794.4]
  wire  _T_1982; // @[package.scala 96:25:@49804.4 package.scala 96:25:@49805.4]
  wire  _T_1988; // @[package.scala 96:25:@49815.4 package.scala 96:25:@49816.4]
  wire  _T_1994; // @[package.scala 96:25:@49826.4 package.scala 96:25:@49827.4]
  wire  _T_2000; // @[package.scala 96:25:@49837.4 package.scala 96:25:@49838.4]
  wire  _T_2006; // @[package.scala 96:25:@49848.4 package.scala 96:25:@49849.4]
  InstrumentationCounter cycles_x593_inr_UnitPipe ( // @[sm_x593_inr_UnitPipe.scala 87:44:@49613.4]
    .clock(cycles_x593_inr_UnitPipe_clock),
    .reset(cycles_x593_inr_UnitPipe_reset),
    .io_enable(cycles_x593_inr_UnitPipe_io_enable),
    .io_count(cycles_x593_inr_UnitPipe_io_count)
  );
  InstrumentationCounter iters_x593_inr_UnitPipe ( // @[sm_x593_inr_UnitPipe.scala 88:43:@49616.4]
    .clock(iters_x593_inr_UnitPipe_clock),
    .reset(iters_x593_inr_UnitPipe_reset),
    .io_enable(iters_x593_inr_UnitPipe_io_enable),
    .io_count(iters_x593_inr_UnitPipe_io_count)
  );
  x586_mul x586_mul_1 ( // @[Math.scala 262:24:@49674.4]
    .clock(x586_mul_1_clock),
    .reset(x586_mul_1_reset),
    .io_a(x586_mul_1_io_a),
    .io_b(x586_mul_1_io_b),
    .io_flow(x586_mul_1_io_flow),
    .io_result(x586_mul_1_io_result)
  );
  RetimeWrapper_529 RetimeWrapper ( // @[package.scala 93:22:@49685.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x748 x748_1 ( // @[Math.scala 860:24:@49694.4]
    .clock(x748_1_clock),
    .reset(x748_1_reset),
    .io_m0(x748_1_io_m0),
    .io_m1(x748_1_io_m1),
    .io_add(x748_1_io_add),
    .io_result(x748_1_io_result)
  );
  cast_x748 cast_x748 ( // @[Math.scala 720:24:@49703.4]
    .io_b(cast_x748_io_b),
    .io_result(cast_x748_io_result)
  );
  RetimeWrapper_534 RetimeWrapper_1 ( // @[package.scala 93:22:@49735.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x748 x749_1 ( // @[Math.scala 860:24:@49744.4]
    .clock(x749_1_clock),
    .reset(x749_1_reset),
    .io_m0(x749_1_io_m0),
    .io_m1(x749_1_io_m1),
    .io_add(x749_1_io_add),
    .io_result(x749_1_io_result)
  );
  cast_x748 cast_x749 ( // @[Math.scala 720:24:@49753.4]
    .io_b(cast_x749_io_b),
    .io_result(cast_x749_io_result)
  );
  RetimeWrapper_521 RetimeWrapper_2 ( // @[package.scala 93:22:@49769.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@49788.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@49799.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@49810.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@49821.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@49832.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@49843.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  assign _T_1828 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@49620.4]
  assign _T_1853 = ~ io_sigsIn_break; // @[sm_x593_inr_UnitPipe.scala 96:114:@49636.4]
  assign _T_1854 = io_rr & _T_1853; // @[sm_x593_inr_UnitPipe.scala 96:111:@49637.4]
  assign _T_1859 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 56:10:@49640.4]
  assign _T_1964 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@49774.4 package.scala 96:25:@49775.4]
  assign _T_1966 = io_rr ? _T_1964 : 1'h0; // @[implicits.scala 56:10:@49776.4]
  assign _T_1967 = _T_1853 & _T_1966; // @[sm_x593_inr_UnitPipe.scala 133:113:@49777.4]
  assign _T_1976 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@49793.4 package.scala 96:25:@49794.4]
  assign _T_1982 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@49804.4 package.scala 96:25:@49805.4]
  assign _T_1988 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@49815.4 package.scala 96:25:@49816.4]
  assign _T_1994 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@49826.4 package.scala 96:25:@49827.4]
  assign _T_2000 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@49837.4 package.scala 96:25:@49838.4]
  assign _T_2006 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@49848.4 package.scala 96:25:@49849.4]
  assign io_in_x555_tmp_1_rPort_0_en_0 = _T_1854 & _T_1859; // @[MemInterfaceType.scala 110:79:@49669.4]
  assign io_in_x555_tmp_1_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@49807.4]
  assign io_in_x555_tmp_1_sDone_1 = io_rr ? _T_1982 : 1'h0; // @[MemInterfaceType.scala 197:17:@49808.4]
  assign io_in_x554_tmp_0_rPort_0_en_0 = _T_1854 & _T_1859; // @[MemInterfaceType.scala 110:79:@49647.4]
  assign io_in_x554_tmp_0_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@49796.4]
  assign io_in_x554_tmp_0_sDone_1 = io_rr ? _T_1976 : 1'h0; // @[MemInterfaceType.scala 197:17:@49797.4]
  assign io_in_x558_tmp_4_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@49840.4]
  assign io_in_x558_tmp_4_sDone_1 = io_rr ? _T_2000 : 1'h0; // @[MemInterfaceType.scala 197:17:@49841.4]
  assign io_in_x557_tmp_3_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@49829.4]
  assign io_in_x557_tmp_3_sDone_1 = io_rr ? _T_1994 : 1'h0; // @[MemInterfaceType.scala 197:17:@49830.4]
  assign io_in_x580_r_0_wPort_0_data_0 = cast_x749_io_result; // @[MemInterfaceType.scala 90:56:@49784.4]
  assign io_in_x580_r_0_wPort_0_en_0 = _T_1967 & _T_1853; // @[MemInterfaceType.scala 93:57:@49786.4]
  assign io_in_x580_r_0_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@49851.4]
  assign io_in_x580_r_0_sDone_0 = io_rr ? _T_2006 : 1'h0; // @[MemInterfaceType.scala 197:17:@49852.4]
  assign io_in_x556_tmp_2_rPort_0_en_0 = _T_1854 & _T_1859; // @[MemInterfaceType.scala 110:79:@49729.4]
  assign io_in_x556_tmp_2_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@49818.4]
  assign io_in_x556_tmp_2_sDone_1 = io_rr ? _T_1988 : 1'h0; // @[MemInterfaceType.scala 197:17:@49819.4]
  assign io_in_instrctrs_9_cycs = cycles_x593_inr_UnitPipe_io_count; // @[Ledger.scala 293:21:@49625.4]
  assign io_in_instrctrs_9_iters = iters_x593_inr_UnitPipe_io_count; // @[Ledger.scala 294:22:@49626.4]
  assign cycles_x593_inr_UnitPipe_clock = clock; // @[:@49614.4]
  assign cycles_x593_inr_UnitPipe_reset = reset; // @[:@49615.4]
  assign cycles_x593_inr_UnitPipe_io_enable = io_sigsIn_baseEn; // @[sm_x593_inr_UnitPipe.scala 89:42:@49619.4]
  assign iters_x593_inr_UnitPipe_clock = clock; // @[:@49617.4]
  assign iters_x593_inr_UnitPipe_reset = reset; // @[:@49618.4]
  assign iters_x593_inr_UnitPipe_io_enable = io_sigsIn_done & _T_1831; // @[sm_x593_inr_UnitPipe.scala 90:41:@49624.4]
  assign x586_mul_1_clock = clock; // @[:@49675.4]
  assign x586_mul_1_reset = reset; // @[:@49676.4]
  assign x586_mul_1_io_a = io_in_x555_tmp_1_rPort_0_output_0; // @[Math.scala 263:17:@49677.4]
  assign x586_mul_1_io_b = io_in_x555_tmp_1_rPort_0_output_0; // @[Math.scala 264:17:@49678.4]
  assign x586_mul_1_io_flow = 1'h1; // @[Math.scala 265:20:@49679.4]
  assign RetimeWrapper_clock = clock; // @[:@49686.4]
  assign RetimeWrapper_reset = reset; // @[:@49687.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@49689.4]
  assign RetimeWrapper_io_in = io_in_x554_tmp_0_rPort_0_output_0; // @[package.scala 94:16:@49688.4]
  assign x748_1_clock = clock; // @[:@49695.4]
  assign x748_1_reset = reset; // @[:@49696.4]
  assign x748_1_io_m0 = RetimeWrapper_io_out; // @[Math.scala 861:18:@49697.4]
  assign x748_1_io_m1 = RetimeWrapper_io_out; // @[Math.scala 862:18:@49698.4]
  assign x748_1_io_add = x586_mul_1_io_result; // @[Math.scala 863:19:@49699.4]
  assign cast_x748_io_b = x748_1_io_result; // @[Math.scala 721:17:@49706.4]
  assign RetimeWrapper_1_clock = clock; // @[:@49736.4]
  assign RetimeWrapper_1_reset = reset; // @[:@49737.4]
  assign RetimeWrapper_1_io_in = io_in_x556_tmp_2_rPort_0_output_0; // @[package.scala 94:16:@49738.4]
  assign x749_1_clock = clock; // @[:@49745.4]
  assign x749_1_reset = reset; // @[:@49746.4]
  assign x749_1_io_m0 = RetimeWrapper_1_io_out; // @[Math.scala 861:18:@49747.4]
  assign x749_1_io_m1 = RetimeWrapper_1_io_out; // @[Math.scala 862:18:@49748.4]
  assign x749_1_io_add = cast_x748_io_result; // @[Math.scala 863:19:@49749.4]
  assign cast_x749_io_b = x749_1_io_result; // @[Math.scala 721:17:@49756.4]
  assign RetimeWrapper_2_clock = clock; // @[:@49770.4]
  assign RetimeWrapper_2_reset = reset; // @[:@49771.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@49773.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@49772.4]
  assign RetimeWrapper_3_clock = clock; // @[:@49789.4]
  assign RetimeWrapper_3_reset = reset; // @[:@49790.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@49792.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_done; // @[package.scala 94:16:@49791.4]
  assign RetimeWrapper_4_clock = clock; // @[:@49800.4]
  assign RetimeWrapper_4_reset = reset; // @[:@49801.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@49803.4]
  assign RetimeWrapper_4_io_in = io_sigsIn_done; // @[package.scala 94:16:@49802.4]
  assign RetimeWrapper_5_clock = clock; // @[:@49811.4]
  assign RetimeWrapper_5_reset = reset; // @[:@49812.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@49814.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_done; // @[package.scala 94:16:@49813.4]
  assign RetimeWrapper_6_clock = clock; // @[:@49822.4]
  assign RetimeWrapper_6_reset = reset; // @[:@49823.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@49825.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_done; // @[package.scala 94:16:@49824.4]
  assign RetimeWrapper_7_clock = clock; // @[:@49833.4]
  assign RetimeWrapper_7_reset = reset; // @[:@49834.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@49836.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_done; // @[package.scala 94:16:@49835.4]
  assign RetimeWrapper_8_clock = clock; // @[:@49844.4]
  assign RetimeWrapper_8_reset = reset; // @[:@49845.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@49847.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_done; // @[package.scala 94:16:@49846.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1831 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1831 <= 1'h0;
    end else begin
      _T_1831 <= _T_1828;
    end
  end
endmodule
module SRAM_74( // @[:@50679.2]
  input         clock, // @[:@50680.4]
  input         reset, // @[:@50681.4]
  input         io_rPort_0_en_0, // @[:@50682.4]
  output [31:0] io_rPort_0_output_0, // @[:@50682.4]
  input  [31:0] io_wPort_0_data_0, // @[:@50682.4]
  input         io_wPort_0_en_0 // @[:@50682.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@50697.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@50697.4]
  wire  Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@50697.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@50697.4]
  wire  Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@50697.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@50697.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@50697.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@50697.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@50723.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@50723.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@50737.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@50737.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@50737.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@50737.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@50737.4]
  wire [33:0] _T_70; // @[Cat.scala 30:58:@50715.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@50727.4]
  wire [2:0] _T_78; // @[Cat.scala 30:58:@50729.4]
  Mem1D_39 Mem1D ( // @[MemPrimitives.scala 64:21:@50697.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@50723.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@50737.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_70 = {io_wPort_0_en_0,io_wPort_0_data_0,1'h0}; // @[Cat.scala 30:58:@50715.4]
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@50727.4]
  assign _T_78 = {_T_76,1'h1,1'h0}; // @[Cat.scala 30:58:@50729.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@50744.4]
  assign Mem1D_clock = clock; // @[:@50698.4]
  assign Mem1D_reset = reset; // @[:@50699.4]
  assign Mem1D_io_r_ofs_0 = _T_78[0]; // @[MemPrimitives.scala 131:28:@50733.4]
  assign Mem1D_io_r_backpressure = _T_78[1]; // @[MemPrimitives.scala 132:32:@50734.4]
  assign Mem1D_io_w_ofs_0 = _T_70[0]; // @[MemPrimitives.scala 94:28:@50719.4]
  assign Mem1D_io_w_data_0 = _T_70[32:1]; // @[MemPrimitives.scala 95:29:@50720.4]
  assign Mem1D_io_w_en_0 = _T_70[33]; // @[MemPrimitives.scala 96:27:@50721.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@50726.4]
  assign RetimeWrapper_clock = clock; // @[:@50738.4]
  assign RetimeWrapper_reset = reset; // @[:@50739.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@50741.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@50740.4]
endmodule
module x594_force_0( // @[:@50947.2]
  input         clock, // @[:@50948.4]
  input         reset, // @[:@50949.4]
  input         io_rPort_0_en_0, // @[:@50950.4]
  output [31:0] io_rPort_0_output_0, // @[:@50950.4]
  input  [31:0] io_wPort_0_data_0, // @[:@50950.4]
  input         io_wPort_0_en_0, // @[:@50950.4]
  input         io_sEn_0, // @[:@50950.4]
  input         io_sEn_1, // @[:@50950.4]
  input         io_sDone_0, // @[:@50950.4]
  input         io_sDone_1 // @[:@50950.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@50959.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@50959.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@50959.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@50959.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@50959.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@50959.4]
  wire [2:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@50959.4]
  wire [2:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@50959.4]
  wire  SRAM_clock; // @[NBuffers.scala 94:23:@50966.4]
  wire  SRAM_reset; // @[NBuffers.scala 94:23:@50966.4]
  wire  SRAM_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@50966.4]
  wire [31:0] SRAM_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@50966.4]
  wire [31:0] SRAM_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@50966.4]
  wire  SRAM_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@50966.4]
  wire  SRAM_1_clock; // @[NBuffers.scala 94:23:@50982.4]
  wire  SRAM_1_reset; // @[NBuffers.scala 94:23:@50982.4]
  wire  SRAM_1_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@50982.4]
  wire [31:0] SRAM_1_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@50982.4]
  wire [31:0] SRAM_1_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@50982.4]
  wire  SRAM_1_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@50982.4]
  wire  _T_110; // @[NBuffers.scala 104:105:@50998.4]
  wire  _T_114; // @[NBuffers.scala 108:92:@51008.4]
  wire  _T_117; // @[NBuffers.scala 104:105:@51014.4]
  wire  _T_121; // @[NBuffers.scala 108:92:@51024.4]
  wire [31:0] _T_129; // @[Mux.scala 19:72:@51032.4]
  wire [31:0] _T_131; // @[Mux.scala 19:72:@51033.4]
  NBufController ctrl ( // @[NBuffers.scala 83:20:@50959.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1)
  );
  SRAM_74 SRAM ( // @[NBuffers.scala 94:23:@50966.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_rPort_0_en_0(SRAM_io_rPort_0_en_0),
    .io_rPort_0_output_0(SRAM_io_rPort_0_output_0),
    .io_wPort_0_data_0(SRAM_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_io_wPort_0_en_0)
  );
  SRAM_74 SRAM_1 ( // @[NBuffers.scala 94:23:@50982.4]
    .clock(SRAM_1_clock),
    .reset(SRAM_1_reset),
    .io_rPort_0_en_0(SRAM_1_io_rPort_0_en_0),
    .io_rPort_0_output_0(SRAM_1_io_rPort_0_output_0),
    .io_wPort_0_data_0(SRAM_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_1_io_wPort_0_en_0)
  );
  assign _T_110 = ctrl_io_statesInW_0 == 3'h0; // @[NBuffers.scala 104:105:@50998.4]
  assign _T_114 = ctrl_io_statesInR_1 == 3'h0; // @[NBuffers.scala 108:92:@51008.4]
  assign _T_117 = ctrl_io_statesInW_0 == 3'h1; // @[NBuffers.scala 104:105:@51014.4]
  assign _T_121 = ctrl_io_statesInR_1 == 3'h1; // @[NBuffers.scala 108:92:@51024.4]
  assign _T_129 = _T_114 ? SRAM_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@51032.4]
  assign _T_131 = _T_121 ? SRAM_1_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@51033.4]
  assign io_rPort_0_output_0 = _T_129 | _T_131; // @[NBuffers.scala 115:66:@51037.4]
  assign ctrl_clock = clock; // @[:@50960.4]
  assign ctrl_reset = reset; // @[:@50961.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@50962.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@50964.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@50963.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@50965.4]
  assign SRAM_clock = clock; // @[:@50967.4]
  assign SRAM_reset = reset; // @[:@50968.4]
  assign SRAM_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_114; // @[MemPrimitives.scala 43:33:@51012.4]
  assign SRAM_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@51001.4]
  assign SRAM_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_110; // @[MemPrimitives.scala 37:29:@51007.4]
  assign SRAM_1_clock = clock; // @[:@50983.4]
  assign SRAM_1_reset = reset; // @[:@50984.4]
  assign SRAM_1_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_121; // @[MemPrimitives.scala 43:33:@51028.4]
  assign SRAM_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@51017.4]
  assign SRAM_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_117; // @[MemPrimitives.scala 37:29:@51023.4]
endmodule
module FF_28( // @[:@51730.2]
  input   clock, // @[:@51731.4]
  input   reset, // @[:@51732.4]
  output  io_rPort_1_output_0, // @[:@51733.4]
  output  io_rPort_0_output_0, // @[:@51733.4]
  input   io_wPort_0_data_0, // @[:@51733.4]
  input   io_wPort_0_reset, // @[:@51733.4]
  input   io_wPort_0_en_0 // @[:@51733.4]
);
  reg  ff; // @[MemPrimitives.scala 321:19:@51753.4]
  reg [31:0] _RAND_0;
  wire  _T_94; // @[MemPrimitives.scala 325:32:@51755.4]
  wire  _T_95; // @[MemPrimitives.scala 325:12:@51756.4]
  assign _T_94 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@51755.4]
  assign _T_95 = io_wPort_0_reset ? 1'h0 : _T_94; // @[MemPrimitives.scala 325:12:@51756.4]
  assign io_rPort_1_output_0 = ff; // @[MemPrimitives.scala 326:34:@51759.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@51758.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 1'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 1'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module x595_reg( // @[:@51792.2]
  input   clock, // @[:@51793.4]
  input   reset, // @[:@51794.4]
  output  io_rPort_1_output_0, // @[:@51795.4]
  output  io_rPort_0_output_0, // @[:@51795.4]
  input   io_wPort_0_data_0, // @[:@51795.4]
  input   io_wPort_0_reset, // @[:@51795.4]
  input   io_wPort_0_en_0, // @[:@51795.4]
  input   io_sEn_0, // @[:@51795.4]
  input   io_sEn_1, // @[:@51795.4]
  input   io_sDone_0, // @[:@51795.4]
  input   io_sDone_1 // @[:@51795.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@51805.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@51805.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@51805.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@51805.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@51805.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@51805.4]
  wire [2:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@51805.4]
  wire [2:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@51805.4]
  wire  FF_clock; // @[NBuffers.scala 146:23:@51812.4]
  wire  FF_reset; // @[NBuffers.scala 146:23:@51812.4]
  wire  FF_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@51812.4]
  wire  FF_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@51812.4]
  wire  FF_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@51812.4]
  wire  FF_io_wPort_0_reset; // @[NBuffers.scala 146:23:@51812.4]
  wire  FF_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@51812.4]
  wire  FF_1_clock; // @[NBuffers.scala 146:23:@51833.4]
  wire  FF_1_reset; // @[NBuffers.scala 146:23:@51833.4]
  wire  FF_1_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@51833.4]
  wire  FF_1_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@51833.4]
  wire  FF_1_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@51833.4]
  wire  FF_1_io_wPort_0_reset; // @[NBuffers.scala 146:23:@51833.4]
  wire  FF_1_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@51833.4]
  wire  _T_140; // @[NBuffers.scala 153:105:@51856.4]
  wire  _T_144; // @[NBuffers.scala 157:92:@51866.4]
  wire  _T_150; // @[NBuffers.scala 153:105:@51878.4]
  wire  _T_154; // @[NBuffers.scala 157:92:@51888.4]
  wire  _T_165; // @[Mux.scala 19:72:@51902.4]
  wire  _T_167; // @[Mux.scala 19:72:@51903.4]
  wire  _T_177; // @[Mux.scala 19:72:@51910.4]
  wire  _T_179; // @[Mux.scala 19:72:@51911.4]
  NBufController ctrl ( // @[NBuffers.scala 83:20:@51805.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1)
  );
  FF_28 FF ( // @[NBuffers.scala 146:23:@51812.4]
    .clock(FF_clock),
    .reset(FF_reset),
    .io_rPort_1_output_0(FF_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_io_wPort_0_en_0)
  );
  FF_28 FF_1 ( // @[NBuffers.scala 146:23:@51833.4]
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_rPort_1_output_0(FF_1_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_1_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_1_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_1_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_1_io_wPort_0_en_0)
  );
  assign _T_140 = ctrl_io_statesInW_0 == 3'h0; // @[NBuffers.scala 153:105:@51856.4]
  assign _T_144 = ctrl_io_statesInR_1 == 3'h0; // @[NBuffers.scala 157:92:@51866.4]
  assign _T_150 = ctrl_io_statesInW_0 == 3'h1; // @[NBuffers.scala 153:105:@51878.4]
  assign _T_154 = ctrl_io_statesInR_1 == 3'h1; // @[NBuffers.scala 157:92:@51888.4]
  assign _T_165 = _T_144 ? FF_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@51902.4]
  assign _T_167 = _T_154 ? FF_1_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@51903.4]
  assign _T_177 = _T_144 ? FF_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@51910.4]
  assign _T_179 = _T_154 ? FF_1_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@51911.4]
  assign io_rPort_1_output_0 = _T_177 | _T_179; // @[NBuffers.scala 163:66:@51915.4]
  assign io_rPort_0_output_0 = _T_165 | _T_167; // @[NBuffers.scala 163:66:@51907.4]
  assign ctrl_clock = clock; // @[:@51806.4]
  assign ctrl_reset = reset; // @[:@51807.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@51808.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@51810.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@51809.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@51811.4]
  assign FF_clock = clock; // @[:@51813.4]
  assign FF_reset = reset; // @[:@51814.4]
  assign FF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@51859.4]
  assign FF_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@51860.4]
  assign FF_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_140; // @[MemPrimitives.scala 37:29:@51865.4]
  assign FF_1_clock = clock; // @[:@51834.4]
  assign FF_1_reset = reset; // @[:@51835.4]
  assign FF_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@51881.4]
  assign FF_1_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@51882.4]
  assign FF_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_150; // @[MemPrimitives.scala 37:29:@51887.4]
endmodule
module FF_30( // @[:@52608.2]
  input   clock, // @[:@52609.4]
  input   reset, // @[:@52610.4]
  output  io_rPort_0_output_0, // @[:@52611.4]
  input   io_wPort_0_data_0, // @[:@52611.4]
  input   io_wPort_0_reset, // @[:@52611.4]
  input   io_wPort_0_en_0 // @[:@52611.4]
);
  reg  ff; // @[MemPrimitives.scala 321:19:@52626.4]
  reg [31:0] _RAND_0;
  wire  _T_68; // @[MemPrimitives.scala 325:32:@52628.4]
  wire  _T_69; // @[MemPrimitives.scala 325:12:@52629.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@52628.4]
  assign _T_69 = io_wPort_0_reset ? 1'h0 : _T_68; // @[MemPrimitives.scala 325:12:@52629.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@52631.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 1'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 1'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module x596_reg( // @[:@52658.2]
  input   clock, // @[:@52659.4]
  input   reset, // @[:@52660.4]
  output  io_rPort_0_output_0, // @[:@52661.4]
  input   io_wPort_0_data_0, // @[:@52661.4]
  input   io_wPort_0_reset, // @[:@52661.4]
  input   io_wPort_0_en_0, // @[:@52661.4]
  input   io_sEn_0, // @[:@52661.4]
  input   io_sEn_1, // @[:@52661.4]
  input   io_sDone_0, // @[:@52661.4]
  input   io_sDone_1 // @[:@52661.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@52670.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@52670.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@52670.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@52670.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@52670.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@52670.4]
  wire [2:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@52670.4]
  wire [2:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@52670.4]
  wire  FF_clock; // @[NBuffers.scala 146:23:@52677.4]
  wire  FF_reset; // @[NBuffers.scala 146:23:@52677.4]
  wire  FF_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@52677.4]
  wire  FF_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@52677.4]
  wire  FF_io_wPort_0_reset; // @[NBuffers.scala 146:23:@52677.4]
  wire  FF_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@52677.4]
  wire  FF_1_clock; // @[NBuffers.scala 146:23:@52693.4]
  wire  FF_1_reset; // @[NBuffers.scala 146:23:@52693.4]
  wire  FF_1_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@52693.4]
  wire  FF_1_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@52693.4]
  wire  FF_1_io_wPort_0_reset; // @[NBuffers.scala 146:23:@52693.4]
  wire  FF_1_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@52693.4]
  wire  _T_110; // @[NBuffers.scala 153:105:@52711.4]
  wire  _T_114; // @[NBuffers.scala 157:92:@52721.4]
  wire  _T_117; // @[NBuffers.scala 153:105:@52727.4]
  wire  _T_121; // @[NBuffers.scala 157:92:@52737.4]
  wire  _T_129; // @[Mux.scala 19:72:@52745.4]
  wire  _T_131; // @[Mux.scala 19:72:@52746.4]
  NBufController ctrl ( // @[NBuffers.scala 83:20:@52670.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1)
  );
  FF_30 FF ( // @[NBuffers.scala 146:23:@52677.4]
    .clock(FF_clock),
    .reset(FF_reset),
    .io_rPort_0_output_0(FF_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_io_wPort_0_en_0)
  );
  FF_30 FF_1 ( // @[NBuffers.scala 146:23:@52693.4]
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_rPort_0_output_0(FF_1_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_1_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_1_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_1_io_wPort_0_en_0)
  );
  assign _T_110 = ctrl_io_statesInW_0 == 3'h0; // @[NBuffers.scala 153:105:@52711.4]
  assign _T_114 = ctrl_io_statesInR_1 == 3'h0; // @[NBuffers.scala 157:92:@52721.4]
  assign _T_117 = ctrl_io_statesInW_0 == 3'h1; // @[NBuffers.scala 153:105:@52727.4]
  assign _T_121 = ctrl_io_statesInR_1 == 3'h1; // @[NBuffers.scala 157:92:@52737.4]
  assign _T_129 = _T_114 ? FF_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@52745.4]
  assign _T_131 = _T_121 ? FF_1_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@52746.4]
  assign io_rPort_0_output_0 = _T_129 | _T_131; // @[NBuffers.scala 163:66:@52750.4]
  assign ctrl_clock = clock; // @[:@52671.4]
  assign ctrl_reset = reset; // @[:@52672.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@52673.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@52675.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@52674.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@52676.4]
  assign FF_clock = clock; // @[:@52678.4]
  assign FF_reset = reset; // @[:@52679.4]
  assign FF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@52714.4]
  assign FF_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@52715.4]
  assign FF_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_110; // @[MemPrimitives.scala 37:29:@52720.4]
  assign FF_1_clock = clock; // @[:@52694.4]
  assign FF_1_reset = reset; // @[:@52695.4]
  assign FF_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@52730.4]
  assign FF_1_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@52731.4]
  assign FF_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_117; // @[MemPrimitives.scala 37:29:@52736.4]
endmodule
module x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1( // @[:@53531.2]
  input         clock, // @[:@53532.4]
  input         reset, // @[:@53533.4]
  output        io_in_x555_tmp_1_sEn_2, // @[:@53534.4]
  output        io_in_x555_tmp_1_sDone_2, // @[:@53534.4]
  output        io_in_x554_tmp_0_sEn_2, // @[:@53534.4]
  output        io_in_x554_tmp_0_sDone_2, // @[:@53534.4]
  output        io_in_x558_tmp_4_sEn_2, // @[:@53534.4]
  output        io_in_x558_tmp_4_sDone_2, // @[:@53534.4]
  output        io_in_x557_tmp_3_sEn_2, // @[:@53534.4]
  output        io_in_x557_tmp_3_sDone_2, // @[:@53534.4]
  output        io_in_x580_r_0_rPort_0_en_0, // @[:@53534.4]
  input  [31:0] io_in_x580_r_0_rPort_0_output_0, // @[:@53534.4]
  output        io_in_x580_r_0_sEn_1, // @[:@53534.4]
  output        io_in_x580_r_0_sDone_1, // @[:@53534.4]
  output        io_in_x595_reg_wPort_0_data_0, // @[:@53534.4]
  output        io_in_x595_reg_wPort_0_reset, // @[:@53534.4]
  output        io_in_x595_reg_wPort_0_en_0, // @[:@53534.4]
  output        io_in_x595_reg_reset, // @[:@53534.4]
  output        io_in_x595_reg_sEn_0, // @[:@53534.4]
  output        io_in_x595_reg_sDone_0, // @[:@53534.4]
  output        io_in_x556_tmp_2_sEn_2, // @[:@53534.4]
  output        io_in_x556_tmp_2_sDone_2, // @[:@53534.4]
  output        io_in_x596_reg_wPort_0_data_0, // @[:@53534.4]
  output        io_in_x596_reg_wPort_0_reset, // @[:@53534.4]
  output        io_in_x596_reg_wPort_0_en_0, // @[:@53534.4]
  output        io_in_x596_reg_reset, // @[:@53534.4]
  output        io_in_x596_reg_sEn_0, // @[:@53534.4]
  output        io_in_x596_reg_sDone_0, // @[:@53534.4]
  output [63:0] io_in_instrctrs_10_cycs, // @[:@53534.4]
  output [63:0] io_in_instrctrs_10_iters, // @[:@53534.4]
  input         io_sigsIn_done, // @[:@53534.4]
  input         io_sigsIn_datapathEn, // @[:@53534.4]
  input         io_sigsIn_baseEn, // @[:@53534.4]
  input         io_sigsIn_break, // @[:@53534.4]
  input         io_rr // @[:@53534.4]
);
  wire  cycles_x605_inr_UnitPipe_clock; // @[sm_x605_inr_UnitPipe.scala 95:44:@53951.4]
  wire  cycles_x605_inr_UnitPipe_reset; // @[sm_x605_inr_UnitPipe.scala 95:44:@53951.4]
  wire  cycles_x605_inr_UnitPipe_io_enable; // @[sm_x605_inr_UnitPipe.scala 95:44:@53951.4]
  wire [63:0] cycles_x605_inr_UnitPipe_io_count; // @[sm_x605_inr_UnitPipe.scala 95:44:@53951.4]
  wire  iters_x605_inr_UnitPipe_clock; // @[sm_x605_inr_UnitPipe.scala 96:43:@53954.4]
  wire  iters_x605_inr_UnitPipe_reset; // @[sm_x605_inr_UnitPipe.scala 96:43:@53954.4]
  wire  iters_x605_inr_UnitPipe_io_enable; // @[sm_x605_inr_UnitPipe.scala 96:43:@53954.4]
  wire [63:0] iters_x605_inr_UnitPipe_io_count; // @[sm_x605_inr_UnitPipe.scala 96:43:@53954.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@54013.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@54013.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@54013.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@54013.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@54013.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@54033.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@54033.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@54033.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@54033.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@54033.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@54050.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@54050.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@54050.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@54050.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@54050.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@54061.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@54061.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@54061.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@54061.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@54061.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@54072.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@54072.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@54072.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@54072.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@54072.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@54083.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@54083.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@54083.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@54083.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@54083.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@54094.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@54094.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@54094.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@54094.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@54094.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@54105.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@54105.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@54105.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@54105.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@54105.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@54116.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@54116.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@54116.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@54116.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@54116.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@54127.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@54127.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@54127.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@54127.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@54127.4]
  wire  _T_2308; // @[package.scala 100:49:@53958.4]
  reg  _T_2311; // @[package.scala 48:56:@53959.4]
  reg [31:0] _RAND_0;
  wire  _T_2333; // @[sm_x605_inr_UnitPipe.scala 104:114:@53974.4]
  wire  _T_2334; // @[sm_x605_inr_UnitPipe.scala 104:111:@53975.4]
  wire  _T_2339; // @[implicits.scala 56:10:@53978.4]
  wire [31:0] _T_2351; // @[Math.scala 476:50:@53993.4]
  wire  x599; // @[Math.scala 476:44:@53994.4]
  wire  x600; // @[Math.scala 476:44:@54001.4]
  wire  x601; // @[sm_x605_inr_UnitPipe.scala 114:20:@54004.4]
  wire  _T_2372; // @[package.scala 96:25:@54018.4 package.scala 96:25:@54019.4]
  wire  _T_2374; // @[implicits.scala 56:10:@54020.4]
  wire  _T_2375; // @[sm_x605_inr_UnitPipe.scala 121:133:@54021.4]
  wire  _T_2387; // @[package.scala 96:25:@54038.4 package.scala 96:25:@54039.4]
  wire  _T_2389; // @[implicits.scala 56:10:@54040.4]
  wire  _T_2390; // @[sm_x605_inr_UnitPipe.scala 126:133:@54041.4]
  wire  _T_2399; // @[package.scala 96:25:@54055.4 package.scala 96:25:@54056.4]
  wire  _T_2405; // @[package.scala 96:25:@54066.4 package.scala 96:25:@54067.4]
  wire  _T_2411; // @[package.scala 96:25:@54077.4 package.scala 96:25:@54078.4]
  wire  _T_2417; // @[package.scala 96:25:@54088.4 package.scala 96:25:@54089.4]
  wire  _T_2423; // @[package.scala 96:25:@54099.4 package.scala 96:25:@54100.4]
  wire  _T_2429; // @[package.scala 96:25:@54110.4 package.scala 96:25:@54111.4]
  wire  _T_2435; // @[package.scala 96:25:@54121.4 package.scala 96:25:@54122.4]
  wire  _T_2441; // @[package.scala 96:25:@54132.4 package.scala 96:25:@54133.4]
  InstrumentationCounter cycles_x605_inr_UnitPipe ( // @[sm_x605_inr_UnitPipe.scala 95:44:@53951.4]
    .clock(cycles_x605_inr_UnitPipe_clock),
    .reset(cycles_x605_inr_UnitPipe_reset),
    .io_enable(cycles_x605_inr_UnitPipe_io_enable),
    .io_count(cycles_x605_inr_UnitPipe_io_count)
  );
  InstrumentationCounter iters_x605_inr_UnitPipe ( // @[sm_x605_inr_UnitPipe.scala 96:43:@53954.4]
    .clock(iters_x605_inr_UnitPipe_clock),
    .reset(iters_x605_inr_UnitPipe_reset),
    .io_enable(iters_x605_inr_UnitPipe_io_enable),
    .io_count(iters_x605_inr_UnitPipe_io_count)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@54013.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@54033.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@54050.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@54061.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@54072.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@54083.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@54094.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@54105.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@54116.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@54127.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  assign _T_2308 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@53958.4]
  assign _T_2333 = ~ io_sigsIn_break; // @[sm_x605_inr_UnitPipe.scala 104:114:@53974.4]
  assign _T_2334 = io_rr & _T_2333; // @[sm_x605_inr_UnitPipe.scala 104:111:@53975.4]
  assign _T_2339 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 56:10:@53978.4]
  assign _T_2351 = $signed(io_in_x580_r_0_rPort_0_output_0); // @[Math.scala 476:50:@53993.4]
  assign x599 = $signed(32'sh0) < $signed(_T_2351); // @[Math.scala 476:44:@53994.4]
  assign x600 = $signed(32'sh400000) < $signed(_T_2351); // @[Math.scala 476:44:@54001.4]
  assign x601 = x599 & x600; // @[sm_x605_inr_UnitPipe.scala 114:20:@54004.4]
  assign _T_2372 = RetimeWrapper_io_out; // @[package.scala 96:25:@54018.4 package.scala 96:25:@54019.4]
  assign _T_2374 = io_rr ? _T_2372 : 1'h0; // @[implicits.scala 56:10:@54020.4]
  assign _T_2375 = _T_2333 & _T_2374; // @[sm_x605_inr_UnitPipe.scala 121:133:@54021.4]
  assign _T_2387 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@54038.4 package.scala 96:25:@54039.4]
  assign _T_2389 = io_rr ? _T_2387 : 1'h0; // @[implicits.scala 56:10:@54040.4]
  assign _T_2390 = _T_2333 & _T_2389; // @[sm_x605_inr_UnitPipe.scala 126:133:@54041.4]
  assign _T_2399 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@54055.4 package.scala 96:25:@54056.4]
  assign _T_2405 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@54066.4 package.scala 96:25:@54067.4]
  assign _T_2411 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@54077.4 package.scala 96:25:@54078.4]
  assign _T_2417 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@54088.4 package.scala 96:25:@54089.4]
  assign _T_2423 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@54099.4 package.scala 96:25:@54100.4]
  assign _T_2429 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@54110.4 package.scala 96:25:@54111.4]
  assign _T_2435 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@54121.4 package.scala 96:25:@54122.4]
  assign _T_2441 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@54132.4 package.scala 96:25:@54133.4]
  assign io_in_x555_tmp_1_sEn_2 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@54069.4]
  assign io_in_x555_tmp_1_sDone_2 = io_rr ? _T_2405 : 1'h0; // @[MemInterfaceType.scala 197:17:@54070.4]
  assign io_in_x554_tmp_0_sEn_2 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@54058.4]
  assign io_in_x554_tmp_0_sDone_2 = io_rr ? _T_2399 : 1'h0; // @[MemInterfaceType.scala 197:17:@54059.4]
  assign io_in_x558_tmp_4_sEn_2 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@54102.4]
  assign io_in_x558_tmp_4_sDone_2 = io_rr ? _T_2423 : 1'h0; // @[MemInterfaceType.scala 197:17:@54103.4]
  assign io_in_x557_tmp_3_sEn_2 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@54091.4]
  assign io_in_x557_tmp_3_sDone_2 = io_rr ? _T_2417 : 1'h0; // @[MemInterfaceType.scala 197:17:@54092.4]
  assign io_in_x580_r_0_rPort_0_en_0 = _T_2334 & _T_2339; // @[MemInterfaceType.scala 110:79:@53985.4]
  assign io_in_x580_r_0_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@54113.4]
  assign io_in_x580_r_0_sDone_1 = io_rr ? _T_2429 : 1'h0; // @[MemInterfaceType.scala 197:17:@54114.4]
  assign io_in_x595_reg_wPort_0_data_0 = x599 & x600; // @[MemInterfaceType.scala 90:56:@54026.4]
  assign io_in_x595_reg_wPort_0_reset = io_in_x595_reg_reset; // @[MemInterfaceType.scala 91:23:@54027.4]
  assign io_in_x595_reg_wPort_0_en_0 = _T_2375 & _T_2333; // @[MemInterfaceType.scala 93:57:@54028.4]
  assign io_in_x595_reg_reset = 1'h0;
  assign io_in_x595_reg_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@54124.4]
  assign io_in_x595_reg_sDone_0 = io_rr ? _T_2435 : 1'h0; // @[MemInterfaceType.scala 197:17:@54125.4]
  assign io_in_x556_tmp_2_sEn_2 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@54080.4]
  assign io_in_x556_tmp_2_sDone_2 = io_rr ? _T_2411 : 1'h0; // @[MemInterfaceType.scala 197:17:@54081.4]
  assign io_in_x596_reg_wPort_0_data_0 = ~ x601; // @[MemInterfaceType.scala 90:56:@54046.4]
  assign io_in_x596_reg_wPort_0_reset = io_in_x596_reg_reset; // @[MemInterfaceType.scala 91:23:@54047.4]
  assign io_in_x596_reg_wPort_0_en_0 = _T_2390 & _T_2333; // @[MemInterfaceType.scala 93:57:@54048.4]
  assign io_in_x596_reg_reset = 1'h0;
  assign io_in_x596_reg_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@54135.4]
  assign io_in_x596_reg_sDone_0 = io_rr ? _T_2441 : 1'h0; // @[MemInterfaceType.scala 197:17:@54136.4]
  assign io_in_instrctrs_10_cycs = cycles_x605_inr_UnitPipe_io_count; // @[Ledger.scala 293:21:@53963.4]
  assign io_in_instrctrs_10_iters = iters_x605_inr_UnitPipe_io_count; // @[Ledger.scala 294:22:@53964.4]
  assign cycles_x605_inr_UnitPipe_clock = clock; // @[:@53952.4]
  assign cycles_x605_inr_UnitPipe_reset = reset; // @[:@53953.4]
  assign cycles_x605_inr_UnitPipe_io_enable = io_sigsIn_baseEn; // @[sm_x605_inr_UnitPipe.scala 97:42:@53957.4]
  assign iters_x605_inr_UnitPipe_clock = clock; // @[:@53955.4]
  assign iters_x605_inr_UnitPipe_reset = reset; // @[:@53956.4]
  assign iters_x605_inr_UnitPipe_io_enable = io_sigsIn_done & _T_2311; // @[sm_x605_inr_UnitPipe.scala 98:41:@53962.4]
  assign RetimeWrapper_clock = clock; // @[:@54014.4]
  assign RetimeWrapper_reset = reset; // @[:@54015.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@54017.4]
  assign RetimeWrapper_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@54016.4]
  assign RetimeWrapper_1_clock = clock; // @[:@54034.4]
  assign RetimeWrapper_1_reset = reset; // @[:@54035.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@54037.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@54036.4]
  assign RetimeWrapper_2_clock = clock; // @[:@54051.4]
  assign RetimeWrapper_2_reset = reset; // @[:@54052.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@54054.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_done; // @[package.scala 94:16:@54053.4]
  assign RetimeWrapper_3_clock = clock; // @[:@54062.4]
  assign RetimeWrapper_3_reset = reset; // @[:@54063.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@54065.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_done; // @[package.scala 94:16:@54064.4]
  assign RetimeWrapper_4_clock = clock; // @[:@54073.4]
  assign RetimeWrapper_4_reset = reset; // @[:@54074.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@54076.4]
  assign RetimeWrapper_4_io_in = io_sigsIn_done; // @[package.scala 94:16:@54075.4]
  assign RetimeWrapper_5_clock = clock; // @[:@54084.4]
  assign RetimeWrapper_5_reset = reset; // @[:@54085.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@54087.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_done; // @[package.scala 94:16:@54086.4]
  assign RetimeWrapper_6_clock = clock; // @[:@54095.4]
  assign RetimeWrapper_6_reset = reset; // @[:@54096.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@54098.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_done; // @[package.scala 94:16:@54097.4]
  assign RetimeWrapper_7_clock = clock; // @[:@54106.4]
  assign RetimeWrapper_7_reset = reset; // @[:@54107.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@54109.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_done; // @[package.scala 94:16:@54108.4]
  assign RetimeWrapper_8_clock = clock; // @[:@54117.4]
  assign RetimeWrapper_8_reset = reset; // @[:@54118.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@54120.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_done; // @[package.scala 94:16:@54119.4]
  assign RetimeWrapper_9_clock = clock; // @[:@54128.4]
  assign RetimeWrapper_9_reset = reset; // @[:@54129.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@54131.4]
  assign RetimeWrapper_9_io_in = io_sigsIn_done; // @[package.scala 94:16:@54130.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2311 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_2311 <= 1'h0;
    end else begin
      _T_2311 <= _T_2308;
    end
  end
endmodule
module x621_inr_Switch_sm( // @[:@54292.2]
  input   clock, // @[:@54293.4]
  input   reset, // @[:@54294.4]
  input   io_enable, // @[:@54295.4]
  output  io_done, // @[:@54295.4]
  input   io_parentAck, // @[:@54295.4]
  input   io_backpressure, // @[:@54295.4]
  input   io_doneIn_0, // @[:@54295.4]
  input   io_doneIn_1, // @[:@54295.4]
  output  io_childAck_0, // @[:@54295.4]
  output  io_childAck_1, // @[:@54295.4]
  input   io_selectsIn_0, // @[:@54295.4]
  input   io_selectsIn_1, // @[:@54295.4]
  output  io_selectsOut_0, // @[:@54295.4]
  output  io_selectsOut_1 // @[:@54295.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@54297.4]
  wire  active_reset; // @[Controllers.scala 261:22:@54297.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@54297.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@54297.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@54297.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@54297.4]
  wire  done_clock; // @[Controllers.scala 262:20:@54300.4]
  wire  done_reset; // @[Controllers.scala 262:20:@54300.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@54300.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@54300.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@54300.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@54300.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@54353.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@54353.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@54353.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@54353.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@54353.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@54361.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@54361.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@54361.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@54361.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@54361.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@54371.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@54371.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@54371.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@54371.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@54371.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@54379.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@54379.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@54379.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@54379.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@54379.4]
  wire  _T_82; // @[Controllers.scala 264:62:@54307.4]
  wire  _T_103; // @[package.scala 100:49:@54333.4]
  reg  _T_120; // @[package.scala 48:56:@54349.4]
  reg [31:0] _RAND_0;
  wire  _T_125; // @[package.scala 96:25:@54358.4 package.scala 96:25:@54359.4]
  wire  _T_131; // @[package.scala 96:25:@54366.4 package.scala 96:25:@54367.4]
  wire  _T_138; // @[package.scala 96:25:@54376.4 package.scala 96:25:@54377.4]
  wire  _T_144; // @[package.scala 96:25:@54384.4 package.scala 96:25:@54385.4]
  SRFF active ( // @[Controllers.scala 261:22:@54297.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@54300.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@54353.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@54361.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@54371.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@54379.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@54307.4]
  assign _T_103 = done_io_output == 1'h0; // @[package.scala 100:49:@54333.4]
  assign _T_125 = RetimeWrapper_io_out; // @[package.scala 96:25:@54358.4 package.scala 96:25:@54359.4]
  assign _T_131 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@54366.4 package.scala 96:25:@54367.4]
  assign _T_138 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@54376.4 package.scala 96:25:@54377.4]
  assign _T_144 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@54384.4 package.scala 96:25:@54385.4]
  assign io_done = done_io_output & _T_120; // @[Controllers.scala 287:13:@54352.4]
  assign io_childAck_0 = _T_125 | _T_131; // @[Controllers.scala 288:56:@54370.4]
  assign io_childAck_1 = _T_138 | _T_144; // @[Controllers.scala 288:56:@54388.4]
  assign io_selectsOut_0 = io_selectsIn_0 & io_enable; // @[Controllers.scala 271:55:@54328.4]
  assign io_selectsOut_1 = io_selectsIn_1 & io_enable; // @[Controllers.scala 271:55:@54330.4]
  assign active_clock = clock; // @[:@54298.4]
  assign active_reset = reset; // @[:@54299.4]
  assign active_io_input_set = io_enable & _T_82; // @[Controllers.scala 264:23:@54310.4]
  assign active_io_input_reset = io_parentAck; // @[Controllers.scala 265:25:@54314.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@54315.4]
  assign done_clock = clock; // @[:@54301.4]
  assign done_reset = reset; // @[:@54302.4]
  assign done_io_input_set = io_doneIn_0 | io_doneIn_1; // @[Controllers.scala 269:50:@54326.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@54323.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@54324.4]
  assign RetimeWrapper_clock = clock; // @[:@54354.4]
  assign RetimeWrapper_reset = reset; // @[:@54355.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@54357.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@54356.4]
  assign RetimeWrapper_1_clock = clock; // @[:@54362.4]
  assign RetimeWrapper_1_reset = reset; // @[:@54363.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@54365.4]
  assign RetimeWrapper_1_io_in = 1'h0; // @[package.scala 94:16:@54364.4]
  assign RetimeWrapper_2_clock = clock; // @[:@54372.4]
  assign RetimeWrapper_2_reset = reset; // @[:@54373.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@54375.4]
  assign RetimeWrapper_2_io_in = io_doneIn_1; // @[package.scala 94:16:@54374.4]
  assign RetimeWrapper_3_clock = clock; // @[:@54380.4]
  assign RetimeWrapper_3_reset = reset; // @[:@54381.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@54383.4]
  assign RetimeWrapper_3_io_in = 1'h0; // @[package.scala 94:16:@54382.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_120 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_120 <= 1'h0;
    end else begin
      _T_120 <= _T_103;
    end
  end
endmodule
module RetimeWrapper_612( // @[:@54599.2]
  input   clock, // @[:@54600.4]
  input   reset, // @[:@54601.4]
  input   io_flow, // @[:@54602.4]
  input   io_in, // @[:@54602.4]
  output  io_out // @[:@54602.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@54604.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@54604.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@54604.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@54604.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@54604.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@54604.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(103)) sr ( // @[RetimeShiftRegister.scala 15:20:@54604.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@54617.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@54616.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@54615.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@54614.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@54613.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@54611.4]
endmodule
module RetimeWrapper_616( // @[:@54727.2]
  input   clock, // @[:@54728.4]
  input   reset, // @[:@54729.4]
  input   io_flow, // @[:@54730.4]
  input   io_in // @[:@54730.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@54732.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@54732.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@54732.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@54732.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@54732.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@54732.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(102)) sr ( // @[RetimeShiftRegister.scala 15:20:@54732.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@54744.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@54743.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@54742.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@54741.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@54739.4]
endmodule
module x619_inr_SwitchCase_sm( // @[:@54747.2]
  input   clock, // @[:@54748.4]
  input   reset, // @[:@54749.4]
  input   io_enable, // @[:@54750.4]
  output  io_done, // @[:@54750.4]
  input   io_ctrDone, // @[:@54750.4]
  output  io_datapathEn, // @[:@54750.4]
  output  io_ctrInc, // @[:@54750.4]
  input   io_parentAck, // @[:@54750.4]
  input   io_break // @[:@54750.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@54752.4]
  wire  active_reset; // @[Controllers.scala 261:22:@54752.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@54752.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@54752.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@54752.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@54752.4]
  wire  done_clock; // @[Controllers.scala 262:20:@54755.4]
  wire  done_reset; // @[Controllers.scala 262:20:@54755.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@54755.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@54755.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@54755.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@54755.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@54789.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@54789.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@54789.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@54789.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@54789.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@54811.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@54811.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@54811.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@54811.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@54811.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@54823.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@54823.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@54823.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@54823.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@54823.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@54831.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@54831.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@54831.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@54831.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@54831.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@54847.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@54847.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@54847.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@54847.4]
  wire  _T_80; // @[Controllers.scala 264:48:@54760.4]
  wire  _T_81; // @[Controllers.scala 264:46:@54761.4]
  wire  _T_82; // @[Controllers.scala 264:62:@54762.4]
  wire  _T_100; // @[package.scala 100:49:@54780.4]
  reg  _T_103; // @[package.scala 48:56:@54781.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@54804.4]
  wire  _T_124; // @[package.scala 96:25:@54816.4 package.scala 96:25:@54817.4]
  wire  _T_126; // @[package.scala 100:49:@54818.4]
  reg  _T_129; // @[package.scala 48:56:@54819.4]
  reg [31:0] _RAND_1;
  wire  _T_150; // @[package.scala 100:49:@54843.4]
  reg  _T_153; // @[package.scala 48:56:@54844.4]
  reg [31:0] _RAND_2;
  SRFF active ( // @[Controllers.scala 261:22:@54752.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@54755.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_612 RetimeWrapper ( // @[package.scala 93:22:@54789.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_612 RetimeWrapper_1 ( // @[package.scala 93:22:@54811.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@54823.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@54831.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_616 RetimeWrapper_4 ( // @[package.scala 93:22:@54847.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@54760.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@54761.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@54762.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@54780.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@54804.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@54816.4 package.scala 96:25:@54817.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@54818.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@54843.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@54822.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@54807.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@54810.4]
  assign active_clock = clock; // @[:@54753.4]
  assign active_reset = reset; // @[:@54754.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@54765.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@54769.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@54770.4]
  assign done_clock = clock; // @[:@54756.4]
  assign done_reset = reset; // @[:@54757.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@54785.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@54778.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@54779.4]
  assign RetimeWrapper_clock = clock; // @[:@54790.4]
  assign RetimeWrapper_reset = reset; // @[:@54791.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@54793.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@54792.4]
  assign RetimeWrapper_1_clock = clock; // @[:@54812.4]
  assign RetimeWrapper_1_reset = reset; // @[:@54813.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@54815.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@54814.4]
  assign RetimeWrapper_2_clock = clock; // @[:@54824.4]
  assign RetimeWrapper_2_reset = reset; // @[:@54825.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@54827.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@54826.4]
  assign RetimeWrapper_3_clock = clock; // @[:@54832.4]
  assign RetimeWrapper_3_reset = reset; // @[:@54833.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@54835.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@54834.4]
  assign RetimeWrapper_4_clock = clock; // @[:@54848.4]
  assign RetimeWrapper_4_reset = reset; // @[:@54849.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@54851.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@54850.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_153 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox_46( // @[:@54892.2]
  input  [31:0] io_a, // @[:@54895.4]
  output [54:0] io_b // @[:@54895.4]
);
  wire [21:0] _T_18; // @[SimBlackBoxes.scala 52:46:@54903.4]
  wire [44:0] tmp_frac; // @[Cat.scala 30:58:@54904.4]
  wire [9:0] new_dec; // @[SimBlackBoxes.scala 92:36:@54907.4]
  assign _T_18 = io_a[21:0]; // @[SimBlackBoxes.scala 52:46:@54903.4]
  assign tmp_frac = {_T_18,23'h0}; // @[Cat.scala 30:58:@54904.4]
  assign new_dec = io_a[31:22]; // @[SimBlackBoxes.scala 92:36:@54907.4]
  assign io_b = {new_dec,tmp_frac}; // @[SimBlackBoxes.scala 98:40:@54910.4]
endmodule
module cast_x611_div( // @[:@54912.2]
  input  [31:0] io_b, // @[:@54915.4]
  output [54:0] io_result // @[:@54915.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@54920.4]
  wire [54:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@54920.4]
  SimBlackBoxesfix2fixBox_46 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@54920.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 717:17:@54933.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@54928.4]
endmodule
module RetimeWrapper_617( // @[:@54947.2]
  input         clock, // @[:@54948.4]
  input         reset, // @[:@54949.4]
  input         io_flow, // @[:@54950.4]
  input  [54:0] io_in, // @[:@54950.4]
  output [54:0] io_out // @[:@54950.4]
);
  wire [54:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@54952.4]
  wire [54:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@54952.4]
  wire [54:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@54952.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@54952.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@54952.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@54952.4]
  RetimeShiftRegister #(.WIDTH(55), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@54952.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@54965.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@54964.4]
  assign sr_init = 55'h0; // @[RetimeShiftRegister.scala 19:16:@54963.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@54962.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@54961.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@54959.4]
endmodule
module fix2fixBox_18( // @[:@55031.2]
  input  [32:0] io_a, // @[:@55034.4]
  output [31:0] io_b // @[:@55034.4]
);
  wire [21:0] tmp_frac; // @[Converter.scala 38:42:@55042.4]
  wire [9:0] new_dec; // @[Converter.scala 88:34:@55045.4]
  assign tmp_frac = io_a[22:1]; // @[Converter.scala 38:42:@55042.4]
  assign new_dec = io_a[32:23]; // @[Converter.scala 88:34:@55045.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@55048.4]
endmodule
module x611_div( // @[:@55050.2]
  input         clock, // @[:@55051.4]
  input         reset, // @[:@55052.4]
  input  [31:0] io_a, // @[:@55053.4]
  input  [31:0] io_b, // @[:@55053.4]
  output [31:0] io_result // @[:@55053.4]
);
  wire [31:0] cast_x611_div_io_b; // @[Math.scala 720:24:@55061.4]
  wire [54:0] cast_x611_div_io_result; // @[Math.scala 720:24:@55061.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@55072.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@55072.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@55072.4]
  wire [54:0] RetimeWrapper_io_in; // @[package.scala 93:22:@55072.4]
  wire [54:0] RetimeWrapper_io_out; // @[package.scala 93:22:@55072.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@55087.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@55087.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@55087.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@55087.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@55087.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@55098.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@55098.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@55098.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@55098.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@55098.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 317:32:@55105.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 317:32:@55105.4]
  wire [54:0] _T_21_number; // @[Math.scala 723:22:@55066.4 Math.scala 724:14:@55067.4]
  wire [54:0] _T_22; // @[FixedPoint.scala 33:34:@55069.4]
  wire [31:0] _T_23; // @[FixedPoint.scala 24:59:@55070.4]
  wire [54:0] _GEN_0; // @[BigIPSim.scala 23:39:@55071.4]
  wire [55:0] _T_24; // @[BigIPSim.scala 23:39:@55071.4]
  wire [55:0] _T_25; // @[package.scala 94:23:@55075.4]
  wire [54:0] _T_28; // @[package.scala 96:25:@55079.4]
  wire [54:0] _T_29; // @[Math.scala 307:88:@55081.4]
  wire  _T_32; // @[FixedPoint.scala 50:25:@55084.4]
  wire  _T_33; // @[FixedPoint.scala 50:25:@55085.4]
  wire  _T_34; // @[Math.scala 315:58:@55086.4]
  cast_x611_div cast_x611_div ( // @[Math.scala 720:24:@55061.4]
    .io_b(cast_x611_div_io_b),
    .io_result(cast_x611_div_io_result)
  );
  RetimeWrapper_617 RetimeWrapper ( // @[package.scala 93:22:@55072.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_521 RetimeWrapper_1 ( // @[package.scala 93:22:@55087.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_521 RetimeWrapper_2 ( // @[package.scala 93:22:@55098.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  fix2fixBox_18 fix2fixBox ( // @[Math.scala 317:32:@55105.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_21_number = cast_x611_div_io_result; // @[Math.scala 723:22:@55066.4 Math.scala 724:14:@55067.4]
  assign _T_22 = $signed(_T_21_number); // @[FixedPoint.scala 33:34:@55069.4]
  assign _T_23 = $signed(io_b); // @[FixedPoint.scala 24:59:@55070.4]
  assign _GEN_0 = {{23{_T_23[31]}},_T_23}; // @[BigIPSim.scala 23:39:@55071.4]
  assign _T_24 = $signed(_T_22) / $signed(_GEN_0); // @[BigIPSim.scala 23:39:@55071.4]
  assign _T_25 = $unsigned(_T_24); // @[package.scala 94:23:@55075.4]
  assign _T_28 = $signed(RetimeWrapper_io_out); // @[package.scala 96:25:@55079.4]
  assign _T_29 = $unsigned(_T_28); // @[Math.scala 307:88:@55081.4]
  assign _T_32 = io_a[31]; // @[FixedPoint.scala 50:25:@55084.4]
  assign _T_33 = io_b[31]; // @[FixedPoint.scala 50:25:@55085.4]
  assign _T_34 = _T_32 ^ _T_33; // @[Math.scala 315:58:@55086.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 323:19:@55113.4]
  assign cast_x611_div_io_b = io_a; // @[Math.scala 721:17:@55064.4]
  assign RetimeWrapper_clock = clock; // @[:@55073.4]
  assign RetimeWrapper_reset = reset; // @[:@55074.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@55077.4]
  assign RetimeWrapper_io_in = _T_25[54:0]; // @[package.scala 94:16:@55076.4]
  assign RetimeWrapper_1_clock = clock; // @[:@55088.4]
  assign RetimeWrapper_1_reset = reset; // @[:@55089.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@55091.4]
  assign RetimeWrapper_1_io_in = _T_32 ^ _T_33; // @[package.scala 94:16:@55090.4]
  assign RetimeWrapper_2_clock = clock; // @[:@55099.4]
  assign RetimeWrapper_2_reset = reset; // @[:@55100.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@55102.4]
  assign RetimeWrapper_2_io_in = _T_34 == 1'h0; // @[package.scala 94:16:@55101.4]
  assign fix2fixBox_io_a = _T_29[32:0]; // @[Math.scala 318:25:@55108.4]
endmodule
module RetimeWrapper_620( // @[:@55127.2]
  input         clock, // @[:@55128.4]
  input         reset, // @[:@55129.4]
  input  [31:0] io_in, // @[:@55130.4]
  output [31:0] io_out // @[:@55130.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@55132.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@55132.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@55132.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@55132.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@55132.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@55132.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@55132.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@55145.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@55144.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@55143.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@55142.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@55141.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@55139.4]
endmodule
module RetimeWrapper_624( // @[:@55382.2]
  input         clock, // @[:@55383.4]
  input         reset, // @[:@55384.4]
  input  [31:0] io_in, // @[:@55385.4]
  output [31:0] io_out // @[:@55385.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@55387.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@55387.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@55387.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@55387.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@55387.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@55387.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(40)) sr ( // @[RetimeShiftRegister.scala 15:20:@55387.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@55400.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@55399.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@55398.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@55397.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@55396.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@55394.4]
endmodule
module RetimeWrapper_628( // @[:@55637.2]
  input         clock, // @[:@55638.4]
  input         reset, // @[:@55639.4]
  input  [31:0] io_in, // @[:@55640.4]
  output [31:0] io_out // @[:@55640.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@55642.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@55642.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@55642.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@55642.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@55642.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@55642.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(60)) sr ( // @[RetimeShiftRegister.scala 15:20:@55642.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@55655.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@55654.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@55653.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@55652.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@55651.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@55649.4]
endmodule
module RetimeWrapper_632( // @[:@55892.2]
  input         clock, // @[:@55893.4]
  input         reset, // @[:@55894.4]
  input  [31:0] io_in, // @[:@55895.4]
  output [31:0] io_out // @[:@55895.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@55897.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@55897.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@55897.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@55897.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@55897.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@55897.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(80)) sr ( // @[RetimeShiftRegister.scala 15:20:@55897.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@55910.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@55909.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@55908.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@55907.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@55906.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@55904.4]
endmodule
module x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1( // @[:@56806.2]
  input         clock, // @[:@56807.4]
  input         reset, // @[:@56808.4]
  output        io_in_x580_r_0_rPort_1_en_0, // @[:@56809.4]
  input  [31:0] io_in_x580_r_0_rPort_1_output_0, // @[:@56809.4]
  input         io_in_x595_reg_rPort_1_output_0, // @[:@56809.4]
  output [63:0] io_in_instrctrs_12_cycs, // @[:@56809.4]
  output [63:0] io_in_instrctrs_12_iters, // @[:@56809.4]
  input         io_sigsIn_done, // @[:@56809.4]
  input         io_sigsIn_datapathEn, // @[:@56809.4]
  input         io_sigsIn_baseEn, // @[:@56809.4]
  input         io_sigsIn_break, // @[:@56809.4]
  input         io_rr, // @[:@56809.4]
  output [31:0] io_ret_number // @[:@56809.4]
);
  wire  cycles_x619_inr_SwitchCase_clock; // @[sm_x619_inr_SwitchCase.scala 63:46:@56983.4]
  wire  cycles_x619_inr_SwitchCase_reset; // @[sm_x619_inr_SwitchCase.scala 63:46:@56983.4]
  wire  cycles_x619_inr_SwitchCase_io_enable; // @[sm_x619_inr_SwitchCase.scala 63:46:@56983.4]
  wire [63:0] cycles_x619_inr_SwitchCase_io_count; // @[sm_x619_inr_SwitchCase.scala 63:46:@56983.4]
  wire  iters_x619_inr_SwitchCase_clock; // @[sm_x619_inr_SwitchCase.scala 64:45:@56986.4]
  wire  iters_x619_inr_SwitchCase_reset; // @[sm_x619_inr_SwitchCase.scala 64:45:@56986.4]
  wire  iters_x619_inr_SwitchCase_io_enable; // @[sm_x619_inr_SwitchCase.scala 64:45:@56986.4]
  wire [63:0] iters_x619_inr_SwitchCase_io_count; // @[sm_x619_inr_SwitchCase.scala 64:45:@56986.4]
  wire  x611_div_1_clock; // @[Math.scala 327:24:@57038.4]
  wire  x611_div_1_reset; // @[Math.scala 327:24:@57038.4]
  wire [31:0] x611_div_1_io_a; // @[Math.scala 327:24:@57038.4]
  wire [31:0] x611_div_1_io_b; // @[Math.scala 327:24:@57038.4]
  wire [31:0] x611_div_1_io_result; // @[Math.scala 327:24:@57038.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@57049.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@57049.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@57049.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@57049.4]
  wire  x612_div_1_clock; // @[Math.scala 327:24:@57058.4]
  wire  x612_div_1_reset; // @[Math.scala 327:24:@57058.4]
  wire [31:0] x612_div_1_io_a; // @[Math.scala 327:24:@57058.4]
  wire [31:0] x612_div_1_io_b; // @[Math.scala 327:24:@57058.4]
  wire [31:0] x612_div_1_io_result; // @[Math.scala 327:24:@57058.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@57069.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@57069.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@57069.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@57069.4]
  wire  x613_div_1_clock; // @[Math.scala 327:24:@57078.4]
  wire  x613_div_1_reset; // @[Math.scala 327:24:@57078.4]
  wire [31:0] x613_div_1_io_a; // @[Math.scala 327:24:@57078.4]
  wire [31:0] x613_div_1_io_b; // @[Math.scala 327:24:@57078.4]
  wire [31:0] x613_div_1_io_result; // @[Math.scala 327:24:@57078.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@57089.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@57089.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@57089.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@57089.4]
  wire  x614_div_1_clock; // @[Math.scala 327:24:@57098.4]
  wire  x614_div_1_reset; // @[Math.scala 327:24:@57098.4]
  wire [31:0] x614_div_1_io_a; // @[Math.scala 327:24:@57098.4]
  wire [31:0] x614_div_1_io_b; // @[Math.scala 327:24:@57098.4]
  wire [31:0] x614_div_1_io_result; // @[Math.scala 327:24:@57098.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@57109.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@57109.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@57109.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@57109.4]
  wire  x615_div_1_clock; // @[Math.scala 327:24:@57118.4]
  wire  x615_div_1_reset; // @[Math.scala 327:24:@57118.4]
  wire [31:0] x615_div_1_io_a; // @[Math.scala 327:24:@57118.4]
  wire [31:0] x615_div_1_io_b; // @[Math.scala 327:24:@57118.4]
  wire [31:0] x615_div_1_io_result; // @[Math.scala 327:24:@57118.4]
  wire  x616_div_1_clock; // @[Math.scala 327:24:@57130.4]
  wire  x616_div_1_reset; // @[Math.scala 327:24:@57130.4]
  wire [31:0] x616_div_1_io_a; // @[Math.scala 327:24:@57130.4]
  wire [31:0] x616_div_1_io_b; // @[Math.scala 327:24:@57130.4]
  wire [31:0] x616_div_1_io_result; // @[Math.scala 327:24:@57130.4]
  wire  x617_div_1_clock; // @[Math.scala 327:24:@57140.4]
  wire  x617_div_1_reset; // @[Math.scala 327:24:@57140.4]
  wire [31:0] x617_div_1_io_a; // @[Math.scala 327:24:@57140.4]
  wire [31:0] x617_div_1_io_b; // @[Math.scala 327:24:@57140.4]
  wire [31:0] x617_div_1_io_result; // @[Math.scala 327:24:@57140.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@57151.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@57151.4]
  wire [31:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@57151.4]
  wire [31:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@57151.4]
  wire  x618_sub_1_clock; // @[Math.scala 191:24:@57160.4]
  wire  x618_sub_1_reset; // @[Math.scala 191:24:@57160.4]
  wire [31:0] x618_sub_1_io_a; // @[Math.scala 191:24:@57160.4]
  wire [31:0] x618_sub_1_io_b; // @[Math.scala 191:24:@57160.4]
  wire [31:0] x618_sub_1_io_result; // @[Math.scala 191:24:@57160.4]
  wire  _T_666; // @[package.scala 100:49:@56990.4]
  reg  _T_669; // @[package.scala 48:56:@56991.4]
  reg [31:0] _RAND_0;
  wire  _T_678; // @[sm_x619_inr_SwitchCase.scala 73:119:@57002.4]
  wire  _T_679; // @[sm_x619_inr_SwitchCase.scala 73:116:@57003.4]
  wire  _T_684; // @[implicits.scala 56:10:@57006.4]
  wire  x608_rd_x595_shared_en; // @[sm_x619_inr_SwitchCase.scala 73:136:@57007.4]
  InstrumentationCounter cycles_x619_inr_SwitchCase ( // @[sm_x619_inr_SwitchCase.scala 63:46:@56983.4]
    .clock(cycles_x619_inr_SwitchCase_clock),
    .reset(cycles_x619_inr_SwitchCase_reset),
    .io_enable(cycles_x619_inr_SwitchCase_io_enable),
    .io_count(cycles_x619_inr_SwitchCase_io_count)
  );
  InstrumentationCounter iters_x619_inr_SwitchCase ( // @[sm_x619_inr_SwitchCase.scala 64:45:@56986.4]
    .clock(iters_x619_inr_SwitchCase_clock),
    .reset(iters_x619_inr_SwitchCase_reset),
    .io_enable(iters_x619_inr_SwitchCase_io_enable),
    .io_count(iters_x619_inr_SwitchCase_io_count)
  );
  x611_div x611_div_1 ( // @[Math.scala 327:24:@57038.4]
    .clock(x611_div_1_clock),
    .reset(x611_div_1_reset),
    .io_a(x611_div_1_io_a),
    .io_b(x611_div_1_io_b),
    .io_result(x611_div_1_io_result)
  );
  RetimeWrapper_620 RetimeWrapper ( // @[package.scala 93:22:@57049.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x611_div x612_div_1 ( // @[Math.scala 327:24:@57058.4]
    .clock(x612_div_1_clock),
    .reset(x612_div_1_reset),
    .io_a(x612_div_1_io_a),
    .io_b(x612_div_1_io_b),
    .io_result(x612_div_1_io_result)
  );
  RetimeWrapper_624 RetimeWrapper_1 ( // @[package.scala 93:22:@57069.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x611_div x613_div_1 ( // @[Math.scala 327:24:@57078.4]
    .clock(x613_div_1_clock),
    .reset(x613_div_1_reset),
    .io_a(x613_div_1_io_a),
    .io_b(x613_div_1_io_b),
    .io_result(x613_div_1_io_result)
  );
  RetimeWrapper_628 RetimeWrapper_2 ( // @[package.scala 93:22:@57089.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x611_div x614_div_1 ( // @[Math.scala 327:24:@57098.4]
    .clock(x614_div_1_clock),
    .reset(x614_div_1_reset),
    .io_a(x614_div_1_io_a),
    .io_b(x614_div_1_io_b),
    .io_result(x614_div_1_io_result)
  );
  RetimeWrapper_632 RetimeWrapper_3 ( // @[package.scala 93:22:@57109.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x611_div x615_div_1 ( // @[Math.scala 327:24:@57118.4]
    .clock(x615_div_1_clock),
    .reset(x615_div_1_reset),
    .io_a(x615_div_1_io_a),
    .io_b(x615_div_1_io_b),
    .io_result(x615_div_1_io_result)
  );
  x611_div x616_div_1 ( // @[Math.scala 327:24:@57130.4]
    .clock(x616_div_1_clock),
    .reset(x616_div_1_reset),
    .io_a(x616_div_1_io_a),
    .io_b(x616_div_1_io_b),
    .io_result(x616_div_1_io_result)
  );
  x611_div x617_div_1 ( // @[Math.scala 327:24:@57140.4]
    .clock(x617_div_1_clock),
    .reset(x617_div_1_reset),
    .io_a(x617_div_1_io_a),
    .io_b(x617_div_1_io_b),
    .io_result(x617_div_1_io_result)
  );
  RetimeWrapper_628 RetimeWrapper_4 ( // @[package.scala 93:22:@57151.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x573_sub x618_sub_1 ( // @[Math.scala 191:24:@57160.4]
    .clock(x618_sub_1_clock),
    .reset(x618_sub_1_reset),
    .io_a(x618_sub_1_io_a),
    .io_b(x618_sub_1_io_b),
    .io_result(x618_sub_1_io_result)
  );
  assign _T_666 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@56990.4]
  assign _T_678 = ~ io_sigsIn_break; // @[sm_x619_inr_SwitchCase.scala 73:119:@57002.4]
  assign _T_679 = io_rr & _T_678; // @[sm_x619_inr_SwitchCase.scala 73:116:@57003.4]
  assign _T_684 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 56:10:@57006.4]
  assign x608_rd_x595_shared_en = _T_679 & _T_684; // @[sm_x619_inr_SwitchCase.scala 73:136:@57007.4]
  assign io_in_x580_r_0_rPort_1_en_0 = x608_rd_x595_shared_en & io_in_x595_reg_rPort_1_output_0; // @[MemInterfaceType.scala 110:79:@57031.4]
  assign io_in_instrctrs_12_cycs = cycles_x619_inr_SwitchCase_io_count; // @[Ledger.scala 293:21:@56995.4]
  assign io_in_instrctrs_12_iters = iters_x619_inr_SwitchCase_io_count; // @[Ledger.scala 294:22:@56996.4]
  assign io_ret_number = x618_sub_1_io_result; // @[sm_x619_inr_SwitchCase.scala 110:16:@57169.4]
  assign cycles_x619_inr_SwitchCase_clock = clock; // @[:@56984.4]
  assign cycles_x619_inr_SwitchCase_reset = reset; // @[:@56985.4]
  assign cycles_x619_inr_SwitchCase_io_enable = io_sigsIn_baseEn; // @[sm_x619_inr_SwitchCase.scala 65:44:@56989.4]
  assign iters_x619_inr_SwitchCase_clock = clock; // @[:@56987.4]
  assign iters_x619_inr_SwitchCase_reset = reset; // @[:@56988.4]
  assign iters_x619_inr_SwitchCase_io_enable = io_sigsIn_done & _T_669; // @[sm_x619_inr_SwitchCase.scala 66:43:@56994.4]
  assign x611_div_1_clock = clock; // @[:@57039.4]
  assign x611_div_1_reset = reset; // @[:@57040.4]
  assign x611_div_1_io_a = 32'h19000000; // @[Math.scala 328:17:@57041.4]
  assign x611_div_1_io_b = io_in_x580_r_0_rPort_1_output_0; // @[Math.scala 329:17:@57042.4]
  assign RetimeWrapper_clock = clock; // @[:@57050.4]
  assign RetimeWrapper_reset = reset; // @[:@57051.4]
  assign RetimeWrapper_io_in = io_in_x580_r_0_rPort_1_output_0; // @[package.scala 94:16:@57052.4]
  assign x612_div_1_clock = clock; // @[:@57059.4]
  assign x612_div_1_reset = reset; // @[:@57060.4]
  assign x612_div_1_io_a = x611_div_1_io_result; // @[Math.scala 328:17:@57061.4]
  assign x612_div_1_io_b = RetimeWrapper_io_out; // @[Math.scala 329:17:@57062.4]
  assign RetimeWrapper_1_clock = clock; // @[:@57070.4]
  assign RetimeWrapper_1_reset = reset; // @[:@57071.4]
  assign RetimeWrapper_1_io_in = io_in_x580_r_0_rPort_1_output_0; // @[package.scala 94:16:@57072.4]
  assign x613_div_1_clock = clock; // @[:@57079.4]
  assign x613_div_1_reset = reset; // @[:@57080.4]
  assign x613_div_1_io_a = x612_div_1_io_result; // @[Math.scala 328:17:@57081.4]
  assign x613_div_1_io_b = RetimeWrapper_1_io_out; // @[Math.scala 329:17:@57082.4]
  assign RetimeWrapper_2_clock = clock; // @[:@57090.4]
  assign RetimeWrapper_2_reset = reset; // @[:@57091.4]
  assign RetimeWrapper_2_io_in = io_in_x580_r_0_rPort_1_output_0; // @[package.scala 94:16:@57092.4]
  assign x614_div_1_clock = clock; // @[:@57099.4]
  assign x614_div_1_reset = reset; // @[:@57100.4]
  assign x614_div_1_io_a = x613_div_1_io_result; // @[Math.scala 328:17:@57101.4]
  assign x614_div_1_io_b = RetimeWrapper_2_io_out; // @[Math.scala 329:17:@57102.4]
  assign RetimeWrapper_3_clock = clock; // @[:@57110.4]
  assign RetimeWrapper_3_reset = reset; // @[:@57111.4]
  assign RetimeWrapper_3_io_in = io_in_x580_r_0_rPort_1_output_0; // @[package.scala 94:16:@57112.4]
  assign x615_div_1_clock = clock; // @[:@57119.4]
  assign x615_div_1_reset = reset; // @[:@57120.4]
  assign x615_div_1_io_a = x614_div_1_io_result; // @[Math.scala 328:17:@57121.4]
  assign x615_div_1_io_b = RetimeWrapper_3_io_out; // @[Math.scala 329:17:@57122.4]
  assign x616_div_1_clock = clock; // @[:@57131.4]
  assign x616_div_1_reset = reset; // @[:@57132.4]
  assign x616_div_1_io_a = 32'h2800000; // @[Math.scala 328:17:@57133.4]
  assign x616_div_1_io_b = io_in_x580_r_0_rPort_1_output_0; // @[Math.scala 329:17:@57134.4]
  assign x617_div_1_clock = clock; // @[:@57141.4]
  assign x617_div_1_reset = reset; // @[:@57142.4]
  assign x617_div_1_io_a = x616_div_1_io_result; // @[Math.scala 328:17:@57143.4]
  assign x617_div_1_io_b = RetimeWrapper_io_out; // @[Math.scala 329:17:@57144.4]
  assign RetimeWrapper_4_clock = clock; // @[:@57152.4]
  assign RetimeWrapper_4_reset = reset; // @[:@57153.4]
  assign RetimeWrapper_4_io_in = x617_div_1_io_result; // @[package.scala 94:16:@57154.4]
  assign x618_sub_1_clock = clock; // @[:@57161.4]
  assign x618_sub_1_reset = reset; // @[:@57162.4]
  assign x618_sub_1_io_a = x615_div_1_io_result; // @[Math.scala 192:17:@57163.4]
  assign x618_sub_1_io_b = RetimeWrapper_4_io_out; // @[Math.scala 193:17:@57164.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_669 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_669 <= 1'h0;
    end else begin
      _T_669 <= _T_666;
    end
  end
endmodule
module x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1( // @[:@57502.2]
  input         clock, // @[:@57503.4]
  input         reset, // @[:@57504.4]
  output [63:0] io_in_instrctrs_13_cycs, // @[:@57505.4]
  output [63:0] io_in_instrctrs_13_iters, // @[:@57505.4]
  input         io_sigsIn_done, // @[:@57505.4]
  input         io_sigsIn_baseEn // @[:@57505.4]
);
  wire  cycles_x620_inr_SwitchCase_clock; // @[sm_x620_inr_SwitchCase.scala 52:46:@57611.4]
  wire  cycles_x620_inr_SwitchCase_reset; // @[sm_x620_inr_SwitchCase.scala 52:46:@57611.4]
  wire  cycles_x620_inr_SwitchCase_io_enable; // @[sm_x620_inr_SwitchCase.scala 52:46:@57611.4]
  wire [63:0] cycles_x620_inr_SwitchCase_io_count; // @[sm_x620_inr_SwitchCase.scala 52:46:@57611.4]
  wire  iters_x620_inr_SwitchCase_clock; // @[sm_x620_inr_SwitchCase.scala 53:45:@57614.4]
  wire  iters_x620_inr_SwitchCase_reset; // @[sm_x620_inr_SwitchCase.scala 53:45:@57614.4]
  wire  iters_x620_inr_SwitchCase_io_enable; // @[sm_x620_inr_SwitchCase.scala 53:45:@57614.4]
  wire [63:0] iters_x620_inr_SwitchCase_io_count; // @[sm_x620_inr_SwitchCase.scala 53:45:@57614.4]
  wire  _T_126; // @[package.scala 100:49:@57618.4]
  reg  _T_129; // @[package.scala 48:56:@57619.4]
  reg [31:0] _RAND_0;
  InstrumentationCounter cycles_x620_inr_SwitchCase ( // @[sm_x620_inr_SwitchCase.scala 52:46:@57611.4]
    .clock(cycles_x620_inr_SwitchCase_clock),
    .reset(cycles_x620_inr_SwitchCase_reset),
    .io_enable(cycles_x620_inr_SwitchCase_io_enable),
    .io_count(cycles_x620_inr_SwitchCase_io_count)
  );
  InstrumentationCounter iters_x620_inr_SwitchCase ( // @[sm_x620_inr_SwitchCase.scala 53:45:@57614.4]
    .clock(iters_x620_inr_SwitchCase_clock),
    .reset(iters_x620_inr_SwitchCase_reset),
    .io_enable(iters_x620_inr_SwitchCase_io_enable),
    .io_count(iters_x620_inr_SwitchCase_io_count)
  );
  assign _T_126 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@57618.4]
  assign io_in_instrctrs_13_cycs = cycles_x620_inr_SwitchCase_io_count; // @[Ledger.scala 293:21:@57623.4]
  assign io_in_instrctrs_13_iters = iters_x620_inr_SwitchCase_io_count; // @[Ledger.scala 294:22:@57624.4]
  assign cycles_x620_inr_SwitchCase_clock = clock; // @[:@57612.4]
  assign cycles_x620_inr_SwitchCase_reset = reset; // @[:@57613.4]
  assign cycles_x620_inr_SwitchCase_io_enable = io_sigsIn_baseEn; // @[sm_x620_inr_SwitchCase.scala 54:44:@57617.4]
  assign iters_x620_inr_SwitchCase_clock = clock; // @[:@57615.4]
  assign iters_x620_inr_SwitchCase_reset = reset; // @[:@57616.4]
  assign iters_x620_inr_SwitchCase_io_enable = io_sigsIn_done & _T_129; // @[sm_x620_inr_SwitchCase.scala 55:43:@57622.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_129 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
  end
endmodule
module x621_inr_Switch_kernelx621_inr_Switch_concrete1( // @[:@57887.2]
  input         clock, // @[:@57888.4]
  input         reset, // @[:@57889.4]
  output        io_in_x555_tmp_1_sEn_3, // @[:@57890.4]
  output        io_in_x555_tmp_1_sDone_3, // @[:@57890.4]
  output        io_in_x554_tmp_0_sEn_3, // @[:@57890.4]
  output        io_in_x554_tmp_0_sDone_3, // @[:@57890.4]
  output        io_in_x558_tmp_4_sEn_3, // @[:@57890.4]
  output        io_in_x558_tmp_4_sDone_3, // @[:@57890.4]
  input         io_in_x736_rd_x596, // @[:@57890.4]
  output        io_in_x557_tmp_3_sEn_3, // @[:@57890.4]
  output        io_in_x557_tmp_3_sDone_3, // @[:@57890.4]
  output        io_in_x580_r_0_rPort_1_en_0, // @[:@57890.4]
  input  [31:0] io_in_x580_r_0_rPort_1_output_0, // @[:@57890.4]
  output        io_in_x580_r_0_sEn_2, // @[:@57890.4]
  output        io_in_x580_r_0_sDone_2, // @[:@57890.4]
  input         io_in_x595_reg_rPort_1_output_0, // @[:@57890.4]
  output        io_in_x595_reg_sEn_1, // @[:@57890.4]
  output        io_in_x595_reg_sDone_1, // @[:@57890.4]
  output        io_in_x556_tmp_2_sEn_3, // @[:@57890.4]
  output        io_in_x556_tmp_2_sDone_3, // @[:@57890.4]
  input         io_in_x735_rd_x595, // @[:@57890.4]
  output        io_in_x596_reg_sEn_1, // @[:@57890.4]
  output        io_in_x596_reg_sDone_1, // @[:@57890.4]
  output [63:0] io_in_instrctrs_11_cycs, // @[:@57890.4]
  output [63:0] io_in_instrctrs_11_iters, // @[:@57890.4]
  output [63:0] io_in_instrctrs_12_cycs, // @[:@57890.4]
  output [63:0] io_in_instrctrs_12_iters, // @[:@57890.4]
  output [63:0] io_in_instrctrs_13_cycs, // @[:@57890.4]
  output [63:0] io_in_instrctrs_13_iters, // @[:@57890.4]
  input         io_sigsIn_done, // @[:@57890.4]
  input         io_sigsIn_baseEn, // @[:@57890.4]
  input         io_sigsIn_smSelectsOut_0, // @[:@57890.4]
  input         io_sigsIn_smSelectsOut_1, // @[:@57890.4]
  input         io_sigsIn_smChildAcks_0, // @[:@57890.4]
  input         io_sigsIn_smChildAcks_1, // @[:@57890.4]
  output        io_sigsOut_smDoneIn_0, // @[:@57890.4]
  output        io_sigsOut_smDoneIn_1, // @[:@57890.4]
  input         io_rr, // @[:@57890.4]
  output [31:0] io_ret_number // @[:@57890.4]
);
  wire  cycles_x621_inr_Switch_clock; // @[sm_x621_inr_Switch.scala 96:42:@58309.4]
  wire  cycles_x621_inr_Switch_reset; // @[sm_x621_inr_Switch.scala 96:42:@58309.4]
  wire  cycles_x621_inr_Switch_io_enable; // @[sm_x621_inr_Switch.scala 96:42:@58309.4]
  wire [63:0] cycles_x621_inr_Switch_io_count; // @[sm_x621_inr_Switch.scala 96:42:@58309.4]
  wire  iters_x621_inr_Switch_clock; // @[sm_x621_inr_Switch.scala 97:41:@58312.4]
  wire  iters_x621_inr_Switch_reset; // @[sm_x621_inr_Switch.scala 97:41:@58312.4]
  wire  iters_x621_inr_Switch_io_enable; // @[sm_x621_inr_Switch.scala 97:41:@58312.4]
  wire [63:0] iters_x621_inr_Switch_io_count; // @[sm_x621_inr_Switch.scala 97:41:@58312.4]
  wire  x619_inr_SwitchCase_sm_clock; // @[sm_x619_inr_SwitchCase.scala 32:18:@58361.4]
  wire  x619_inr_SwitchCase_sm_reset; // @[sm_x619_inr_SwitchCase.scala 32:18:@58361.4]
  wire  x619_inr_SwitchCase_sm_io_enable; // @[sm_x619_inr_SwitchCase.scala 32:18:@58361.4]
  wire  x619_inr_SwitchCase_sm_io_done; // @[sm_x619_inr_SwitchCase.scala 32:18:@58361.4]
  wire  x619_inr_SwitchCase_sm_io_ctrDone; // @[sm_x619_inr_SwitchCase.scala 32:18:@58361.4]
  wire  x619_inr_SwitchCase_sm_io_datapathEn; // @[sm_x619_inr_SwitchCase.scala 32:18:@58361.4]
  wire  x619_inr_SwitchCase_sm_io_ctrInc; // @[sm_x619_inr_SwitchCase.scala 32:18:@58361.4]
  wire  x619_inr_SwitchCase_sm_io_parentAck; // @[sm_x619_inr_SwitchCase.scala 32:18:@58361.4]
  wire  x619_inr_SwitchCase_sm_io_break; // @[sm_x619_inr_SwitchCase.scala 32:18:@58361.4]
  wire  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_clock; // @[sm_x619_inr_SwitchCase.scala 112:24:@58439.4]
  wire  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_reset; // @[sm_x619_inr_SwitchCase.scala 112:24:@58439.4]
  wire  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x580_r_0_rPort_1_en_0; // @[sm_x619_inr_SwitchCase.scala 112:24:@58439.4]
  wire [31:0] x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x580_r_0_rPort_1_output_0; // @[sm_x619_inr_SwitchCase.scala 112:24:@58439.4]
  wire  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x595_reg_rPort_1_output_0; // @[sm_x619_inr_SwitchCase.scala 112:24:@58439.4]
  wire [63:0] x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_instrctrs_12_cycs; // @[sm_x619_inr_SwitchCase.scala 112:24:@58439.4]
  wire [63:0] x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_instrctrs_12_iters; // @[sm_x619_inr_SwitchCase.scala 112:24:@58439.4]
  wire  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_done; // @[sm_x619_inr_SwitchCase.scala 112:24:@58439.4]
  wire  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_datapathEn; // @[sm_x619_inr_SwitchCase.scala 112:24:@58439.4]
  wire  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_baseEn; // @[sm_x619_inr_SwitchCase.scala 112:24:@58439.4]
  wire  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_break; // @[sm_x619_inr_SwitchCase.scala 112:24:@58439.4]
  wire  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_rr; // @[sm_x619_inr_SwitchCase.scala 112:24:@58439.4]
  wire [31:0] x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_ret_number; // @[sm_x619_inr_SwitchCase.scala 112:24:@58439.4]
  wire  x620_inr_SwitchCase_sm_clock; // @[sm_x620_inr_SwitchCase.scala 31:18:@58745.4]
  wire  x620_inr_SwitchCase_sm_reset; // @[sm_x620_inr_SwitchCase.scala 31:18:@58745.4]
  wire  x620_inr_SwitchCase_sm_io_enable; // @[sm_x620_inr_SwitchCase.scala 31:18:@58745.4]
  wire  x620_inr_SwitchCase_sm_io_done; // @[sm_x620_inr_SwitchCase.scala 31:18:@58745.4]
  wire  x620_inr_SwitchCase_sm_io_ctrDone; // @[sm_x620_inr_SwitchCase.scala 31:18:@58745.4]
  wire  x620_inr_SwitchCase_sm_io_datapathEn; // @[sm_x620_inr_SwitchCase.scala 31:18:@58745.4]
  wire  x620_inr_SwitchCase_sm_io_ctrInc; // @[sm_x620_inr_SwitchCase.scala 31:18:@58745.4]
  wire  x620_inr_SwitchCase_sm_io_parentAck; // @[sm_x620_inr_SwitchCase.scala 31:18:@58745.4]
  wire  x620_inr_SwitchCase_sm_io_break; // @[sm_x620_inr_SwitchCase.scala 31:18:@58745.4]
  wire  x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_clock; // @[sm_x620_inr_SwitchCase.scala 60:24:@58823.4]
  wire  x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_reset; // @[sm_x620_inr_SwitchCase.scala 60:24:@58823.4]
  wire [63:0] x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_io_in_instrctrs_13_cycs; // @[sm_x620_inr_SwitchCase.scala 60:24:@58823.4]
  wire [63:0] x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_io_in_instrctrs_13_iters; // @[sm_x620_inr_SwitchCase.scala 60:24:@58823.4]
  wire  x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_io_sigsIn_done; // @[sm_x620_inr_SwitchCase.scala 60:24:@58823.4]
  wire  x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_io_sigsIn_baseEn; // @[sm_x620_inr_SwitchCase.scala 60:24:@58823.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@58999.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@58999.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@58999.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@58999.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@58999.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@59010.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@59010.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@59010.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@59010.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@59010.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@59021.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@59021.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@59021.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@59021.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@59021.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@59032.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@59032.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@59032.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@59032.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@59032.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@59043.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@59043.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@59043.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@59043.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@59043.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@59054.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@59054.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@59054.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@59054.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@59054.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@59065.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@59065.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@59065.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@59065.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@59065.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@59076.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@59076.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@59076.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@59076.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@59076.4]
  wire  _T_2310; // @[package.scala 100:49:@58316.4]
  reg  _T_2313; // @[package.scala 48:56:@58317.4]
  reg [31:0] _RAND_0;
  wire  _T_2375; // @[package.scala 100:49:@58390.4]
  reg  _T_2378; // @[package.scala 48:56:@58391.4]
  reg [31:0] _RAND_1;
  wire  _T_2458; // @[package.scala 100:49:@58774.4]
  reg  _T_2461; // @[package.scala 48:56:@58775.4]
  reg [31:0] _RAND_2;
  wire [31:0] x619_inr_SwitchCase_number; // @[sm_x621_inr_Switch.scala 108:37:@58402.4 sm_x621_inr_Switch.scala 111:29:@58708.4]
  wire [31:0] _T_2499; // @[Mux.scala 19:72:@58989.4]
  wire [31:0] _T_2501; // @[Mux.scala 19:72:@58990.4]
  wire  _T_2511; // @[package.scala 96:25:@59004.4 package.scala 96:25:@59005.4]
  wire  _T_2517; // @[package.scala 96:25:@59015.4 package.scala 96:25:@59016.4]
  wire  _T_2523; // @[package.scala 96:25:@59026.4 package.scala 96:25:@59027.4]
  wire  _T_2529; // @[package.scala 96:25:@59037.4 package.scala 96:25:@59038.4]
  wire  _T_2535; // @[package.scala 96:25:@59048.4 package.scala 96:25:@59049.4]
  wire  _T_2541; // @[package.scala 96:25:@59059.4 package.scala 96:25:@59060.4]
  wire  _T_2547; // @[package.scala 96:25:@59070.4 package.scala 96:25:@59071.4]
  wire  _T_2553; // @[package.scala 96:25:@59081.4 package.scala 96:25:@59082.4]
  InstrumentationCounter cycles_x621_inr_Switch ( // @[sm_x621_inr_Switch.scala 96:42:@58309.4]
    .clock(cycles_x621_inr_Switch_clock),
    .reset(cycles_x621_inr_Switch_reset),
    .io_enable(cycles_x621_inr_Switch_io_enable),
    .io_count(cycles_x621_inr_Switch_io_count)
  );
  InstrumentationCounter iters_x621_inr_Switch ( // @[sm_x621_inr_Switch.scala 97:41:@58312.4]
    .clock(iters_x621_inr_Switch_clock),
    .reset(iters_x621_inr_Switch_reset),
    .io_enable(iters_x621_inr_Switch_io_enable),
    .io_count(iters_x621_inr_Switch_io_count)
  );
  x619_inr_SwitchCase_sm x619_inr_SwitchCase_sm ( // @[sm_x619_inr_SwitchCase.scala 32:18:@58361.4]
    .clock(x619_inr_SwitchCase_sm_clock),
    .reset(x619_inr_SwitchCase_sm_reset),
    .io_enable(x619_inr_SwitchCase_sm_io_enable),
    .io_done(x619_inr_SwitchCase_sm_io_done),
    .io_ctrDone(x619_inr_SwitchCase_sm_io_ctrDone),
    .io_datapathEn(x619_inr_SwitchCase_sm_io_datapathEn),
    .io_ctrInc(x619_inr_SwitchCase_sm_io_ctrInc),
    .io_parentAck(x619_inr_SwitchCase_sm_io_parentAck),
    .io_break(x619_inr_SwitchCase_sm_io_break)
  );
  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1 x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1 ( // @[sm_x619_inr_SwitchCase.scala 112:24:@58439.4]
    .clock(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_clock),
    .reset(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_reset),
    .io_in_x580_r_0_rPort_1_en_0(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x580_r_0_rPort_1_en_0),
    .io_in_x580_r_0_rPort_1_output_0(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x580_r_0_rPort_1_output_0),
    .io_in_x595_reg_rPort_1_output_0(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x595_reg_rPort_1_output_0),
    .io_in_instrctrs_12_cycs(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_instrctrs_12_cycs),
    .io_in_instrctrs_12_iters(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_instrctrs_12_iters),
    .io_sigsIn_done(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_done),
    .io_sigsIn_datapathEn(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_break),
    .io_rr(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_rr),
    .io_ret_number(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_ret_number)
  );
  x619_inr_SwitchCase_sm x620_inr_SwitchCase_sm ( // @[sm_x620_inr_SwitchCase.scala 31:18:@58745.4]
    .clock(x620_inr_SwitchCase_sm_clock),
    .reset(x620_inr_SwitchCase_sm_reset),
    .io_enable(x620_inr_SwitchCase_sm_io_enable),
    .io_done(x620_inr_SwitchCase_sm_io_done),
    .io_ctrDone(x620_inr_SwitchCase_sm_io_ctrDone),
    .io_datapathEn(x620_inr_SwitchCase_sm_io_datapathEn),
    .io_ctrInc(x620_inr_SwitchCase_sm_io_ctrInc),
    .io_parentAck(x620_inr_SwitchCase_sm_io_parentAck),
    .io_break(x620_inr_SwitchCase_sm_io_break)
  );
  x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1 x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1 ( // @[sm_x620_inr_SwitchCase.scala 60:24:@58823.4]
    .clock(x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_clock),
    .reset(x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_reset),
    .io_in_instrctrs_13_cycs(x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_io_in_instrctrs_13_cycs),
    .io_in_instrctrs_13_iters(x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_io_in_instrctrs_13_iters),
    .io_sigsIn_done(x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_io_sigsIn_baseEn)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@58999.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@59010.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@59021.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@59032.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@59043.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@59054.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@59065.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@59076.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign _T_2310 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@58316.4]
  assign _T_2375 = x619_inr_SwitchCase_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@58390.4]
  assign _T_2458 = x620_inr_SwitchCase_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@58774.4]
  assign x619_inr_SwitchCase_number = x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_ret_number; // @[sm_x621_inr_Switch.scala 108:37:@58402.4 sm_x621_inr_Switch.scala 111:29:@58708.4]
  assign _T_2499 = io_in_x735_rd_x595 ? x619_inr_SwitchCase_number : 32'h0; // @[Mux.scala 19:72:@58989.4]
  assign _T_2501 = io_in_x736_rd_x596 ? 32'h16800000 : 32'h0; // @[Mux.scala 19:72:@58990.4]
  assign _T_2511 = RetimeWrapper_io_out; // @[package.scala 96:25:@59004.4 package.scala 96:25:@59005.4]
  assign _T_2517 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@59015.4 package.scala 96:25:@59016.4]
  assign _T_2523 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@59026.4 package.scala 96:25:@59027.4]
  assign _T_2529 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@59037.4 package.scala 96:25:@59038.4]
  assign _T_2535 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@59048.4 package.scala 96:25:@59049.4]
  assign _T_2541 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@59059.4 package.scala 96:25:@59060.4]
  assign _T_2547 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@59070.4 package.scala 96:25:@59071.4]
  assign _T_2553 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@59081.4 package.scala 96:25:@59082.4]
  assign io_in_x555_tmp_1_sEn_3 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@59018.4]
  assign io_in_x555_tmp_1_sDone_3 = io_rr ? _T_2517 : 1'h0; // @[MemInterfaceType.scala 197:17:@59019.4]
  assign io_in_x554_tmp_0_sEn_3 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@59007.4]
  assign io_in_x554_tmp_0_sDone_3 = io_rr ? _T_2511 : 1'h0; // @[MemInterfaceType.scala 197:17:@59008.4]
  assign io_in_x558_tmp_4_sEn_3 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@59051.4]
  assign io_in_x558_tmp_4_sDone_3 = io_rr ? _T_2535 : 1'h0; // @[MemInterfaceType.scala 197:17:@59052.4]
  assign io_in_x557_tmp_3_sEn_3 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@59040.4]
  assign io_in_x557_tmp_3_sDone_3 = io_rr ? _T_2529 : 1'h0; // @[MemInterfaceType.scala 197:17:@59041.4]
  assign io_in_x580_r_0_rPort_1_en_0 = x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x580_r_0_rPort_1_en_0; // @[MemInterfaceType.scala 66:44:@58653.4]
  assign io_in_x580_r_0_sEn_2 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@59062.4]
  assign io_in_x580_r_0_sDone_2 = io_rr ? _T_2541 : 1'h0; // @[MemInterfaceType.scala 197:17:@59063.4]
  assign io_in_x595_reg_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@59073.4]
  assign io_in_x595_reg_sDone_1 = io_rr ? _T_2547 : 1'h0; // @[MemInterfaceType.scala 197:17:@59074.4]
  assign io_in_x556_tmp_2_sEn_3 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@59029.4]
  assign io_in_x556_tmp_2_sDone_3 = io_rr ? _T_2523 : 1'h0; // @[MemInterfaceType.scala 197:17:@59030.4]
  assign io_in_x596_reg_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@59084.4]
  assign io_in_x596_reg_sDone_1 = io_rr ? _T_2553 : 1'h0; // @[MemInterfaceType.scala 197:17:@59085.4]
  assign io_in_instrctrs_11_cycs = cycles_x621_inr_Switch_io_count; // @[Ledger.scala 293:21:@58321.4]
  assign io_in_instrctrs_11_iters = iters_x621_inr_Switch_io_count; // @[Ledger.scala 294:22:@58322.4]
  assign io_in_instrctrs_12_cycs = x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_instrctrs_12_cycs; // @[Ledger.scala 302:78:@58680.4]
  assign io_in_instrctrs_12_iters = x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_instrctrs_12_iters; // @[Ledger.scala 302:78:@58679.4]
  assign io_in_instrctrs_13_cycs = x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_io_in_instrctrs_13_cycs; // @[Ledger.scala 302:78:@58954.4]
  assign io_in_instrctrs_13_iters = x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_io_in_instrctrs_13_iters; // @[Ledger.scala 302:78:@58953.4]
  assign io_sigsOut_smDoneIn_0 = x619_inr_SwitchCase_sm_io_done; // @[SpatialBlocks.scala 155:56:@58425.4]
  assign io_sigsOut_smDoneIn_1 = x620_inr_SwitchCase_sm_io_done; // @[SpatialBlocks.scala 155:56:@58809.4]
  assign io_ret_number = _T_2499 | _T_2501; // @[sm_x621_inr_Switch.scala 129:16:@58997.4]
  assign cycles_x621_inr_Switch_clock = clock; // @[:@58310.4]
  assign cycles_x621_inr_Switch_reset = reset; // @[:@58311.4]
  assign cycles_x621_inr_Switch_io_enable = io_sigsIn_baseEn; // @[sm_x621_inr_Switch.scala 98:40:@58315.4]
  assign iters_x621_inr_Switch_clock = clock; // @[:@58313.4]
  assign iters_x621_inr_Switch_reset = reset; // @[:@58314.4]
  assign iters_x621_inr_Switch_io_enable = io_sigsIn_done & _T_2313; // @[sm_x621_inr_Switch.scala 99:39:@58320.4]
  assign x619_inr_SwitchCase_sm_clock = clock; // @[:@58362.4]
  assign x619_inr_SwitchCase_sm_reset = reset; // @[:@58363.4]
  assign x619_inr_SwitchCase_sm_io_enable = io_sigsIn_smSelectsOut_0; // @[SpatialBlocks.scala 139:18:@58422.4]
  assign x619_inr_SwitchCase_sm_io_ctrDone = x619_inr_SwitchCase_sm_io_ctrInc & _T_2378; // @[sm_x621_inr_Switch.scala 103:45:@58394.4]
  assign x619_inr_SwitchCase_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@58424.4]
  assign x619_inr_SwitchCase_sm_io_break = 1'h0; // @[sm_x621_inr_Switch.scala 107:43:@58401.4]
  assign x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_clock = clock; // @[:@58440.4]
  assign x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_reset = reset; // @[:@58441.4]
  assign x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x580_r_0_rPort_1_output_0 = io_in_x580_r_0_rPort_1_output_0; // @[MemInterfaceType.scala 66:44:@58651.4]
  assign x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x595_reg_rPort_1_output_0 = io_in_x595_reg_rPort_1_output_0; // @[MemInterfaceType.scala 66:44:@58672.4]
  assign x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_done = x619_inr_SwitchCase_sm_io_done; // @[sm_x619_inr_SwitchCase.scala 118:22:@58700.4]
  assign x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_datapathEn = x619_inr_SwitchCase_sm_io_datapathEn; // @[sm_x619_inr_SwitchCase.scala 118:22:@58693.4]
  assign x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_baseEn = io_sigsIn_smSelectsOut_0; // @[sm_x619_inr_SwitchCase.scala 118:22:@58692.4]
  assign x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_break = x619_inr_SwitchCase_sm_io_break; // @[sm_x619_inr_SwitchCase.scala 118:22:@58691.4]
  assign x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_rr = io_rr; // @[sm_x619_inr_SwitchCase.scala 117:18:@58681.4]
  assign x620_inr_SwitchCase_sm_clock = clock; // @[:@58746.4]
  assign x620_inr_SwitchCase_sm_reset = reset; // @[:@58747.4]
  assign x620_inr_SwitchCase_sm_io_enable = io_sigsIn_smSelectsOut_1; // @[SpatialBlocks.scala 139:18:@58806.4]
  assign x620_inr_SwitchCase_sm_io_ctrDone = x620_inr_SwitchCase_sm_io_ctrInc & _T_2461; // @[sm_x621_inr_Switch.scala 114:45:@58778.4]
  assign x620_inr_SwitchCase_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 141:21:@58808.4]
  assign x620_inr_SwitchCase_sm_io_break = 1'h0; // @[sm_x621_inr_Switch.scala 118:43:@58785.4]
  assign x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_clock = clock; // @[:@58824.4]
  assign x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_reset = reset; // @[:@58825.4]
  assign x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_io_sigsIn_done = x620_inr_SwitchCase_sm_io_done; // @[sm_x620_inr_SwitchCase.scala 65:22:@58974.4]
  assign x620_inr_SwitchCase_kernelx620_inr_SwitchCase_concrete1_io_sigsIn_baseEn = io_sigsIn_smSelectsOut_1; // @[sm_x620_inr_SwitchCase.scala 65:22:@58966.4]
  assign RetimeWrapper_clock = clock; // @[:@59000.4]
  assign RetimeWrapper_reset = reset; // @[:@59001.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@59003.4]
  assign RetimeWrapper_io_in = io_sigsIn_done; // @[package.scala 94:16:@59002.4]
  assign RetimeWrapper_1_clock = clock; // @[:@59011.4]
  assign RetimeWrapper_1_reset = reset; // @[:@59012.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@59014.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_done; // @[package.scala 94:16:@59013.4]
  assign RetimeWrapper_2_clock = clock; // @[:@59022.4]
  assign RetimeWrapper_2_reset = reset; // @[:@59023.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@59025.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_done; // @[package.scala 94:16:@59024.4]
  assign RetimeWrapper_3_clock = clock; // @[:@59033.4]
  assign RetimeWrapper_3_reset = reset; // @[:@59034.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@59036.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_done; // @[package.scala 94:16:@59035.4]
  assign RetimeWrapper_4_clock = clock; // @[:@59044.4]
  assign RetimeWrapper_4_reset = reset; // @[:@59045.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@59047.4]
  assign RetimeWrapper_4_io_in = io_sigsIn_done; // @[package.scala 94:16:@59046.4]
  assign RetimeWrapper_5_clock = clock; // @[:@59055.4]
  assign RetimeWrapper_5_reset = reset; // @[:@59056.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@59058.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_done; // @[package.scala 94:16:@59057.4]
  assign RetimeWrapper_6_clock = clock; // @[:@59066.4]
  assign RetimeWrapper_6_reset = reset; // @[:@59067.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@59069.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_done; // @[package.scala 94:16:@59068.4]
  assign RetimeWrapper_7_clock = clock; // @[:@59077.4]
  assign RetimeWrapper_7_reset = reset; // @[:@59078.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@59080.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_done; // @[package.scala 94:16:@59079.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2313 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_2378 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2461 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_2313 <= 1'h0;
    end else begin
      _T_2313 <= _T_2310;
    end
    if (reset) begin
      _T_2378 <= 1'h0;
    end else begin
      _T_2378 <= _T_2375;
    end
    if (reset) begin
      _T_2461 <= 1'h0;
    end else begin
      _T_2461 <= _T_2458;
    end
  end
endmodule
module x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1( // @[:@59699.2]
  input         clock, // @[:@59700.4]
  input         reset, // @[:@59701.4]
  output        io_in_x555_tmp_1_sEn_4, // @[:@59702.4]
  output        io_in_x555_tmp_1_sDone_4, // @[:@59702.4]
  output        io_in_x554_tmp_0_sEn_4, // @[:@59702.4]
  output        io_in_x554_tmp_0_sDone_4, // @[:@59702.4]
  output        io_in_x558_tmp_4_sEn_4, // @[:@59702.4]
  output        io_in_x558_tmp_4_sDone_4, // @[:@59702.4]
  output [31:0] io_in_x594_force_0_wPort_0_data_0, // @[:@59702.4]
  output        io_in_x594_force_0_wPort_0_en_0, // @[:@59702.4]
  output        io_in_x594_force_0_sEn_0, // @[:@59702.4]
  output        io_in_x594_force_0_sDone_0, // @[:@59702.4]
  input  [31:0] io_in_x621_inr_Switch_number, // @[:@59702.4]
  output        io_in_x557_tmp_3_sEn_4, // @[:@59702.4]
  output        io_in_x557_tmp_3_sDone_4, // @[:@59702.4]
  output        io_in_x556_tmp_2_sEn_4, // @[:@59702.4]
  output        io_in_x556_tmp_2_sDone_4, // @[:@59702.4]
  output [63:0] io_in_instrctrs_14_cycs, // @[:@59702.4]
  output [63:0] io_in_instrctrs_14_iters, // @[:@59702.4]
  input         io_sigsIn_done, // @[:@59702.4]
  input         io_sigsIn_datapathEn, // @[:@59702.4]
  input         io_sigsIn_baseEn, // @[:@59702.4]
  input         io_sigsIn_break, // @[:@59702.4]
  input         io_rr // @[:@59702.4]
);
  wire  cycles_x623_inr_UnitPipe_clock; // @[sm_x623_inr_UnitPipe.scala 92:44:@60051.4]
  wire  cycles_x623_inr_UnitPipe_reset; // @[sm_x623_inr_UnitPipe.scala 92:44:@60051.4]
  wire  cycles_x623_inr_UnitPipe_io_enable; // @[sm_x623_inr_UnitPipe.scala 92:44:@60051.4]
  wire [63:0] cycles_x623_inr_UnitPipe_io_count; // @[sm_x623_inr_UnitPipe.scala 92:44:@60051.4]
  wire  iters_x623_inr_UnitPipe_clock; // @[sm_x623_inr_UnitPipe.scala 93:43:@60054.4]
  wire  iters_x623_inr_UnitPipe_reset; // @[sm_x623_inr_UnitPipe.scala 93:43:@60054.4]
  wire  iters_x623_inr_UnitPipe_io_enable; // @[sm_x623_inr_UnitPipe.scala 93:43:@60054.4]
  wire [63:0] iters_x623_inr_UnitPipe_io_count; // @[sm_x623_inr_UnitPipe.scala 93:43:@60054.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@60087.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@60087.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@60087.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@60087.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@60087.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@60098.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@60098.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@60098.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@60098.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@60098.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@60109.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@60109.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@60109.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@60109.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@60109.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@60120.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@60120.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@60120.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@60120.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@60120.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@60131.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@60131.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@60131.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@60131.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@60131.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@60142.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@60142.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@60142.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@60142.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@60142.4]
  wire  _T_1770; // @[package.scala 100:49:@60058.4]
  reg  _T_1773; // @[package.scala 48:56:@60059.4]
  reg [31:0] _RAND_0;
  wire  _T_1785; // @[sm_x623_inr_UnitPipe.scala 101:100:@60071.4]
  wire  _T_1791; // @[implicits.scala 56:10:@60075.4]
  wire  _T_1792; // @[sm_x623_inr_UnitPipe.scala 101:117:@60076.4]
  wire  _T_1801; // @[package.scala 96:25:@60092.4 package.scala 96:25:@60093.4]
  wire  _T_1807; // @[package.scala 96:25:@60103.4 package.scala 96:25:@60104.4]
  wire  _T_1813; // @[package.scala 96:25:@60114.4 package.scala 96:25:@60115.4]
  wire  _T_1819; // @[package.scala 96:25:@60125.4 package.scala 96:25:@60126.4]
  wire  _T_1825; // @[package.scala 96:25:@60136.4 package.scala 96:25:@60137.4]
  wire  _T_1831; // @[package.scala 96:25:@60147.4 package.scala 96:25:@60148.4]
  InstrumentationCounter cycles_x623_inr_UnitPipe ( // @[sm_x623_inr_UnitPipe.scala 92:44:@60051.4]
    .clock(cycles_x623_inr_UnitPipe_clock),
    .reset(cycles_x623_inr_UnitPipe_reset),
    .io_enable(cycles_x623_inr_UnitPipe_io_enable),
    .io_count(cycles_x623_inr_UnitPipe_io_count)
  );
  InstrumentationCounter iters_x623_inr_UnitPipe ( // @[sm_x623_inr_UnitPipe.scala 93:43:@60054.4]
    .clock(iters_x623_inr_UnitPipe_clock),
    .reset(iters_x623_inr_UnitPipe_reset),
    .io_enable(iters_x623_inr_UnitPipe_io_enable),
    .io_count(iters_x623_inr_UnitPipe_io_count)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@60087.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@60098.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@60109.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@60120.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@60131.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@60142.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  assign _T_1770 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@60058.4]
  assign _T_1785 = ~ io_sigsIn_break; // @[sm_x623_inr_UnitPipe.scala 101:100:@60071.4]
  assign _T_1791 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 56:10:@60075.4]
  assign _T_1792 = _T_1785 & _T_1791; // @[sm_x623_inr_UnitPipe.scala 101:117:@60076.4]
  assign _T_1801 = RetimeWrapper_io_out; // @[package.scala 96:25:@60092.4 package.scala 96:25:@60093.4]
  assign _T_1807 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@60103.4 package.scala 96:25:@60104.4]
  assign _T_1813 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@60114.4 package.scala 96:25:@60115.4]
  assign _T_1819 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@60125.4 package.scala 96:25:@60126.4]
  assign _T_1825 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@60136.4 package.scala 96:25:@60137.4]
  assign _T_1831 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@60147.4 package.scala 96:25:@60148.4]
  assign io_in_x555_tmp_1_sEn_4 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@60106.4]
  assign io_in_x555_tmp_1_sDone_4 = io_rr ? _T_1807 : 1'h0; // @[MemInterfaceType.scala 197:17:@60107.4]
  assign io_in_x554_tmp_0_sEn_4 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@60095.4]
  assign io_in_x554_tmp_0_sDone_4 = io_rr ? _T_1801 : 1'h0; // @[MemInterfaceType.scala 197:17:@60096.4]
  assign io_in_x558_tmp_4_sEn_4 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@60139.4]
  assign io_in_x558_tmp_4_sDone_4 = io_rr ? _T_1825 : 1'h0; // @[MemInterfaceType.scala 197:17:@60140.4]
  assign io_in_x594_force_0_wPort_0_data_0 = io_in_x621_inr_Switch_number; // @[MemInterfaceType.scala 90:56:@60083.4]
  assign io_in_x594_force_0_wPort_0_en_0 = _T_1792 & _T_1785; // @[MemInterfaceType.scala 93:57:@60085.4]
  assign io_in_x594_force_0_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@60150.4]
  assign io_in_x594_force_0_sDone_0 = io_rr ? _T_1831 : 1'h0; // @[MemInterfaceType.scala 197:17:@60151.4]
  assign io_in_x557_tmp_3_sEn_4 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@60128.4]
  assign io_in_x557_tmp_3_sDone_4 = io_rr ? _T_1819 : 1'h0; // @[MemInterfaceType.scala 197:17:@60129.4]
  assign io_in_x556_tmp_2_sEn_4 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@60117.4]
  assign io_in_x556_tmp_2_sDone_4 = io_rr ? _T_1813 : 1'h0; // @[MemInterfaceType.scala 197:17:@60118.4]
  assign io_in_instrctrs_14_cycs = cycles_x623_inr_UnitPipe_io_count; // @[Ledger.scala 293:21:@60063.4]
  assign io_in_instrctrs_14_iters = iters_x623_inr_UnitPipe_io_count; // @[Ledger.scala 294:22:@60064.4]
  assign cycles_x623_inr_UnitPipe_clock = clock; // @[:@60052.4]
  assign cycles_x623_inr_UnitPipe_reset = reset; // @[:@60053.4]
  assign cycles_x623_inr_UnitPipe_io_enable = io_sigsIn_baseEn; // @[sm_x623_inr_UnitPipe.scala 94:42:@60057.4]
  assign iters_x623_inr_UnitPipe_clock = clock; // @[:@60055.4]
  assign iters_x623_inr_UnitPipe_reset = reset; // @[:@60056.4]
  assign iters_x623_inr_UnitPipe_io_enable = io_sigsIn_done & _T_1773; // @[sm_x623_inr_UnitPipe.scala 95:41:@60062.4]
  assign RetimeWrapper_clock = clock; // @[:@60088.4]
  assign RetimeWrapper_reset = reset; // @[:@60089.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@60091.4]
  assign RetimeWrapper_io_in = io_sigsIn_done; // @[package.scala 94:16:@60090.4]
  assign RetimeWrapper_1_clock = clock; // @[:@60099.4]
  assign RetimeWrapper_1_reset = reset; // @[:@60100.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@60102.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_done; // @[package.scala 94:16:@60101.4]
  assign RetimeWrapper_2_clock = clock; // @[:@60110.4]
  assign RetimeWrapper_2_reset = reset; // @[:@60111.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@60113.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_done; // @[package.scala 94:16:@60112.4]
  assign RetimeWrapper_3_clock = clock; // @[:@60121.4]
  assign RetimeWrapper_3_reset = reset; // @[:@60122.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@60124.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_done; // @[package.scala 94:16:@60123.4]
  assign RetimeWrapper_4_clock = clock; // @[:@60132.4]
  assign RetimeWrapper_4_reset = reset; // @[:@60133.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@60135.4]
  assign RetimeWrapper_4_io_in = io_sigsIn_done; // @[package.scala 94:16:@60134.4]
  assign RetimeWrapper_5_clock = clock; // @[:@60143.4]
  assign RetimeWrapper_5_reset = reset; // @[:@60144.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@60146.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_done; // @[package.scala 94:16:@60145.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1773 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1773 <= 1'h0;
    end else begin
      _T_1773 <= _T_1770;
    end
  end
endmodule
module RetimeWrapper_671( // @[:@60354.2]
  input   clock, // @[:@60355.4]
  input   reset, // @[:@60356.4]
  input   io_in, // @[:@60357.4]
  output  io_out // @[:@60357.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@60359.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@60359.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@60359.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@60359.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@60359.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@60359.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(15)) sr ( // @[RetimeShiftRegister.scala 15:20:@60359.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@60372.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@60371.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@60370.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@60369.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@60368.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@60366.4]
endmodule
module RetimeWrapper_675( // @[:@60482.2]
  input   clock, // @[:@60483.4]
  input   reset, // @[:@60484.4]
  input   io_in, // @[:@60485.4]
  output  io_out // @[:@60485.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@60487.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@60487.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@60487.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@60487.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@60487.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@60487.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(14)) sr ( // @[RetimeShiftRegister.scala 15:20:@60487.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@60500.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@60499.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@60498.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@60497.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@60496.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@60494.4]
endmodule
module x639_inr_Foreach_sm( // @[:@60502.2]
  input   clock, // @[:@60503.4]
  input   reset, // @[:@60504.4]
  input   io_enable, // @[:@60505.4]
  output  io_done, // @[:@60505.4]
  input   io_rst, // @[:@60505.4]
  input   io_ctrDone, // @[:@60505.4]
  output  io_datapathEn, // @[:@60505.4]
  output  io_ctrInc, // @[:@60505.4]
  output  io_ctrRst, // @[:@60505.4]
  input   io_parentAck, // @[:@60505.4]
  input   io_backpressure, // @[:@60505.4]
  input   io_break // @[:@60505.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@60507.4]
  wire  active_reset; // @[Controllers.scala 261:22:@60507.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@60507.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@60507.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@60507.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@60507.4]
  wire  done_clock; // @[Controllers.scala 262:20:@60510.4]
  wire  done_reset; // @[Controllers.scala 262:20:@60510.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@60510.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@60510.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@60510.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@60510.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@60544.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@60544.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@60544.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@60544.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@60566.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@60566.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@60566.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@60566.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@60578.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@60578.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@60578.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@60578.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@60578.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@60586.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@60586.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@60586.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@60586.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@60586.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@60602.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@60602.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@60602.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@60602.4]
  wire  _T_80; // @[Controllers.scala 264:48:@60515.4]
  wire  _T_81; // @[Controllers.scala 264:46:@60516.4]
  wire  _T_82; // @[Controllers.scala 264:62:@60517.4]
  wire  _T_100; // @[package.scala 100:49:@60535.4]
  reg  _T_103; // @[package.scala 48:56:@60536.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@60549.4 package.scala 96:25:@60550.4]
  wire  _T_110; // @[package.scala 100:49:@60551.4]
  reg  _T_113; // @[package.scala 48:56:@60552.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@60554.4]
  wire  _T_118; // @[Controllers.scala 283:41:@60559.4]
  wire  _T_124; // @[package.scala 96:25:@60571.4 package.scala 96:25:@60572.4]
  wire  _T_126; // @[package.scala 100:49:@60573.4]
  reg  _T_129; // @[package.scala 48:56:@60574.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@60598.4]
  reg  _T_153; // @[package.scala 48:56:@60599.4]
  reg [31:0] _RAND_3;
  SRFF active ( // @[Controllers.scala 261:22:@60507.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@60510.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_671 RetimeWrapper ( // @[package.scala 93:22:@60544.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_671 RetimeWrapper_1 ( // @[package.scala 93:22:@60566.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@60578.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@60586.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_675 RetimeWrapper_4 ( // @[package.scala 93:22:@60602.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@60515.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@60516.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@60517.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@60535.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@60549.4 package.scala 96:25:@60550.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@60551.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@60554.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@60559.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@60571.4 package.scala 96:25:@60572.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@60573.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@60598.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@60577.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@60562.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@60565.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@60557.4]
  assign active_clock = clock; // @[:@60508.4]
  assign active_reset = reset; // @[:@60509.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@60520.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@60524.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@60525.4]
  assign done_clock = clock; // @[:@60511.4]
  assign done_reset = reset; // @[:@60512.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@60540.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@60533.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@60534.4]
  assign RetimeWrapper_clock = clock; // @[:@60545.4]
  assign RetimeWrapper_reset = reset; // @[:@60546.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@60547.4]
  assign RetimeWrapper_1_clock = clock; // @[:@60567.4]
  assign RetimeWrapper_1_reset = reset; // @[:@60568.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@60569.4]
  assign RetimeWrapper_2_clock = clock; // @[:@60579.4]
  assign RetimeWrapper_2_reset = reset; // @[:@60580.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@60582.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@60581.4]
  assign RetimeWrapper_3_clock = clock; // @[:@60587.4]
  assign RetimeWrapper_3_reset = reset; // @[:@60588.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@60590.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@60589.4]
  assign RetimeWrapper_4_clock = clock; // @[:@60603.4]
  assign RetimeWrapper_4_reset = reset; // @[:@60604.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@60605.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x639_inr_Foreach_iiCtr( // @[:@60615.2]
  input   clock, // @[:@60616.4]
  input   reset, // @[:@60617.4]
  input   io_input_enable, // @[:@60618.4]
  input   io_input_reset, // @[:@60618.4]
  output  io_output_issue, // @[:@60618.4]
  output  io_output_done // @[:@60618.4]
);
  reg [5:0] _T_15; // @[Counter.scala 135:22:@60620.4]
  reg [31:0] _RAND_0;
  wire  _T_17; // @[Counter.scala 138:24:@60621.4]
  wire  _T_20; // @[Counter.scala 139:23:@60623.4]
  wire [6:0] _T_26; // @[Counter.scala 141:68:@60626.4]
  wire [5:0] _T_27; // @[Counter.scala 141:68:@60627.4]
  wire [5:0] _T_28; // @[Counter.scala 141:68:@60628.4]
  wire [5:0] _T_29; // @[Counter.scala 141:23:@60629.4]
  wire [5:0] _T_30; // @[Counter.scala 142:19:@60630.4]
  wire [5:0] _T_32; // @[Counter.scala 143:15:@60631.4]
  assign _T_17 = $signed(_T_15) == $signed(6'she); // @[Counter.scala 138:24:@60621.4]
  assign _T_20 = $signed(_T_15) == $signed(6'sh0); // @[Counter.scala 139:23:@60623.4]
  assign _T_26 = $signed(_T_15) - $signed(6'sh1); // @[Counter.scala 141:68:@60626.4]
  assign _T_27 = $signed(_T_15) - $signed(6'sh1); // @[Counter.scala 141:68:@60627.4]
  assign _T_28 = $signed(_T_27); // @[Counter.scala 141:68:@60628.4]
  assign _T_29 = _T_20 ? $signed(6'she) : $signed(_T_28); // @[Counter.scala 141:23:@60629.4]
  assign _T_30 = io_input_enable ? $signed(_T_29) : $signed(_T_15); // @[Counter.scala 142:19:@60630.4]
  assign _T_32 = io_input_reset ? $signed(6'she) : $signed(_T_30); // @[Counter.scala 143:15:@60631.4]
  assign io_output_issue = _T_17 & io_input_enable; // @[Counter.scala 146:21:@60634.4]
  assign io_output_done = _T_20 & io_input_enable; // @[Counter.scala 145:20:@60633.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 6'she;
    end else begin
      if (io_input_reset) begin
        _T_15 <= 6'she;
      end else begin
        if (io_input_enable) begin
          if (_T_20) begin
            _T_15 <= 6'she;
          end else begin
            _T_15 <= _T_28;
          end
        end
      end
    end
  end
endmodule
module RetimeWrapper_689( // @[:@61285.2]
  input         clock, // @[:@61286.4]
  input         reset, // @[:@61287.4]
  input  [31:0] io_in, // @[:@61288.4]
  output [31:0] io_out // @[:@61288.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@61290.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@61290.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@61290.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@61290.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@61290.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@61290.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(14)) sr ( // @[RetimeShiftRegister.scala 15:20:@61290.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@61303.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@61302.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@61301.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@61300.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@61299.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@61297.4]
endmodule
module x639_inr_Foreach_kernelx639_inr_Foreach_concrete1( // @[:@61721.2]
  input         clock, // @[:@61722.4]
  input         reset, // @[:@61723.4]
  output [1:0]  io_in_x555_tmp_1_wPort_1_ofs_0, // @[:@61724.4]
  output [31:0] io_in_x555_tmp_1_wPort_1_data_0, // @[:@61724.4]
  output        io_in_x555_tmp_1_wPort_1_en_0, // @[:@61724.4]
  output        io_in_x555_tmp_1_sEn_5, // @[:@61724.4]
  output        io_in_x555_tmp_1_sDone_5, // @[:@61724.4]
  output [1:0]  io_in_x554_tmp_0_wPort_1_ofs_0, // @[:@61724.4]
  output [31:0] io_in_x554_tmp_0_wPort_1_data_0, // @[:@61724.4]
  output        io_in_x554_tmp_0_wPort_1_en_0, // @[:@61724.4]
  output        io_in_x554_tmp_0_sEn_5, // @[:@61724.4]
  output        io_in_x554_tmp_0_sDone_5, // @[:@61724.4]
  output [1:0]  io_in_x558_tmp_4_wPort_1_ofs_0, // @[:@61724.4]
  output [31:0] io_in_x558_tmp_4_wPort_1_data_0, // @[:@61724.4]
  output        io_in_x558_tmp_4_wPort_1_en_0, // @[:@61724.4]
  output        io_in_x558_tmp_4_sEn_5, // @[:@61724.4]
  output        io_in_x558_tmp_4_sDone_5, // @[:@61724.4]
  input         io_in_b552, // @[:@61724.4]
  output        io_in_x594_force_0_rPort_0_en_0, // @[:@61724.4]
  input  [31:0] io_in_x594_force_0_rPort_0_output_0, // @[:@61724.4]
  output        io_in_x594_force_0_sEn_1, // @[:@61724.4]
  output        io_in_x594_force_0_sDone_1, // @[:@61724.4]
  output [1:0]  io_in_x557_tmp_3_rPort_0_ofs_0, // @[:@61724.4]
  output        io_in_x557_tmp_3_rPort_0_en_0, // @[:@61724.4]
  input  [31:0] io_in_x557_tmp_3_rPort_0_output_0, // @[:@61724.4]
  output [1:0]  io_in_x557_tmp_3_wPort_1_ofs_0, // @[:@61724.4]
  output [31:0] io_in_x557_tmp_3_wPort_1_data_0, // @[:@61724.4]
  output        io_in_x557_tmp_3_wPort_1_en_0, // @[:@61724.4]
  output        io_in_x557_tmp_3_sEn_5, // @[:@61724.4]
  output        io_in_x557_tmp_3_sDone_5, // @[:@61724.4]
  output [1:0]  io_in_x556_tmp_2_wPort_1_ofs_0, // @[:@61724.4]
  output [31:0] io_in_x556_tmp_2_wPort_1_data_0, // @[:@61724.4]
  output        io_in_x556_tmp_2_wPort_1_en_0, // @[:@61724.4]
  output        io_in_x556_tmp_2_sEn_5, // @[:@61724.4]
  output        io_in_x556_tmp_2_sDone_5, // @[:@61724.4]
  input         io_in_b543, // @[:@61724.4]
  output [63:0] io_in_instrctrs_15_cycs, // @[:@61724.4]
  output [63:0] io_in_instrctrs_15_iters, // @[:@61724.4]
  input         io_sigsIn_done, // @[:@61724.4]
  input         io_sigsIn_iiIssue, // @[:@61724.4]
  input         io_sigsIn_datapathEn, // @[:@61724.4]
  input         io_sigsIn_baseEn, // @[:@61724.4]
  input         io_sigsIn_break, // @[:@61724.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@61724.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@61724.4]
  input         io_rr // @[:@61724.4]
);
  wire  cycles_x639_inr_Foreach_clock; // @[sm_x639_inr_Foreach.scala 87:43:@62073.4]
  wire  cycles_x639_inr_Foreach_reset; // @[sm_x639_inr_Foreach.scala 87:43:@62073.4]
  wire  cycles_x639_inr_Foreach_io_enable; // @[sm_x639_inr_Foreach.scala 87:43:@62073.4]
  wire [63:0] cycles_x639_inr_Foreach_io_count; // @[sm_x639_inr_Foreach.scala 87:43:@62073.4]
  wire  iters_x639_inr_Foreach_clock; // @[sm_x639_inr_Foreach.scala 88:42:@62076.4]
  wire  iters_x639_inr_Foreach_reset; // @[sm_x639_inr_Foreach.scala 88:42:@62076.4]
  wire  iters_x639_inr_Foreach_io_enable; // @[sm_x639_inr_Foreach.scala 88:42:@62076.4]
  wire [63:0] iters_x639_inr_Foreach_io_count; // @[sm_x639_inr_Foreach.scala 88:42:@62076.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@62093.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@62093.4]
  wire  x630_mul_1_clock; // @[Math.scala 262:24:@62127.4]
  wire  x630_mul_1_reset; // @[Math.scala 262:24:@62127.4]
  wire [31:0] x630_mul_1_io_a; // @[Math.scala 262:24:@62127.4]
  wire [31:0] x630_mul_1_io_b; // @[Math.scala 262:24:@62127.4]
  wire  x630_mul_1_io_flow; // @[Math.scala 262:24:@62127.4]
  wire [31:0] x630_mul_1_io_result; // @[Math.scala 262:24:@62127.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@62162.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@62162.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@62162.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@62162.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@62162.4]
  wire  x633_mul_1_clock; // @[Math.scala 262:24:@62171.4]
  wire  x633_mul_1_reset; // @[Math.scala 262:24:@62171.4]
  wire [31:0] x633_mul_1_io_a; // @[Math.scala 262:24:@62171.4]
  wire [31:0] x633_mul_1_io_b; // @[Math.scala 262:24:@62171.4]
  wire  x633_mul_1_io_flow; // @[Math.scala 262:24:@62171.4]
  wire [31:0] x633_mul_1_io_result; // @[Math.scala 262:24:@62171.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@62182.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@62182.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@62182.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@62182.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@62192.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@62192.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@62192.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@62192.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@62202.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@62202.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@62202.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@62202.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@62212.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@62212.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@62212.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@62212.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@62226.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@62226.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@62226.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@62226.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@62252.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@62252.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@62252.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@62252.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@62278.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@62278.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@62278.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@62278.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@62304.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@62304.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@62304.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@62304.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@62330.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@62330.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@62330.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@62330.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@62351.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@62351.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@62351.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@62351.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@62351.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@62362.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@62362.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@62362.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@62362.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@62362.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@62373.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@62373.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@62373.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@62373.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@62373.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@62384.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@62384.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@62384.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@62384.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@62384.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@62395.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@62395.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@62395.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@62395.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@62395.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@62406.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@62406.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@62406.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@62406.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@62406.4]
  wire  _T_1768; // @[package.scala 100:49:@62080.4]
  reg  _T_1771; // @[package.scala 48:56:@62081.4]
  reg [31:0] _RAND_0;
  wire  b627; // @[sm_x639_inr_Foreach.scala 93:18:@62101.4]
  wire  _T_1796; // @[sm_x639_inr_Foreach.scala 98:114:@62107.4]
  wire  _T_1797; // @[sm_x639_inr_Foreach.scala 98:111:@62108.4]
  wire  _T_1798; // @[sm_x639_inr_Foreach.scala 98:156:@62109.4]
  wire  _T_1802; // @[implicits.scala 56:10:@62111.4]
  wire  _T_1803; // @[sm_x639_inr_Foreach.scala 98:131:@62112.4]
  wire  _T_1804; // @[sm_x639_inr_Foreach.scala 98:228:@62113.4]
  wire  _T_1805; // @[sm_x639_inr_Foreach.scala 98:236:@62114.4]
  wire  _T_1885; // @[package.scala 96:25:@62231.4 package.scala 96:25:@62232.4]
  wire  _T_1887; // @[implicits.scala 56:10:@62233.4]
  wire  _T_1888; // @[sm_x639_inr_Foreach.scala 130:115:@62234.4]
  wire  _T_1890; // @[sm_x639_inr_Foreach.scala 130:213:@62236.4]
  wire  x787_b627_D14; // @[package.scala 96:25:@62207.4 package.scala 96:25:@62208.4]
  wire  _T_1892; // @[sm_x639_inr_Foreach.scala 130:258:@62238.4]
  wire  x785_b552_D14; // @[package.scala 96:25:@62187.4 package.scala 96:25:@62188.4]
  wire  _T_1893; // @[sm_x639_inr_Foreach.scala 130:266:@62239.4]
  wire  x788_b543_D14; // @[package.scala 96:25:@62217.4 package.scala 96:25:@62218.4]
  wire  _T_1905; // @[package.scala 96:25:@62257.4 package.scala 96:25:@62258.4]
  wire  _T_1907; // @[implicits.scala 56:10:@62259.4]
  wire  _T_1908; // @[sm_x639_inr_Foreach.scala 135:115:@62260.4]
  wire  _T_1910; // @[sm_x639_inr_Foreach.scala 135:213:@62262.4]
  wire  _T_1912; // @[sm_x639_inr_Foreach.scala 135:258:@62264.4]
  wire  _T_1913; // @[sm_x639_inr_Foreach.scala 135:266:@62265.4]
  wire  _T_1925; // @[package.scala 96:25:@62283.4 package.scala 96:25:@62284.4]
  wire  _T_1927; // @[implicits.scala 56:10:@62285.4]
  wire  _T_1928; // @[sm_x639_inr_Foreach.scala 140:115:@62286.4]
  wire  _T_1930; // @[sm_x639_inr_Foreach.scala 140:213:@62288.4]
  wire  _T_1932; // @[sm_x639_inr_Foreach.scala 140:258:@62290.4]
  wire  _T_1933; // @[sm_x639_inr_Foreach.scala 140:266:@62291.4]
  wire  _T_1945; // @[package.scala 96:25:@62309.4 package.scala 96:25:@62310.4]
  wire  _T_1947; // @[implicits.scala 56:10:@62311.4]
  wire  _T_1948; // @[sm_x639_inr_Foreach.scala 145:115:@62312.4]
  wire  _T_1950; // @[sm_x639_inr_Foreach.scala 145:213:@62314.4]
  wire  _T_1952; // @[sm_x639_inr_Foreach.scala 145:258:@62316.4]
  wire  _T_1953; // @[sm_x639_inr_Foreach.scala 145:266:@62317.4]
  wire  _T_1965; // @[package.scala 96:25:@62335.4 package.scala 96:25:@62336.4]
  wire  _T_1967; // @[implicits.scala 56:10:@62337.4]
  wire  _T_1968; // @[sm_x639_inr_Foreach.scala 150:115:@62338.4]
  wire  _T_1970; // @[sm_x639_inr_Foreach.scala 150:213:@62340.4]
  wire  _T_1972; // @[sm_x639_inr_Foreach.scala 150:258:@62342.4]
  wire  _T_1973; // @[sm_x639_inr_Foreach.scala 150:266:@62343.4]
  wire  _T_1978; // @[package.scala 96:25:@62356.4 package.scala 96:25:@62357.4]
  wire  _T_1984; // @[package.scala 96:25:@62367.4 package.scala 96:25:@62368.4]
  wire  _T_1990; // @[package.scala 96:25:@62378.4 package.scala 96:25:@62379.4]
  wire  _T_1996; // @[package.scala 96:25:@62389.4 package.scala 96:25:@62390.4]
  wire  _T_2002; // @[package.scala 96:25:@62400.4 package.scala 96:25:@62401.4]
  wire  _T_2008; // @[package.scala 96:25:@62411.4 package.scala 96:25:@62412.4]
  wire [31:0] b626_number; // @[Math.scala 723:22:@62098.4 Math.scala 724:14:@62099.4]
  wire [31:0] x786_b626_D14_number; // @[package.scala 96:25:@62197.4 package.scala 96:25:@62198.4]
  InstrumentationCounter cycles_x639_inr_Foreach ( // @[sm_x639_inr_Foreach.scala 87:43:@62073.4]
    .clock(cycles_x639_inr_Foreach_clock),
    .reset(cycles_x639_inr_Foreach_reset),
    .io_enable(cycles_x639_inr_Foreach_io_enable),
    .io_count(cycles_x639_inr_Foreach_io_count)
  );
  InstrumentationCounter iters_x639_inr_Foreach ( // @[sm_x639_inr_Foreach.scala 88:42:@62076.4]
    .clock(iters_x639_inr_Foreach_clock),
    .reset(iters_x639_inr_Foreach_reset),
    .io_enable(iters_x639_inr_Foreach_io_enable),
    .io_count(iters_x639_inr_Foreach_io_count)
  );
  _ _ ( // @[Math.scala 720:24:@62093.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x586_mul x630_mul_1 ( // @[Math.scala 262:24:@62127.4]
    .clock(x630_mul_1_clock),
    .reset(x630_mul_1_reset),
    .io_a(x630_mul_1_io_a),
    .io_b(x630_mul_1_io_b),
    .io_flow(x630_mul_1_io_flow),
    .io_result(x630_mul_1_io_result)
  );
  RetimeWrapper_529 RetimeWrapper ( // @[package.scala 93:22:@62162.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x586_mul x633_mul_1 ( // @[Math.scala 262:24:@62171.4]
    .clock(x633_mul_1_clock),
    .reset(x633_mul_1_reset),
    .io_a(x633_mul_1_io_a),
    .io_b(x633_mul_1_io_b),
    .io_flow(x633_mul_1_io_flow),
    .io_result(x633_mul_1_io_result)
  );
  RetimeWrapper_675 RetimeWrapper_1 ( // @[package.scala 93:22:@62182.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_689 RetimeWrapper_2 ( // @[package.scala 93:22:@62192.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_675 RetimeWrapper_3 ( // @[package.scala 93:22:@62202.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_675 RetimeWrapper_4 ( // @[package.scala 93:22:@62212.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_675 RetimeWrapper_5 ( // @[package.scala 93:22:@62226.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_675 RetimeWrapper_6 ( // @[package.scala 93:22:@62252.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_675 RetimeWrapper_7 ( // @[package.scala 93:22:@62278.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_675 RetimeWrapper_8 ( // @[package.scala 93:22:@62304.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_675 RetimeWrapper_9 ( // @[package.scala 93:22:@62330.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@62351.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 ( // @[package.scala 93:22:@62362.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper RetimeWrapper_12 ( // @[package.scala 93:22:@62373.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 ( // @[package.scala 93:22:@62384.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@62395.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@62406.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  assign _T_1768 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@62080.4]
  assign b627 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x639_inr_Foreach.scala 93:18:@62101.4]
  assign _T_1796 = ~ io_sigsIn_break; // @[sm_x639_inr_Foreach.scala 98:114:@62107.4]
  assign _T_1797 = io_rr & _T_1796; // @[sm_x639_inr_Foreach.scala 98:111:@62108.4]
  assign _T_1798 = io_sigsIn_datapathEn & io_sigsIn_iiIssue; // @[sm_x639_inr_Foreach.scala 98:156:@62109.4]
  assign _T_1802 = io_rr ? _T_1798 : 1'h0; // @[implicits.scala 56:10:@62111.4]
  assign _T_1803 = _T_1797 & _T_1802; // @[sm_x639_inr_Foreach.scala 98:131:@62112.4]
  assign _T_1804 = _T_1803 & b627; // @[sm_x639_inr_Foreach.scala 98:228:@62113.4]
  assign _T_1805 = _T_1804 & io_in_b552; // @[sm_x639_inr_Foreach.scala 98:236:@62114.4]
  assign _T_1885 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@62231.4 package.scala 96:25:@62232.4]
  assign _T_1887 = io_rr ? _T_1885 : 1'h0; // @[implicits.scala 56:10:@62233.4]
  assign _T_1888 = _T_1796 & _T_1887; // @[sm_x639_inr_Foreach.scala 130:115:@62234.4]
  assign _T_1890 = _T_1888 & _T_1796; // @[sm_x639_inr_Foreach.scala 130:213:@62236.4]
  assign x787_b627_D14 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@62207.4 package.scala 96:25:@62208.4]
  assign _T_1892 = _T_1890 & x787_b627_D14; // @[sm_x639_inr_Foreach.scala 130:258:@62238.4]
  assign x785_b552_D14 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@62187.4 package.scala 96:25:@62188.4]
  assign _T_1893 = _T_1892 & x785_b552_D14; // @[sm_x639_inr_Foreach.scala 130:266:@62239.4]
  assign x788_b543_D14 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@62217.4 package.scala 96:25:@62218.4]
  assign _T_1905 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@62257.4 package.scala 96:25:@62258.4]
  assign _T_1907 = io_rr ? _T_1905 : 1'h0; // @[implicits.scala 56:10:@62259.4]
  assign _T_1908 = _T_1796 & _T_1907; // @[sm_x639_inr_Foreach.scala 135:115:@62260.4]
  assign _T_1910 = _T_1908 & _T_1796; // @[sm_x639_inr_Foreach.scala 135:213:@62262.4]
  assign _T_1912 = _T_1910 & x787_b627_D14; // @[sm_x639_inr_Foreach.scala 135:258:@62264.4]
  assign _T_1913 = _T_1912 & x785_b552_D14; // @[sm_x639_inr_Foreach.scala 135:266:@62265.4]
  assign _T_1925 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@62283.4 package.scala 96:25:@62284.4]
  assign _T_1927 = io_rr ? _T_1925 : 1'h0; // @[implicits.scala 56:10:@62285.4]
  assign _T_1928 = _T_1796 & _T_1927; // @[sm_x639_inr_Foreach.scala 140:115:@62286.4]
  assign _T_1930 = _T_1928 & _T_1796; // @[sm_x639_inr_Foreach.scala 140:213:@62288.4]
  assign _T_1932 = _T_1930 & x787_b627_D14; // @[sm_x639_inr_Foreach.scala 140:258:@62290.4]
  assign _T_1933 = _T_1932 & x785_b552_D14; // @[sm_x639_inr_Foreach.scala 140:266:@62291.4]
  assign _T_1945 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@62309.4 package.scala 96:25:@62310.4]
  assign _T_1947 = io_rr ? _T_1945 : 1'h0; // @[implicits.scala 56:10:@62311.4]
  assign _T_1948 = _T_1796 & _T_1947; // @[sm_x639_inr_Foreach.scala 145:115:@62312.4]
  assign _T_1950 = _T_1948 & _T_1796; // @[sm_x639_inr_Foreach.scala 145:213:@62314.4]
  assign _T_1952 = _T_1950 & x787_b627_D14; // @[sm_x639_inr_Foreach.scala 145:258:@62316.4]
  assign _T_1953 = _T_1952 & x785_b552_D14; // @[sm_x639_inr_Foreach.scala 145:266:@62317.4]
  assign _T_1965 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@62335.4 package.scala 96:25:@62336.4]
  assign _T_1967 = io_rr ? _T_1965 : 1'h0; // @[implicits.scala 56:10:@62337.4]
  assign _T_1968 = _T_1796 & _T_1967; // @[sm_x639_inr_Foreach.scala 150:115:@62338.4]
  assign _T_1970 = _T_1968 & _T_1796; // @[sm_x639_inr_Foreach.scala 150:213:@62340.4]
  assign _T_1972 = _T_1970 & x787_b627_D14; // @[sm_x639_inr_Foreach.scala 150:258:@62342.4]
  assign _T_1973 = _T_1972 & x785_b552_D14; // @[sm_x639_inr_Foreach.scala 150:266:@62343.4]
  assign _T_1978 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@62356.4 package.scala 96:25:@62357.4]
  assign _T_1984 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@62367.4 package.scala 96:25:@62368.4]
  assign _T_1990 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@62378.4 package.scala 96:25:@62379.4]
  assign _T_1996 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@62389.4 package.scala 96:25:@62390.4]
  assign _T_2002 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@62400.4 package.scala 96:25:@62401.4]
  assign _T_2008 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@62411.4 package.scala 96:25:@62412.4]
  assign b626_number = __io_result; // @[Math.scala 723:22:@62098.4 Math.scala 724:14:@62099.4]
  assign x786_b626_D14_number = RetimeWrapper_2_io_out; // @[package.scala 96:25:@62197.4 package.scala 96:25:@62198.4]
  assign io_in_x555_tmp_1_wPort_1_ofs_0 = x786_b626_D14_number[1:0]; // @[MemInterfaceType.scala 89:54:@62242.4]
  assign io_in_x555_tmp_1_wPort_1_data_0 = x633_mul_1_io_result; // @[MemInterfaceType.scala 90:56:@62243.4]
  assign io_in_x555_tmp_1_wPort_1_en_0 = _T_1893 & x788_b543_D14; // @[MemInterfaceType.scala 93:57:@62245.4]
  assign io_in_x555_tmp_1_sEn_5 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@62370.4]
  assign io_in_x555_tmp_1_sDone_5 = io_rr ? _T_1984 : 1'h0; // @[MemInterfaceType.scala 197:17:@62371.4]
  assign io_in_x554_tmp_0_wPort_1_ofs_0 = x786_b626_D14_number[1:0]; // @[MemInterfaceType.scala 89:54:@62268.4]
  assign io_in_x554_tmp_0_wPort_1_data_0 = x633_mul_1_io_result; // @[MemInterfaceType.scala 90:56:@62269.4]
  assign io_in_x554_tmp_0_wPort_1_en_0 = _T_1913 & x788_b543_D14; // @[MemInterfaceType.scala 93:57:@62271.4]
  assign io_in_x554_tmp_0_sEn_5 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@62359.4]
  assign io_in_x554_tmp_0_sDone_5 = io_rr ? _T_1978 : 1'h0; // @[MemInterfaceType.scala 197:17:@62360.4]
  assign io_in_x558_tmp_4_wPort_1_ofs_0 = x786_b626_D14_number[1:0]; // @[MemInterfaceType.scala 89:54:@62294.4]
  assign io_in_x558_tmp_4_wPort_1_data_0 = x633_mul_1_io_result; // @[MemInterfaceType.scala 90:56:@62295.4]
  assign io_in_x558_tmp_4_wPort_1_en_0 = _T_1933 & x788_b543_D14; // @[MemInterfaceType.scala 93:57:@62297.4]
  assign io_in_x558_tmp_4_sEn_5 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@62403.4]
  assign io_in_x558_tmp_4_sDone_5 = io_rr ? _T_2002 : 1'h0; // @[MemInterfaceType.scala 197:17:@62404.4]
  assign io_in_x594_force_0_rPort_0_en_0 = _T_1805 & io_in_b543; // @[MemInterfaceType.scala 110:79:@62156.4]
  assign io_in_x594_force_0_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@62414.4]
  assign io_in_x594_force_0_sDone_1 = io_rr ? _T_2008 : 1'h0; // @[MemInterfaceType.scala 197:17:@62415.4]
  assign io_in_x557_tmp_3_rPort_0_ofs_0 = b626_number[1:0]; // @[MemInterfaceType.scala 107:54:@62118.4]
  assign io_in_x557_tmp_3_rPort_0_en_0 = _T_1805 & io_in_b543; // @[MemInterfaceType.scala 110:79:@62120.4]
  assign io_in_x557_tmp_3_wPort_1_ofs_0 = x786_b626_D14_number[1:0]; // @[MemInterfaceType.scala 89:54:@62320.4]
  assign io_in_x557_tmp_3_wPort_1_data_0 = x633_mul_1_io_result; // @[MemInterfaceType.scala 90:56:@62321.4]
  assign io_in_x557_tmp_3_wPort_1_en_0 = _T_1953 & x788_b543_D14; // @[MemInterfaceType.scala 93:57:@62323.4]
  assign io_in_x557_tmp_3_sEn_5 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@62392.4]
  assign io_in_x557_tmp_3_sDone_5 = io_rr ? _T_1996 : 1'h0; // @[MemInterfaceType.scala 197:17:@62393.4]
  assign io_in_x556_tmp_2_wPort_1_ofs_0 = x786_b626_D14_number[1:0]; // @[MemInterfaceType.scala 89:54:@62346.4]
  assign io_in_x556_tmp_2_wPort_1_data_0 = x633_mul_1_io_result; // @[MemInterfaceType.scala 90:56:@62347.4]
  assign io_in_x556_tmp_2_wPort_1_en_0 = _T_1973 & x788_b543_D14; // @[MemInterfaceType.scala 93:57:@62349.4]
  assign io_in_x556_tmp_2_sEn_5 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@62381.4]
  assign io_in_x556_tmp_2_sDone_5 = io_rr ? _T_1990 : 1'h0; // @[MemInterfaceType.scala 197:17:@62382.4]
  assign io_in_instrctrs_15_cycs = cycles_x639_inr_Foreach_io_count; // @[Ledger.scala 293:21:@62085.4]
  assign io_in_instrctrs_15_iters = iters_x639_inr_Foreach_io_count; // @[Ledger.scala 294:22:@62086.4]
  assign cycles_x639_inr_Foreach_clock = clock; // @[:@62074.4]
  assign cycles_x639_inr_Foreach_reset = reset; // @[:@62075.4]
  assign cycles_x639_inr_Foreach_io_enable = io_sigsIn_baseEn; // @[sm_x639_inr_Foreach.scala 89:41:@62079.4]
  assign iters_x639_inr_Foreach_clock = clock; // @[:@62077.4]
  assign iters_x639_inr_Foreach_reset = reset; // @[:@62078.4]
  assign iters_x639_inr_Foreach_io_enable = io_sigsIn_done & _T_1771; // @[sm_x639_inr_Foreach.scala 90:40:@62084.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@62096.4]
  assign x630_mul_1_clock = clock; // @[:@62128.4]
  assign x630_mul_1_reset = reset; // @[:@62129.4]
  assign x630_mul_1_io_a = io_in_x557_tmp_3_rPort_0_output_0; // @[Math.scala 263:17:@62130.4]
  assign x630_mul_1_io_b = 32'h66666; // @[Math.scala 264:17:@62131.4]
  assign x630_mul_1_io_flow = 1'h1; // @[Math.scala 265:20:@62132.4]
  assign RetimeWrapper_clock = clock; // @[:@62163.4]
  assign RetimeWrapper_reset = reset; // @[:@62164.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@62166.4]
  assign RetimeWrapper_io_in = io_in_x594_force_0_rPort_0_output_0; // @[package.scala 94:16:@62165.4]
  assign x633_mul_1_clock = clock; // @[:@62172.4]
  assign x633_mul_1_reset = reset; // @[:@62173.4]
  assign x633_mul_1_io_a = x630_mul_1_io_result; // @[Math.scala 263:17:@62174.4]
  assign x633_mul_1_io_b = RetimeWrapper_io_out; // @[Math.scala 264:17:@62175.4]
  assign x633_mul_1_io_flow = 1'h1; // @[Math.scala 265:20:@62176.4]
  assign RetimeWrapper_1_clock = clock; // @[:@62183.4]
  assign RetimeWrapper_1_reset = reset; // @[:@62184.4]
  assign RetimeWrapper_1_io_in = io_in_b552; // @[package.scala 94:16:@62185.4]
  assign RetimeWrapper_2_clock = clock; // @[:@62193.4]
  assign RetimeWrapper_2_reset = reset; // @[:@62194.4]
  assign RetimeWrapper_2_io_in = __io_result; // @[package.scala 94:16:@62195.4]
  assign RetimeWrapper_3_clock = clock; // @[:@62203.4]
  assign RetimeWrapper_3_reset = reset; // @[:@62204.4]
  assign RetimeWrapper_3_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@62205.4]
  assign RetimeWrapper_4_clock = clock; // @[:@62213.4]
  assign RetimeWrapper_4_reset = reset; // @[:@62214.4]
  assign RetimeWrapper_4_io_in = io_in_b543; // @[package.scala 94:16:@62215.4]
  assign RetimeWrapper_5_clock = clock; // @[:@62227.4]
  assign RetimeWrapper_5_reset = reset; // @[:@62228.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_datapathEn & io_sigsIn_iiIssue; // @[package.scala 94:16:@62229.4]
  assign RetimeWrapper_6_clock = clock; // @[:@62253.4]
  assign RetimeWrapper_6_reset = reset; // @[:@62254.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn & io_sigsIn_iiIssue; // @[package.scala 94:16:@62255.4]
  assign RetimeWrapper_7_clock = clock; // @[:@62279.4]
  assign RetimeWrapper_7_reset = reset; // @[:@62280.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_datapathEn & io_sigsIn_iiIssue; // @[package.scala 94:16:@62281.4]
  assign RetimeWrapper_8_clock = clock; // @[:@62305.4]
  assign RetimeWrapper_8_reset = reset; // @[:@62306.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_datapathEn & io_sigsIn_iiIssue; // @[package.scala 94:16:@62307.4]
  assign RetimeWrapper_9_clock = clock; // @[:@62331.4]
  assign RetimeWrapper_9_reset = reset; // @[:@62332.4]
  assign RetimeWrapper_9_io_in = io_sigsIn_datapathEn & io_sigsIn_iiIssue; // @[package.scala 94:16:@62333.4]
  assign RetimeWrapper_10_clock = clock; // @[:@62352.4]
  assign RetimeWrapper_10_reset = reset; // @[:@62353.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@62355.4]
  assign RetimeWrapper_10_io_in = io_sigsIn_done; // @[package.scala 94:16:@62354.4]
  assign RetimeWrapper_11_clock = clock; // @[:@62363.4]
  assign RetimeWrapper_11_reset = reset; // @[:@62364.4]
  assign RetimeWrapper_11_io_flow = 1'h1; // @[package.scala 95:18:@62366.4]
  assign RetimeWrapper_11_io_in = io_sigsIn_done; // @[package.scala 94:16:@62365.4]
  assign RetimeWrapper_12_clock = clock; // @[:@62374.4]
  assign RetimeWrapper_12_reset = reset; // @[:@62375.4]
  assign RetimeWrapper_12_io_flow = 1'h1; // @[package.scala 95:18:@62377.4]
  assign RetimeWrapper_12_io_in = io_sigsIn_done; // @[package.scala 94:16:@62376.4]
  assign RetimeWrapper_13_clock = clock; // @[:@62385.4]
  assign RetimeWrapper_13_reset = reset; // @[:@62386.4]
  assign RetimeWrapper_13_io_flow = 1'h1; // @[package.scala 95:18:@62388.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_done; // @[package.scala 94:16:@62387.4]
  assign RetimeWrapper_14_clock = clock; // @[:@62396.4]
  assign RetimeWrapper_14_reset = reset; // @[:@62397.4]
  assign RetimeWrapper_14_io_flow = 1'h1; // @[package.scala 95:18:@62399.4]
  assign RetimeWrapper_14_io_in = io_sigsIn_done; // @[package.scala 94:16:@62398.4]
  assign RetimeWrapper_15_clock = clock; // @[:@62407.4]
  assign RetimeWrapper_15_reset = reset; // @[:@62408.4]
  assign RetimeWrapper_15_io_flow = 1'h1; // @[package.scala 95:18:@62410.4]
  assign RetimeWrapper_15_io_in = io_sigsIn_done; // @[package.scala 94:16:@62409.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1771 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1771 <= 1'h0;
    end else begin
      _T_1771 <= _T_1768;
    end
  end
endmodule
module x652_inr_Foreach_sm( // @[:@62603.2]
  input   clock, // @[:@62604.4]
  input   reset, // @[:@62605.4]
  input   io_enable, // @[:@62606.4]
  output  io_done, // @[:@62606.4]
  output  io_doneLatch, // @[:@62606.4]
  input   io_ctrDone, // @[:@62606.4]
  output  io_datapathEn, // @[:@62606.4]
  output  io_ctrInc, // @[:@62606.4]
  output  io_ctrRst, // @[:@62606.4]
  input   io_parentAck, // @[:@62606.4]
  input   io_backpressure, // @[:@62606.4]
  input   io_break // @[:@62606.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@62608.4]
  wire  active_reset; // @[Controllers.scala 261:22:@62608.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@62608.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@62608.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@62608.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@62608.4]
  wire  done_clock; // @[Controllers.scala 262:20:@62611.4]
  wire  done_reset; // @[Controllers.scala 262:20:@62611.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@62611.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@62611.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@62611.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@62611.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@62645.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@62645.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@62645.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@62645.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@62645.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@62667.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@62667.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@62667.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@62667.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@62667.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@62679.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@62679.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@62679.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@62679.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@62679.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@62687.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@62687.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@62687.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@62687.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@62687.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@62703.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@62703.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@62703.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@62703.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@62703.4]
  wire  _T_80; // @[Controllers.scala 264:48:@62616.4]
  wire  _T_81; // @[Controllers.scala 264:46:@62617.4]
  wire  _T_82; // @[Controllers.scala 264:62:@62618.4]
  wire  _T_83; // @[Controllers.scala 264:60:@62619.4]
  wire  _T_100; // @[package.scala 100:49:@62636.4]
  reg  _T_103; // @[package.scala 48:56:@62637.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@62650.4 package.scala 96:25:@62651.4]
  wire  _T_110; // @[package.scala 100:49:@62652.4]
  reg  _T_113; // @[package.scala 48:56:@62653.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@62655.4]
  wire  _T_118; // @[Controllers.scala 283:41:@62660.4]
  wire  _T_119; // @[Controllers.scala 283:59:@62661.4]
  wire  _T_121; // @[Controllers.scala 284:37:@62664.4]
  wire  _T_124; // @[package.scala 96:25:@62672.4 package.scala 96:25:@62673.4]
  wire  _T_126; // @[package.scala 100:49:@62674.4]
  reg  _T_129; // @[package.scala 48:56:@62675.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@62697.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@62699.4]
  reg  _T_153; // @[package.scala 48:56:@62700.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@62708.4 package.scala 96:25:@62709.4]
  wire  _T_158; // @[Controllers.scala 292:61:@62710.4]
  wire  _T_159; // @[Controllers.scala 292:24:@62711.4]
  SRFF active ( // @[Controllers.scala 261:22:@62608.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@62611.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_25 RetimeWrapper ( // @[package.scala 93:22:@62645.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@62667.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@62679.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@62687.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_59 RetimeWrapper_4 ( // @[package.scala 93:22:@62703.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@62616.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@62617.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@62618.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@62619.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@62636.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@62650.4 package.scala 96:25:@62651.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@62652.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@62655.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@62660.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@62661.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@62664.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@62672.4 package.scala 96:25:@62673.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@62674.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@62699.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@62708.4 package.scala 96:25:@62709.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@62710.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@62711.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@62678.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@62713.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@62663.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@62666.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@62658.4]
  assign active_clock = clock; // @[:@62609.4]
  assign active_reset = reset; // @[:@62610.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@62621.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@62625.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@62626.4]
  assign done_clock = clock; // @[:@62612.4]
  assign done_reset = reset; // @[:@62613.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@62641.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@62634.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@62635.4]
  assign RetimeWrapper_clock = clock; // @[:@62646.4]
  assign RetimeWrapper_reset = reset; // @[:@62647.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@62649.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@62648.4]
  assign RetimeWrapper_1_clock = clock; // @[:@62668.4]
  assign RetimeWrapper_1_reset = reset; // @[:@62669.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@62671.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@62670.4]
  assign RetimeWrapper_2_clock = clock; // @[:@62680.4]
  assign RetimeWrapper_2_reset = reset; // @[:@62681.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@62683.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@62682.4]
  assign RetimeWrapper_3_clock = clock; // @[:@62688.4]
  assign RetimeWrapper_3_reset = reset; // @[:@62689.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@62691.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@62690.4]
  assign RetimeWrapper_4_clock = clock; // @[:@62704.4]
  assign RetimeWrapper_4_reset = reset; // @[:@62705.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@62707.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@62706.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x648_sum( // @[:@63095.2]
  input         clock, // @[:@63096.4]
  input         reset, // @[:@63097.4]
  input  [31:0] io_a, // @[:@63098.4]
  input  [31:0] io_b, // @[:@63098.4]
  output [31:0] io_result // @[:@63098.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@63106.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@63106.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@63113.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@63113.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@63131.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@63131.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@63131.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@63131.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@63131.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@63111.4 Math.scala 724:14:@63112.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@63118.4 Math.scala 724:14:@63119.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@63120.4]
  __37 _ ( // @[Math.scala 720:24:@63106.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __37 __1 ( // @[Math.scala 720:24:@63113.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_12 fix2fixBox ( // @[Math.scala 141:30:@63131.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@63111.4 Math.scala 724:14:@63112.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@63118.4 Math.scala 724:14:@63119.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@63120.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@63139.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@63109.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@63116.4]
  assign fix2fixBox_clock = clock; // @[:@63132.4]
  assign fix2fixBox_reset = reset; // @[:@63133.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@63134.4]
  assign fix2fixBox_io_flow = 1'h1; // @[Math.scala 145:26:@63137.4]
endmodule
module RetimeWrapper_718( // @[:@63281.2]
  input         clock, // @[:@63282.4]
  input         reset, // @[:@63283.4]
  input  [31:0] io_in, // @[:@63284.4]
  output [31:0] io_out // @[:@63284.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@63286.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@63286.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@63286.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@63286.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@63286.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@63286.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@63286.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@63299.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@63298.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@63297.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@63296.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@63295.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@63293.4]
endmodule
module x652_inr_Foreach_kernelx652_inr_Foreach_concrete1( // @[:@63397.2]
  input         clock, // @[:@63398.4]
  input         reset, // @[:@63399.4]
  input  [31:0] io_in_b550_number, // @[:@63400.4]
  output [1:0]  io_in_x558_tmp_4_rPort_0_ofs_0, // @[:@63400.4]
  output        io_in_x558_tmp_4_rPort_0_en_0, // @[:@63400.4]
  input  [31:0] io_in_x558_tmp_4_rPort_0_output_0, // @[:@63400.4]
  output        io_in_x558_tmp_4_sEn_6, // @[:@63400.4]
  output        io_in_x558_tmp_4_sDone_6, // @[:@63400.4]
  output [1:0]  io_in_x545_accum_1_wPort_0_ofs_0, // @[:@63400.4]
  output [31:0] io_in_x545_accum_1_wPort_0_data_0, // @[:@63400.4]
  output        io_in_x545_accum_1_wPort_0_en_0, // @[:@63400.4]
  output [1:0]  io_in_x544_accum_0_rPort_0_ofs_0, // @[:@63400.4]
  output        io_in_x544_accum_0_rPort_0_en_0, // @[:@63400.4]
  input  [31:0] io_in_x544_accum_0_rPort_0_output_0, // @[:@63400.4]
  output [1:0]  io_in_x544_accum_0_wPort_0_ofs_0, // @[:@63400.4]
  output [31:0] io_in_x544_accum_0_wPort_0_data_0, // @[:@63400.4]
  output        io_in_x544_accum_0_wPort_0_en_0, // @[:@63400.4]
  input         io_in_b543, // @[:@63400.4]
  output [63:0] io_in_instrctrs_16_cycs, // @[:@63400.4]
  output [63:0] io_in_instrctrs_16_iters, // @[:@63400.4]
  input         io_sigsIn_done, // @[:@63400.4]
  input         io_sigsIn_datapathEn, // @[:@63400.4]
  input         io_sigsIn_baseEn, // @[:@63400.4]
  input         io_sigsIn_break, // @[:@63400.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@63400.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@63400.4]
  input         io_rr // @[:@63400.4]
);
  wire  cycles_x652_inr_Foreach_clock; // @[sm_x652_inr_Foreach.scala 77:43:@63590.4]
  wire  cycles_x652_inr_Foreach_reset; // @[sm_x652_inr_Foreach.scala 77:43:@63590.4]
  wire  cycles_x652_inr_Foreach_io_enable; // @[sm_x652_inr_Foreach.scala 77:43:@63590.4]
  wire [63:0] cycles_x652_inr_Foreach_io_count; // @[sm_x652_inr_Foreach.scala 77:43:@63590.4]
  wire  iters_x652_inr_Foreach_clock; // @[sm_x652_inr_Foreach.scala 78:42:@63593.4]
  wire  iters_x652_inr_Foreach_reset; // @[sm_x652_inr_Foreach.scala 78:42:@63593.4]
  wire  iters_x652_inr_Foreach_io_enable; // @[sm_x652_inr_Foreach.scala 78:42:@63593.4]
  wire [63:0] iters_x652_inr_Foreach_io_count; // @[sm_x652_inr_Foreach.scala 78:42:@63593.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@63610.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@63610.4]
  wire  x648_sum_1_clock; // @[Math.scala 150:24:@63669.4]
  wire  x648_sum_1_reset; // @[Math.scala 150:24:@63669.4]
  wire [31:0] x648_sum_1_io_a; // @[Math.scala 150:24:@63669.4]
  wire [31:0] x648_sum_1_io_b; // @[Math.scala 150:24:@63669.4]
  wire [31:0] x648_sum_1_io_result; // @[Math.scala 150:24:@63669.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@63680.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@63680.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@63680.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@63680.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@63680.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@63690.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@63690.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@63690.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@63690.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@63690.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@63703.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@63703.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@63703.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@63703.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@63703.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@63713.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@63713.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@63713.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@63713.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@63713.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@63723.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@63723.4]
  wire [31:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@63723.4]
  wire [31:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@63723.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@63737.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@63737.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@63737.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@63737.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@63737.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@63762.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@63762.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@63762.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@63762.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@63762.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@63782.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@63782.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@63782.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@63782.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@63782.4]
  wire  _T_750; // @[package.scala 100:49:@63597.4]
  reg  _T_753; // @[package.scala 48:56:@63598.4]
  reg [31:0] _RAND_0;
  wire  b553; // @[sm_x652_inr_Foreach.scala 83:18:@63618.4]
  wire  _T_778; // @[sm_x652_inr_Foreach.scala 88:114:@63624.4]
  wire  _T_779; // @[sm_x652_inr_Foreach.scala 88:111:@63625.4]
  wire  _T_784; // @[implicits.scala 56:10:@63628.4]
  wire  _T_785; // @[sm_x652_inr_Foreach.scala 88:131:@63629.4]
  wire  _T_786; // @[sm_x652_inr_Foreach.scala 88:228:@63630.4]
  wire [31:0] _T_820; // @[Math.scala 510:37:@63664.4]
  wire  x790_x647_D3; // @[package.scala 96:25:@63695.4 package.scala 96:25:@63696.4]
  wire [31:0] x789_x641_elem_0_D1_number; // @[package.scala 96:25:@63685.4 package.scala 96:25:@63686.4]
  wire [31:0] x648_sum_number; // @[Math.scala 154:22:@63675.4 Math.scala 155:14:@63676.4]
  wire  _T_864; // @[package.scala 96:25:@63742.4 package.scala 96:25:@63743.4]
  wire  _T_866; // @[implicits.scala 56:10:@63744.4]
  wire  _T_867; // @[sm_x652_inr_Foreach.scala 122:117:@63745.4]
  wire  _T_869; // @[sm_x652_inr_Foreach.scala 122:214:@63747.4]
  wire  x792_b553_D3; // @[package.scala 96:25:@63718.4 package.scala 96:25:@63719.4]
  wire  _T_871; // @[sm_x652_inr_Foreach.scala 122:259:@63749.4]
  wire  x791_b543_D3; // @[package.scala 96:25:@63708.4 package.scala 96:25:@63709.4]
  wire  _T_883; // @[package.scala 96:25:@63767.4 package.scala 96:25:@63768.4]
  wire  _T_885; // @[implicits.scala 56:10:@63769.4]
  wire  _T_886; // @[sm_x652_inr_Foreach.scala 127:117:@63770.4]
  wire  _T_888; // @[sm_x652_inr_Foreach.scala 127:214:@63772.4]
  wire  _T_890; // @[sm_x652_inr_Foreach.scala 127:259:@63774.4]
  wire  _T_895; // @[package.scala 96:25:@63787.4 package.scala 96:25:@63788.4]
  wire [31:0] b551_number; // @[Math.scala 723:22:@63615.4 Math.scala 724:14:@63616.4]
  wire [31:0] x793_b551_D3_number; // @[package.scala 96:25:@63728.4 package.scala 96:25:@63729.4]
  InstrumentationCounter cycles_x652_inr_Foreach ( // @[sm_x652_inr_Foreach.scala 77:43:@63590.4]
    .clock(cycles_x652_inr_Foreach_clock),
    .reset(cycles_x652_inr_Foreach_reset),
    .io_enable(cycles_x652_inr_Foreach_io_enable),
    .io_count(cycles_x652_inr_Foreach_io_count)
  );
  InstrumentationCounter iters_x652_inr_Foreach ( // @[sm_x652_inr_Foreach.scala 78:42:@63593.4]
    .clock(iters_x652_inr_Foreach_clock),
    .reset(iters_x652_inr_Foreach_reset),
    .io_enable(iters_x652_inr_Foreach_io_enable),
    .io_count(iters_x652_inr_Foreach_io_count)
  );
  _ _ ( // @[Math.scala 720:24:@63610.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x648_sum x648_sum_1 ( // @[Math.scala 150:24:@63669.4]
    .clock(x648_sum_1_clock),
    .reset(x648_sum_1_reset),
    .io_a(x648_sum_1_io_a),
    .io_b(x648_sum_1_io_b),
    .io_result(x648_sum_1_io_result)
  );
  RetimeWrapper_32 RetimeWrapper ( // @[package.scala 93:22:@63680.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_59 RetimeWrapper_1 ( // @[package.scala 93:22:@63690.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_59 RetimeWrapper_2 ( // @[package.scala 93:22:@63703.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_59 RetimeWrapper_3 ( // @[package.scala 93:22:@63713.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_718 RetimeWrapper_4 ( // @[package.scala 93:22:@63723.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_59 RetimeWrapper_5 ( // @[package.scala 93:22:@63737.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_59 RetimeWrapper_6 ( // @[package.scala 93:22:@63762.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@63782.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign _T_750 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@63597.4]
  assign b553 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x652_inr_Foreach.scala 83:18:@63618.4]
  assign _T_778 = ~ io_sigsIn_break; // @[sm_x652_inr_Foreach.scala 88:114:@63624.4]
  assign _T_779 = io_rr & _T_778; // @[sm_x652_inr_Foreach.scala 88:111:@63625.4]
  assign _T_784 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 56:10:@63628.4]
  assign _T_785 = _T_779 & _T_784; // @[sm_x652_inr_Foreach.scala 88:131:@63629.4]
  assign _T_786 = _T_785 & b553; // @[sm_x652_inr_Foreach.scala 88:228:@63630.4]
  assign _T_820 = $signed(io_in_b550_number); // @[Math.scala 510:37:@63664.4]
  assign x790_x647_D3 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@63695.4 package.scala 96:25:@63696.4]
  assign x789_x641_elem_0_D1_number = RetimeWrapper_io_out; // @[package.scala 96:25:@63685.4 package.scala 96:25:@63686.4]
  assign x648_sum_number = x648_sum_1_io_result; // @[Math.scala 154:22:@63675.4 Math.scala 155:14:@63676.4]
  assign _T_864 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@63742.4 package.scala 96:25:@63743.4]
  assign _T_866 = io_rr ? _T_864 : 1'h0; // @[implicits.scala 56:10:@63744.4]
  assign _T_867 = _T_778 & _T_866; // @[sm_x652_inr_Foreach.scala 122:117:@63745.4]
  assign _T_869 = _T_867 & _T_778; // @[sm_x652_inr_Foreach.scala 122:214:@63747.4]
  assign x792_b553_D3 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@63718.4 package.scala 96:25:@63719.4]
  assign _T_871 = _T_869 & x792_b553_D3; // @[sm_x652_inr_Foreach.scala 122:259:@63749.4]
  assign x791_b543_D3 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@63708.4 package.scala 96:25:@63709.4]
  assign _T_883 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@63767.4 package.scala 96:25:@63768.4]
  assign _T_885 = io_rr ? _T_883 : 1'h0; // @[implicits.scala 56:10:@63769.4]
  assign _T_886 = _T_778 & _T_885; // @[sm_x652_inr_Foreach.scala 127:117:@63770.4]
  assign _T_888 = _T_886 & _T_778; // @[sm_x652_inr_Foreach.scala 127:214:@63772.4]
  assign _T_890 = _T_888 & x792_b553_D3; // @[sm_x652_inr_Foreach.scala 127:259:@63774.4]
  assign _T_895 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@63787.4 package.scala 96:25:@63788.4]
  assign b551_number = __io_result; // @[Math.scala 723:22:@63615.4 Math.scala 724:14:@63616.4]
  assign x793_b551_D3_number = RetimeWrapper_4_io_out; // @[package.scala 96:25:@63728.4 package.scala 96:25:@63729.4]
  assign io_in_x558_tmp_4_rPort_0_ofs_0 = b551_number[1:0]; // @[MemInterfaceType.scala 107:54:@63634.4]
  assign io_in_x558_tmp_4_rPort_0_en_0 = _T_786 & io_in_b543; // @[MemInterfaceType.scala 110:79:@63636.4]
  assign io_in_x558_tmp_4_sEn_6 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@63790.4]
  assign io_in_x558_tmp_4_sDone_6 = io_rr ? _T_895 : 1'h0; // @[MemInterfaceType.scala 197:17:@63791.4]
  assign io_in_x545_accum_1_wPort_0_ofs_0 = x793_b551_D3_number[1:0]; // @[MemInterfaceType.scala 89:54:@63752.4]
  assign io_in_x545_accum_1_wPort_0_data_0 = x790_x647_D3 ? x789_x641_elem_0_D1_number : x648_sum_number; // @[MemInterfaceType.scala 90:56:@63753.4]
  assign io_in_x545_accum_1_wPort_0_en_0 = _T_871 & x791_b543_D3; // @[MemInterfaceType.scala 93:57:@63755.4]
  assign io_in_x544_accum_0_rPort_0_ofs_0 = b551_number[1:0]; // @[MemInterfaceType.scala 107:54:@63655.4]
  assign io_in_x544_accum_0_rPort_0_en_0 = _T_786 & io_in_b543; // @[MemInterfaceType.scala 110:79:@63657.4]
  assign io_in_x544_accum_0_wPort_0_ofs_0 = x793_b551_D3_number[1:0]; // @[MemInterfaceType.scala 89:54:@63777.4]
  assign io_in_x544_accum_0_wPort_0_data_0 = x790_x647_D3 ? x789_x641_elem_0_D1_number : x648_sum_number; // @[MemInterfaceType.scala 90:56:@63778.4]
  assign io_in_x544_accum_0_wPort_0_en_0 = _T_890 & x791_b543_D3; // @[MemInterfaceType.scala 93:57:@63780.4]
  assign io_in_instrctrs_16_cycs = cycles_x652_inr_Foreach_io_count; // @[Ledger.scala 293:21:@63602.4]
  assign io_in_instrctrs_16_iters = iters_x652_inr_Foreach_io_count; // @[Ledger.scala 294:22:@63603.4]
  assign cycles_x652_inr_Foreach_clock = clock; // @[:@63591.4]
  assign cycles_x652_inr_Foreach_reset = reset; // @[:@63592.4]
  assign cycles_x652_inr_Foreach_io_enable = io_sigsIn_baseEn; // @[sm_x652_inr_Foreach.scala 79:41:@63596.4]
  assign iters_x652_inr_Foreach_clock = clock; // @[:@63594.4]
  assign iters_x652_inr_Foreach_reset = reset; // @[:@63595.4]
  assign iters_x652_inr_Foreach_io_enable = io_sigsIn_done & _T_753; // @[sm_x652_inr_Foreach.scala 80:40:@63601.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@63613.4]
  assign x648_sum_1_clock = clock; // @[:@63670.4]
  assign x648_sum_1_reset = reset; // @[:@63671.4]
  assign x648_sum_1_io_a = io_in_x558_tmp_4_rPort_0_output_0; // @[Math.scala 151:17:@63672.4]
  assign x648_sum_1_io_b = io_in_x544_accum_0_rPort_0_output_0; // @[Math.scala 152:17:@63673.4]
  assign RetimeWrapper_clock = clock; // @[:@63681.4]
  assign RetimeWrapper_reset = reset; // @[:@63682.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@63684.4]
  assign RetimeWrapper_io_in = io_in_x558_tmp_4_rPort_0_output_0; // @[package.scala 94:16:@63683.4]
  assign RetimeWrapper_1_clock = clock; // @[:@63691.4]
  assign RetimeWrapper_1_reset = reset; // @[:@63692.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@63694.4]
  assign RetimeWrapper_1_io_in = $signed(_T_820) == $signed(32'sh0); // @[package.scala 94:16:@63693.4]
  assign RetimeWrapper_2_clock = clock; // @[:@63704.4]
  assign RetimeWrapper_2_reset = reset; // @[:@63705.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@63707.4]
  assign RetimeWrapper_2_io_in = io_in_b543; // @[package.scala 94:16:@63706.4]
  assign RetimeWrapper_3_clock = clock; // @[:@63714.4]
  assign RetimeWrapper_3_reset = reset; // @[:@63715.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@63717.4]
  assign RetimeWrapper_3_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@63716.4]
  assign RetimeWrapper_4_clock = clock; // @[:@63724.4]
  assign RetimeWrapper_4_reset = reset; // @[:@63725.4]
  assign RetimeWrapper_4_io_in = __io_result; // @[package.scala 94:16:@63726.4]
  assign RetimeWrapper_5_clock = clock; // @[:@63738.4]
  assign RetimeWrapper_5_reset = reset; // @[:@63739.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@63741.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@63740.4]
  assign RetimeWrapper_6_clock = clock; // @[:@63763.4]
  assign RetimeWrapper_6_reset = reset; // @[:@63764.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@63766.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@63765.4]
  assign RetimeWrapper_7_clock = clock; // @[:@63783.4]
  assign RetimeWrapper_7_reset = reset; // @[:@63784.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@63786.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_done; // @[package.scala 94:16:@63785.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_753 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_753 <= 1'h0;
    end else begin
      _T_753 <= _T_750;
    end
  end
endmodule
module x653_outr_Reduce_kernelx653_outr_Reduce_concrete1( // @[:@63825.2]
  input         clock, // @[:@63826.4]
  input         reset, // @[:@63827.4]
  output [8:0]  io_in_x472_A_sram_1_rPort_0_ofs_0, // @[:@63828.4]
  output        io_in_x472_A_sram_1_rPort_0_en_0, // @[:@63828.4]
  input  [31:0] io_in_x472_A_sram_1_rPort_0_output_0, // @[:@63828.4]
  input  [31:0] io_in_b542_number, // @[:@63828.4]
  output [8:0]  io_in_x471_A_sram_0_rPort_0_ofs_0, // @[:@63828.4]
  output        io_in_x471_A_sram_0_rPort_0_en_0, // @[:@63828.4]
  input  [31:0] io_in_x471_A_sram_0_rPort_0_output_0, // @[:@63828.4]
  output [1:0]  io_in_x545_accum_1_wPort_0_ofs_0, // @[:@63828.4]
  output [31:0] io_in_x545_accum_1_wPort_0_data_0, // @[:@63828.4]
  output        io_in_x545_accum_1_wPort_0_en_0, // @[:@63828.4]
  output        io_in_x545_accum_1_sEn_0, // @[:@63828.4]
  output        io_in_x545_accum_1_sDone_0, // @[:@63828.4]
  output [1:0]  io_in_x544_accum_0_rPort_0_ofs_0, // @[:@63828.4]
  output        io_in_x544_accum_0_rPort_0_en_0, // @[:@63828.4]
  input  [31:0] io_in_x544_accum_0_rPort_0_output_0, // @[:@63828.4]
  output [1:0]  io_in_x544_accum_0_wPort_0_ofs_0, // @[:@63828.4]
  output [31:0] io_in_x544_accum_0_wPort_0_data_0, // @[:@63828.4]
  output        io_in_x544_accum_0_wPort_0_en_0, // @[:@63828.4]
  output        io_in_x549_ctrchain_input_reset, // @[:@63828.4]
  output        io_in_x549_ctrchain_input_enable, // @[:@63828.4]
  input  [3:0]  io_in_x549_ctrchain_output_counts_0, // @[:@63828.4]
  input         io_in_x549_ctrchain_output_oobs_0, // @[:@63828.4]
  input         io_in_x549_ctrchain_output_done, // @[:@63828.4]
  input         io_in_b543, // @[:@63828.4]
  output [63:0] io_in_instrctrs_7_cycs, // @[:@63828.4]
  output [63:0] io_in_instrctrs_7_iters, // @[:@63828.4]
  output [63:0] io_in_instrctrs_8_cycs, // @[:@63828.4]
  output [63:0] io_in_instrctrs_8_iters, // @[:@63828.4]
  output [63:0] io_in_instrctrs_9_cycs, // @[:@63828.4]
  output [63:0] io_in_instrctrs_9_iters, // @[:@63828.4]
  output [63:0] io_in_instrctrs_10_cycs, // @[:@63828.4]
  output [63:0] io_in_instrctrs_10_iters, // @[:@63828.4]
  output [63:0] io_in_instrctrs_11_cycs, // @[:@63828.4]
  output [63:0] io_in_instrctrs_11_iters, // @[:@63828.4]
  output [63:0] io_in_instrctrs_12_cycs, // @[:@63828.4]
  output [63:0] io_in_instrctrs_12_iters, // @[:@63828.4]
  output [63:0] io_in_instrctrs_13_cycs, // @[:@63828.4]
  output [63:0] io_in_instrctrs_13_iters, // @[:@63828.4]
  output [63:0] io_in_instrctrs_14_cycs, // @[:@63828.4]
  output [63:0] io_in_instrctrs_14_iters, // @[:@63828.4]
  output [63:0] io_in_instrctrs_15_cycs, // @[:@63828.4]
  output [63:0] io_in_instrctrs_15_iters, // @[:@63828.4]
  output [63:0] io_in_instrctrs_16_cycs, // @[:@63828.4]
  output [63:0] io_in_instrctrs_16_iters, // @[:@63828.4]
  input         io_sigsIn_done, // @[:@63828.4]
  input         io_sigsIn_baseEn, // @[:@63828.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@63828.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@63828.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@63828.4]
  input         io_sigsIn_smEnableOuts_3, // @[:@63828.4]
  input         io_sigsIn_smEnableOuts_4, // @[:@63828.4]
  input         io_sigsIn_smEnableOuts_5, // @[:@63828.4]
  input         io_sigsIn_smEnableOuts_6, // @[:@63828.4]
  input         io_sigsIn_smChildAcks_0, // @[:@63828.4]
  input         io_sigsIn_smChildAcks_1, // @[:@63828.4]
  input         io_sigsIn_smChildAcks_2, // @[:@63828.4]
  input         io_sigsIn_smChildAcks_3, // @[:@63828.4]
  input         io_sigsIn_smChildAcks_4, // @[:@63828.4]
  input         io_sigsIn_smChildAcks_5, // @[:@63828.4]
  input         io_sigsIn_smChildAcks_6, // @[:@63828.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@63828.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@63828.4]
  output        io_sigsOut_smDoneIn_0, // @[:@63828.4]
  output        io_sigsOut_smDoneIn_1, // @[:@63828.4]
  output        io_sigsOut_smDoneIn_2, // @[:@63828.4]
  output        io_sigsOut_smDoneIn_3, // @[:@63828.4]
  output        io_sigsOut_smDoneIn_4, // @[:@63828.4]
  output        io_sigsOut_smDoneIn_5, // @[:@63828.4]
  output        io_sigsOut_smDoneIn_6, // @[:@63828.4]
  output        io_sigsOut_smMaskIn_0, // @[:@63828.4]
  output        io_sigsOut_smMaskIn_1, // @[:@63828.4]
  output        io_sigsOut_smMaskIn_2, // @[:@63828.4]
  output        io_sigsOut_smMaskIn_4, // @[:@63828.4]
  output        io_sigsOut_smMaskIn_5, // @[:@63828.4]
  input         io_rr // @[:@63828.4]
);
  wire  cycles_x653_outr_Reduce_clock; // @[sm_x653_outr_Reduce.scala 86:43:@64023.4]
  wire  cycles_x653_outr_Reduce_reset; // @[sm_x653_outr_Reduce.scala 86:43:@64023.4]
  wire  cycles_x653_outr_Reduce_io_enable; // @[sm_x653_outr_Reduce.scala 86:43:@64023.4]
  wire [63:0] cycles_x653_outr_Reduce_io_count; // @[sm_x653_outr_Reduce.scala 86:43:@64023.4]
  wire  iters_x653_outr_Reduce_clock; // @[sm_x653_outr_Reduce.scala 87:42:@64026.4]
  wire  iters_x653_outr_Reduce_reset; // @[sm_x653_outr_Reduce.scala 87:42:@64026.4]
  wire  iters_x653_outr_Reduce_io_enable; // @[sm_x653_outr_Reduce.scala 87:42:@64026.4]
  wire [63:0] iters_x653_outr_Reduce_io_count; // @[sm_x653_outr_Reduce.scala 87:42:@64026.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@64043.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@64043.4]
  wire  b550_chain_clock; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_reset; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire [31:0] b550_chain_io_rPort_5_output_0; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire [31:0] b550_chain_io_rPort_4_output_0; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire [31:0] b550_chain_io_rPort_3_output_0; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire [31:0] b550_chain_io_rPort_2_output_0; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire [31:0] b550_chain_io_rPort_1_output_0; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire [31:0] b550_chain_io_rPort_0_output_0; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire [31:0] b550_chain_io_wPort_0_data_0; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_io_wPort_0_reset; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_io_wPort_0_en_0; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_io_sEn_0; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_io_sEn_1; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_io_sEn_2; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_io_sEn_3; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_io_sEn_4; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_io_sEn_5; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_io_sEn_6; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_io_sDone_0; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_io_sDone_1; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_io_sDone_2; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_io_sDone_3; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_io_sDone_4; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_io_sDone_5; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  b550_chain_io_sDone_6; // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@64115.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@64115.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@64115.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@64115.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@64115.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@64127.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@64127.4]
  wire [31:0] __2_io_b; // @[Math.scala 720:24:@64138.4]
  wire [31:0] __2_io_result; // @[Math.scala 720:24:@64138.4]
  wire [31:0] __3_io_b; // @[Math.scala 720:24:@64149.4]
  wire [31:0] __3_io_result; // @[Math.scala 720:24:@64149.4]
  wire [31:0] __4_io_b; // @[Math.scala 720:24:@64160.4]
  wire [31:0] __4_io_result; // @[Math.scala 720:24:@64160.4]
  wire [31:0] __5_io_b; // @[Math.scala 720:24:@64171.4]
  wire [31:0] __5_io_result; // @[Math.scala 720:24:@64171.4]
  wire [31:0] __6_io_b; // @[Math.scala 720:24:@64182.4]
  wire [31:0] __6_io_result; // @[Math.scala 720:24:@64182.4]
  wire  b552_chain_clock; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_reset; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_rPort_4_output_0; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_rPort_3_output_0; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_rPort_1_output_0; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_rPort_0_output_0; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_wPort_0_data_0; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_wPort_0_reset; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_wPort_0_en_0; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_sEn_0; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_sEn_1; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_sEn_2; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_sEn_3; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_sEn_4; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_sEn_5; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_sEn_6; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_sDone_0; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_sDone_1; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_sDone_2; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_sDone_3; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_sDone_4; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_sDone_5; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  b552_chain_io_sDone_6; // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@64255.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@64255.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@64255.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@64255.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@64255.4]
  wire  x554_tmp_0_clock; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x554_tmp_0_reset; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire [1:0] x554_tmp_0_io_rPort_0_ofs_0; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x554_tmp_0_io_rPort_0_en_0; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire [31:0] x554_tmp_0_io_rPort_0_output_0; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire [1:0] x554_tmp_0_io_wPort_1_ofs_0; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire [31:0] x554_tmp_0_io_wPort_1_data_0; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x554_tmp_0_io_wPort_1_en_0; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire [1:0] x554_tmp_0_io_wPort_0_ofs_0; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire [31:0] x554_tmp_0_io_wPort_0_data_0; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x554_tmp_0_io_wPort_0_en_0; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x554_tmp_0_io_sEn_0; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x554_tmp_0_io_sEn_1; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x554_tmp_0_io_sEn_2; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x554_tmp_0_io_sEn_3; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x554_tmp_0_io_sEn_4; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x554_tmp_0_io_sEn_5; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x554_tmp_0_io_sDone_0; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x554_tmp_0_io_sDone_1; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x554_tmp_0_io_sDone_2; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x554_tmp_0_io_sDone_3; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x554_tmp_0_io_sDone_4; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x554_tmp_0_io_sDone_5; // @[m_x554_tmp_0.scala 28:22:@64270.4]
  wire  x555_tmp_1_clock; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x555_tmp_1_reset; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire [1:0] x555_tmp_1_io_rPort_0_ofs_0; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x555_tmp_1_io_rPort_0_en_0; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire [31:0] x555_tmp_1_io_rPort_0_output_0; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire [1:0] x555_tmp_1_io_wPort_1_ofs_0; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire [31:0] x555_tmp_1_io_wPort_1_data_0; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x555_tmp_1_io_wPort_1_en_0; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire [1:0] x555_tmp_1_io_wPort_0_ofs_0; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire [31:0] x555_tmp_1_io_wPort_0_data_0; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x555_tmp_1_io_wPort_0_en_0; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x555_tmp_1_io_sEn_0; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x555_tmp_1_io_sEn_1; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x555_tmp_1_io_sEn_2; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x555_tmp_1_io_sEn_3; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x555_tmp_1_io_sEn_4; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x555_tmp_1_io_sEn_5; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x555_tmp_1_io_sDone_0; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x555_tmp_1_io_sDone_1; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x555_tmp_1_io_sDone_2; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x555_tmp_1_io_sDone_3; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x555_tmp_1_io_sDone_4; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x555_tmp_1_io_sDone_5; // @[m_x555_tmp_1.scala 28:22:@64317.4]
  wire  x556_tmp_2_clock; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x556_tmp_2_reset; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire [1:0] x556_tmp_2_io_rPort_0_ofs_0; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x556_tmp_2_io_rPort_0_en_0; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire [31:0] x556_tmp_2_io_rPort_0_output_0; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire [1:0] x556_tmp_2_io_wPort_1_ofs_0; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire [31:0] x556_tmp_2_io_wPort_1_data_0; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x556_tmp_2_io_wPort_1_en_0; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire [1:0] x556_tmp_2_io_wPort_0_ofs_0; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire [31:0] x556_tmp_2_io_wPort_0_data_0; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x556_tmp_2_io_wPort_0_en_0; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x556_tmp_2_io_sEn_0; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x556_tmp_2_io_sEn_1; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x556_tmp_2_io_sEn_2; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x556_tmp_2_io_sEn_3; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x556_tmp_2_io_sEn_4; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x556_tmp_2_io_sEn_5; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x556_tmp_2_io_sDone_0; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x556_tmp_2_io_sDone_1; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x556_tmp_2_io_sDone_2; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x556_tmp_2_io_sDone_3; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x556_tmp_2_io_sDone_4; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x556_tmp_2_io_sDone_5; // @[m_x556_tmp_2.scala 28:22:@64364.4]
  wire  x557_tmp_3_clock; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x557_tmp_3_reset; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire [1:0] x557_tmp_3_io_rPort_0_ofs_0; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x557_tmp_3_io_rPort_0_en_0; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire [31:0] x557_tmp_3_io_rPort_0_output_0; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire [1:0] x557_tmp_3_io_wPort_1_ofs_0; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire [31:0] x557_tmp_3_io_wPort_1_data_0; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x557_tmp_3_io_wPort_1_en_0; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire [1:0] x557_tmp_3_io_wPort_0_ofs_0; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire [31:0] x557_tmp_3_io_wPort_0_data_0; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x557_tmp_3_io_wPort_0_en_0; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x557_tmp_3_io_sEn_0; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x557_tmp_3_io_sEn_1; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x557_tmp_3_io_sEn_2; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x557_tmp_3_io_sEn_3; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x557_tmp_3_io_sEn_4; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x557_tmp_3_io_sEn_5; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x557_tmp_3_io_sDone_0; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x557_tmp_3_io_sDone_1; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x557_tmp_3_io_sDone_2; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x557_tmp_3_io_sDone_3; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x557_tmp_3_io_sDone_4; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x557_tmp_3_io_sDone_5; // @[m_x557_tmp_3.scala 28:22:@64411.4]
  wire  x558_tmp_4_clock; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_reset; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire [1:0] x558_tmp_4_io_rPort_0_ofs_0; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_rPort_0_en_0; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire [31:0] x558_tmp_4_io_rPort_0_output_0; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire [1:0] x558_tmp_4_io_wPort_1_ofs_0; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire [31:0] x558_tmp_4_io_wPort_1_data_0; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_wPort_1_en_0; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire [1:0] x558_tmp_4_io_wPort_0_ofs_0; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire [31:0] x558_tmp_4_io_wPort_0_data_0; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_wPort_0_en_0; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_sEn_0; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_sEn_1; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_sEn_2; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_sEn_3; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_sEn_4; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_sEn_5; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_sEn_6; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_sDone_0; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_sDone_1; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_sDone_2; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_sDone_3; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_sDone_4; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_sDone_5; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x558_tmp_4_io_sDone_6; // @[m_x558_tmp_4.scala 28:22:@64458.4]
  wire  x560_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@64507.4]
  wire  x560_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@64507.4]
  wire  x560_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@64507.4]
  wire  x560_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@64507.4]
  wire [3:0] x560_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@64507.4]
  wire  x560_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@64507.4]
  wire  x560_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@64507.4]
  wire  x579_inr_Foreach_sm_clock; // @[sm_x579_inr_Foreach.scala 35:18:@64560.4]
  wire  x579_inr_Foreach_sm_reset; // @[sm_x579_inr_Foreach.scala 35:18:@64560.4]
  wire  x579_inr_Foreach_sm_io_enable; // @[sm_x579_inr_Foreach.scala 35:18:@64560.4]
  wire  x579_inr_Foreach_sm_io_done; // @[sm_x579_inr_Foreach.scala 35:18:@64560.4]
  wire  x579_inr_Foreach_sm_io_ctrDone; // @[sm_x579_inr_Foreach.scala 35:18:@64560.4]
  wire  x579_inr_Foreach_sm_io_datapathEn; // @[sm_x579_inr_Foreach.scala 35:18:@64560.4]
  wire  x579_inr_Foreach_sm_io_ctrInc; // @[sm_x579_inr_Foreach.scala 35:18:@64560.4]
  wire  x579_inr_Foreach_sm_io_ctrRst; // @[sm_x579_inr_Foreach.scala 35:18:@64560.4]
  wire  x579_inr_Foreach_sm_io_parentAck; // @[sm_x579_inr_Foreach.scala 35:18:@64560.4]
  wire  x579_inr_Foreach_sm_io_backpressure; // @[sm_x579_inr_Foreach.scala 35:18:@64560.4]
  wire  x579_inr_Foreach_sm_io_break; // @[sm_x579_inr_Foreach.scala 35:18:@64560.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@64589.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@64589.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@64589.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@64589.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@64589.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@64598.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@64598.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@64598.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@64598.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@64598.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@64608.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@64608.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@64608.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@64608.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@64608.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@64650.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@64650.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@64650.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@64650.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@64650.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@64658.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@64658.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@64658.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@64658.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@64658.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_clock; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_reset; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [1:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_ofs_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_data_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_en_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_sEn_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_sDone_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b550_number; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [8:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_en_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_output_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b542_number; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [8:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_en_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_output_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [1:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_ofs_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_data_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_en_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_sEn_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_sDone_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [1:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_ofs_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_data_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_en_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b552; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [1:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_ofs_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_data_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_en_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_sEn_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_sDone_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [1:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_ofs_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_data_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_en_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_sEn_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_sDone_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b543; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [63:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_instrctrs_8_cycs; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [63:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_instrctrs_8_iters; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_done; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_rr; // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
  wire  x580_r_0_clock; // @[m_x580_r_0.scala 28:22:@65236.4]
  wire  x580_r_0_reset; // @[m_x580_r_0.scala 28:22:@65236.4]
  wire  x580_r_0_io_rPort_1_en_0; // @[m_x580_r_0.scala 28:22:@65236.4]
  wire [31:0] x580_r_0_io_rPort_1_output_0; // @[m_x580_r_0.scala 28:22:@65236.4]
  wire  x580_r_0_io_rPort_0_en_0; // @[m_x580_r_0.scala 28:22:@65236.4]
  wire [31:0] x580_r_0_io_rPort_0_output_0; // @[m_x580_r_0.scala 28:22:@65236.4]
  wire [31:0] x580_r_0_io_wPort_0_data_0; // @[m_x580_r_0.scala 28:22:@65236.4]
  wire  x580_r_0_io_wPort_0_en_0; // @[m_x580_r_0.scala 28:22:@65236.4]
  wire  x580_r_0_io_sEn_0; // @[m_x580_r_0.scala 28:22:@65236.4]
  wire  x580_r_0_io_sEn_1; // @[m_x580_r_0.scala 28:22:@65236.4]
  wire  x580_r_0_io_sEn_2; // @[m_x580_r_0.scala 28:22:@65236.4]
  wire  x580_r_0_io_sDone_0; // @[m_x580_r_0.scala 28:22:@65236.4]
  wire  x580_r_0_io_sDone_1; // @[m_x580_r_0.scala 28:22:@65236.4]
  wire  x580_r_0_io_sDone_2; // @[m_x580_r_0.scala 28:22:@65236.4]
  wire  x593_inr_UnitPipe_sm_clock; // @[sm_x593_inr_UnitPipe.scala 33:18:@65311.4]
  wire  x593_inr_UnitPipe_sm_reset; // @[sm_x593_inr_UnitPipe.scala 33:18:@65311.4]
  wire  x593_inr_UnitPipe_sm_io_enable; // @[sm_x593_inr_UnitPipe.scala 33:18:@65311.4]
  wire  x593_inr_UnitPipe_sm_io_done; // @[sm_x593_inr_UnitPipe.scala 33:18:@65311.4]
  wire  x593_inr_UnitPipe_sm_io_ctrDone; // @[sm_x593_inr_UnitPipe.scala 33:18:@65311.4]
  wire  x593_inr_UnitPipe_sm_io_datapathEn; // @[sm_x593_inr_UnitPipe.scala 33:18:@65311.4]
  wire  x593_inr_UnitPipe_sm_io_ctrInc; // @[sm_x593_inr_UnitPipe.scala 33:18:@65311.4]
  wire  x593_inr_UnitPipe_sm_io_parentAck; // @[sm_x593_inr_UnitPipe.scala 33:18:@65311.4]
  wire  x593_inr_UnitPipe_sm_io_backpressure; // @[sm_x593_inr_UnitPipe.scala 33:18:@65311.4]
  wire  x593_inr_UnitPipe_sm_io_break; // @[sm_x593_inr_UnitPipe.scala 33:18:@65311.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@65344.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@65344.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@65344.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@65344.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@65344.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@65354.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@65354.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@65354.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@65354.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@65354.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@65390.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@65390.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@65390.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@65390.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@65390.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@65398.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@65398.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@65398.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@65398.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@65398.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_clock; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_reset; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_rPort_0_en_0; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire [31:0] x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_rPort_0_output_0; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_1; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_1; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_rPort_0_en_0; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire [31:0] x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_rPort_0_output_0; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_1; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_1; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_1; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_1; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_1; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_1; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire [31:0] x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_wPort_0_data_0; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_wPort_0_en_0; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_sEn_0; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_sDone_0; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_rPort_0_en_0; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire [31:0] x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_rPort_0_output_0; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_1; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_1; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire [63:0] x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_instrctrs_9_cycs; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire [63:0] x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_instrctrs_9_iters; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_done; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_baseEn; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_break; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_rr; // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
  wire  x594_force_0_clock; // @[m_x594_force_0.scala 27:22:@65971.4]
  wire  x594_force_0_reset; // @[m_x594_force_0.scala 27:22:@65971.4]
  wire  x594_force_0_io_rPort_0_en_0; // @[m_x594_force_0.scala 27:22:@65971.4]
  wire [31:0] x594_force_0_io_rPort_0_output_0; // @[m_x594_force_0.scala 27:22:@65971.4]
  wire [31:0] x594_force_0_io_wPort_0_data_0; // @[m_x594_force_0.scala 27:22:@65971.4]
  wire  x594_force_0_io_wPort_0_en_0; // @[m_x594_force_0.scala 27:22:@65971.4]
  wire  x594_force_0_io_sEn_0; // @[m_x594_force_0.scala 27:22:@65971.4]
  wire  x594_force_0_io_sEn_1; // @[m_x594_force_0.scala 27:22:@65971.4]
  wire  x594_force_0_io_sDone_0; // @[m_x594_force_0.scala 27:22:@65971.4]
  wire  x594_force_0_io_sDone_1; // @[m_x594_force_0.scala 27:22:@65971.4]
  wire  x595_reg_clock; // @[m_x595_reg.scala 28:22:@66001.4]
  wire  x595_reg_reset; // @[m_x595_reg.scala 28:22:@66001.4]
  wire  x595_reg_io_rPort_1_output_0; // @[m_x595_reg.scala 28:22:@66001.4]
  wire  x595_reg_io_rPort_0_output_0; // @[m_x595_reg.scala 28:22:@66001.4]
  wire  x595_reg_io_wPort_0_data_0; // @[m_x595_reg.scala 28:22:@66001.4]
  wire  x595_reg_io_wPort_0_reset; // @[m_x595_reg.scala 28:22:@66001.4]
  wire  x595_reg_io_wPort_0_en_0; // @[m_x595_reg.scala 28:22:@66001.4]
  wire  x595_reg_io_sEn_0; // @[m_x595_reg.scala 28:22:@66001.4]
  wire  x595_reg_io_sEn_1; // @[m_x595_reg.scala 28:22:@66001.4]
  wire  x595_reg_io_sDone_0; // @[m_x595_reg.scala 28:22:@66001.4]
  wire  x595_reg_io_sDone_1; // @[m_x595_reg.scala 28:22:@66001.4]
  wire  x596_reg_clock; // @[m_x596_reg.scala 27:22:@66038.4]
  wire  x596_reg_reset; // @[m_x596_reg.scala 27:22:@66038.4]
  wire  x596_reg_io_rPort_0_output_0; // @[m_x596_reg.scala 27:22:@66038.4]
  wire  x596_reg_io_wPort_0_data_0; // @[m_x596_reg.scala 27:22:@66038.4]
  wire  x596_reg_io_wPort_0_reset; // @[m_x596_reg.scala 27:22:@66038.4]
  wire  x596_reg_io_wPort_0_en_0; // @[m_x596_reg.scala 27:22:@66038.4]
  wire  x596_reg_io_sEn_0; // @[m_x596_reg.scala 27:22:@66038.4]
  wire  x596_reg_io_sEn_1; // @[m_x596_reg.scala 27:22:@66038.4]
  wire  x596_reg_io_sDone_0; // @[m_x596_reg.scala 27:22:@66038.4]
  wire  x596_reg_io_sDone_1; // @[m_x596_reg.scala 27:22:@66038.4]
  wire  x605_inr_UnitPipe_sm_clock; // @[sm_x605_inr_UnitPipe.scala 33:18:@66104.4]
  wire  x605_inr_UnitPipe_sm_reset; // @[sm_x605_inr_UnitPipe.scala 33:18:@66104.4]
  wire  x605_inr_UnitPipe_sm_io_enable; // @[sm_x605_inr_UnitPipe.scala 33:18:@66104.4]
  wire  x605_inr_UnitPipe_sm_io_done; // @[sm_x605_inr_UnitPipe.scala 33:18:@66104.4]
  wire  x605_inr_UnitPipe_sm_io_doneLatch; // @[sm_x605_inr_UnitPipe.scala 33:18:@66104.4]
  wire  x605_inr_UnitPipe_sm_io_ctrDone; // @[sm_x605_inr_UnitPipe.scala 33:18:@66104.4]
  wire  x605_inr_UnitPipe_sm_io_datapathEn; // @[sm_x605_inr_UnitPipe.scala 33:18:@66104.4]
  wire  x605_inr_UnitPipe_sm_io_ctrInc; // @[sm_x605_inr_UnitPipe.scala 33:18:@66104.4]
  wire  x605_inr_UnitPipe_sm_io_ctrRst; // @[sm_x605_inr_UnitPipe.scala 33:18:@66104.4]
  wire  x605_inr_UnitPipe_sm_io_parentAck; // @[sm_x605_inr_UnitPipe.scala 33:18:@66104.4]
  wire  x605_inr_UnitPipe_sm_io_backpressure; // @[sm_x605_inr_UnitPipe.scala 33:18:@66104.4]
  wire  x605_inr_UnitPipe_sm_io_break; // @[sm_x605_inr_UnitPipe.scala 33:18:@66104.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@66137.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@66137.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@66137.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@66137.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@66137.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@66147.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@66147.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@66147.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@66147.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@66147.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@66183.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@66183.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@66183.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@66183.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@66183.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@66191.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@66191.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@66191.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@66191.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@66191.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_clock; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_reset; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_2; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_2; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_2; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_2; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_2; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_2; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_2; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_2; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_rPort_0_en_0; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire [31:0] x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_rPort_0_output_0; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_sEn_1; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_sDone_1; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_data_0; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_reset; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_en_0; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_reset; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_sEn_0; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_sDone_0; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_2; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_2; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_data_0; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_reset; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_en_0; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_reset; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_sEn_0; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_sDone_0; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire [63:0] x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_instrctrs_10_cycs; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire [63:0] x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_instrctrs_10_iters; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_done; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_baseEn; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_break; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_rr; // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
  wire  x621_inr_Switch_sm_clock; // @[sm_x621_inr_Switch.scala 33:18:@66923.4]
  wire  x621_inr_Switch_sm_reset; // @[sm_x621_inr_Switch.scala 33:18:@66923.4]
  wire  x621_inr_Switch_sm_io_enable; // @[sm_x621_inr_Switch.scala 33:18:@66923.4]
  wire  x621_inr_Switch_sm_io_done; // @[sm_x621_inr_Switch.scala 33:18:@66923.4]
  wire  x621_inr_Switch_sm_io_parentAck; // @[sm_x621_inr_Switch.scala 33:18:@66923.4]
  wire  x621_inr_Switch_sm_io_backpressure; // @[sm_x621_inr_Switch.scala 33:18:@66923.4]
  wire  x621_inr_Switch_sm_io_doneIn_0; // @[sm_x621_inr_Switch.scala 33:18:@66923.4]
  wire  x621_inr_Switch_sm_io_doneIn_1; // @[sm_x621_inr_Switch.scala 33:18:@66923.4]
  wire  x621_inr_Switch_sm_io_childAck_0; // @[sm_x621_inr_Switch.scala 33:18:@66923.4]
  wire  x621_inr_Switch_sm_io_childAck_1; // @[sm_x621_inr_Switch.scala 33:18:@66923.4]
  wire  x621_inr_Switch_sm_io_selectsIn_0; // @[sm_x621_inr_Switch.scala 33:18:@66923.4]
  wire  x621_inr_Switch_sm_io_selectsIn_1; // @[sm_x621_inr_Switch.scala 33:18:@66923.4]
  wire  x621_inr_Switch_sm_io_selectsOut_0; // @[sm_x621_inr_Switch.scala 33:18:@66923.4]
  wire  x621_inr_Switch_sm_io_selectsOut_1; // @[sm_x621_inr_Switch.scala 33:18:@66923.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@66960.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@66960.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@66960.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@66960.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@66960.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@66970.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@66970.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@66970.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@66970.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@66970.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@67012.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@67012.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@67012.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@67012.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@67012.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@67020.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@67020.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@67020.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@67020.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@67020.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_clock; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_reset; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x555_tmp_1_sEn_3; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x555_tmp_1_sDone_3; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x554_tmp_0_sEn_3; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x554_tmp_0_sDone_3; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x558_tmp_4_sEn_3; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x558_tmp_4_sDone_3; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x736_rd_x596; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x557_tmp_3_sEn_3; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x557_tmp_3_sDone_3; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_rPort_1_en_0; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire [31:0] x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_rPort_1_output_0; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_sEn_2; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_sDone_2; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_rPort_1_output_0; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_sEn_1; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_sDone_1; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x556_tmp_2_sEn_3; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x556_tmp_2_sDone_3; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x735_rd_x595; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x596_reg_sEn_1; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x596_reg_sDone_1; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire [63:0] x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_11_cycs; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire [63:0] x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_11_iters; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire [63:0] x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_12_cycs; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire [63:0] x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_12_iters; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire [63:0] x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_13_cycs; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire [63:0] x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_13_iters; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_done; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_baseEn; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smSelectsOut_0; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smSelectsOut_1; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_rr; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire [31:0] x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_ret_number; // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
  wire  x623_inr_UnitPipe_sm_clock; // @[sm_x623_inr_UnitPipe.scala 34:18:@67730.4]
  wire  x623_inr_UnitPipe_sm_reset; // @[sm_x623_inr_UnitPipe.scala 34:18:@67730.4]
  wire  x623_inr_UnitPipe_sm_io_enable; // @[sm_x623_inr_UnitPipe.scala 34:18:@67730.4]
  wire  x623_inr_UnitPipe_sm_io_done; // @[sm_x623_inr_UnitPipe.scala 34:18:@67730.4]
  wire  x623_inr_UnitPipe_sm_io_doneLatch; // @[sm_x623_inr_UnitPipe.scala 34:18:@67730.4]
  wire  x623_inr_UnitPipe_sm_io_ctrDone; // @[sm_x623_inr_UnitPipe.scala 34:18:@67730.4]
  wire  x623_inr_UnitPipe_sm_io_datapathEn; // @[sm_x623_inr_UnitPipe.scala 34:18:@67730.4]
  wire  x623_inr_UnitPipe_sm_io_ctrInc; // @[sm_x623_inr_UnitPipe.scala 34:18:@67730.4]
  wire  x623_inr_UnitPipe_sm_io_parentAck; // @[sm_x623_inr_UnitPipe.scala 34:18:@67730.4]
  wire  x623_inr_UnitPipe_sm_io_backpressure; // @[sm_x623_inr_UnitPipe.scala 34:18:@67730.4]
  wire  x623_inr_UnitPipe_sm_io_break; // @[sm_x623_inr_UnitPipe.scala 34:18:@67730.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@67763.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@67763.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@67763.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@67763.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@67763.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@67773.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@67773.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@67773.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@67773.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@67773.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@67809.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@67809.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@67809.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@67809.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@67809.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@67817.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@67817.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@67817.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@67817.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@67817.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_clock; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_reset; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_4; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_4; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_4; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_4; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_4; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_4; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire [31:0] x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_wPort_0_data_0; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_wPort_0_en_0; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_sEn_0; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_sDone_0; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire [31:0] x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x621_inr_Switch_number; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_4; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_4; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_4; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_4; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire [63:0] x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_instrctrs_14_cycs; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire [63:0] x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_instrctrs_14_iters; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_done; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_baseEn; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_break; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_rr; // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
  wire  x625_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@68366.4]
  wire  x625_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@68366.4]
  wire  x625_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@68366.4]
  wire  x625_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@68366.4]
  wire [3:0] x625_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@68366.4]
  wire  x625_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@68366.4]
  wire  x625_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@68366.4]
  wire  x639_inr_Foreach_sm_clock; // @[sm_x639_inr_Foreach.scala 33:18:@68419.4]
  wire  x639_inr_Foreach_sm_reset; // @[sm_x639_inr_Foreach.scala 33:18:@68419.4]
  wire  x639_inr_Foreach_sm_io_enable; // @[sm_x639_inr_Foreach.scala 33:18:@68419.4]
  wire  x639_inr_Foreach_sm_io_done; // @[sm_x639_inr_Foreach.scala 33:18:@68419.4]
  wire  x639_inr_Foreach_sm_io_rst; // @[sm_x639_inr_Foreach.scala 33:18:@68419.4]
  wire  x639_inr_Foreach_sm_io_ctrDone; // @[sm_x639_inr_Foreach.scala 33:18:@68419.4]
  wire  x639_inr_Foreach_sm_io_datapathEn; // @[sm_x639_inr_Foreach.scala 33:18:@68419.4]
  wire  x639_inr_Foreach_sm_io_ctrInc; // @[sm_x639_inr_Foreach.scala 33:18:@68419.4]
  wire  x639_inr_Foreach_sm_io_ctrRst; // @[sm_x639_inr_Foreach.scala 33:18:@68419.4]
  wire  x639_inr_Foreach_sm_io_parentAck; // @[sm_x639_inr_Foreach.scala 33:18:@68419.4]
  wire  x639_inr_Foreach_sm_io_backpressure; // @[sm_x639_inr_Foreach.scala 33:18:@68419.4]
  wire  x639_inr_Foreach_sm_io_break; // @[sm_x639_inr_Foreach.scala 33:18:@68419.4]
  wire  x639_inr_Foreach_iiCtr_clock; // @[sm_x639_inr_Foreach.scala 34:21:@68444.4]
  wire  x639_inr_Foreach_iiCtr_reset; // @[sm_x639_inr_Foreach.scala 34:21:@68444.4]
  wire  x639_inr_Foreach_iiCtr_io_input_enable; // @[sm_x639_inr_Foreach.scala 34:21:@68444.4]
  wire  x639_inr_Foreach_iiCtr_io_input_reset; // @[sm_x639_inr_Foreach.scala 34:21:@68444.4]
  wire  x639_inr_Foreach_iiCtr_io_output_issue; // @[sm_x639_inr_Foreach.scala 34:21:@68444.4]
  wire  x639_inr_Foreach_iiCtr_io_output_done; // @[sm_x639_inr_Foreach.scala 34:21:@68444.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@68448.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@68448.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@68448.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@68448.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@68448.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@68457.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@68457.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@68457.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@68457.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@68457.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@68467.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@68467.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@68467.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@68467.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@68467.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@68509.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@68509.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@68509.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@68509.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@68509.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@68517.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@68517.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@68517.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@68517.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@68517.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_clock; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_reset; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire [1:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_ofs_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire [31:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_data_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_en_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_sEn_5; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_sDone_5; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire [1:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_ofs_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire [31:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_data_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_en_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_sEn_5; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_sDone_5; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire [1:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_ofs_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire [31:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_data_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_en_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_5; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_5; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_b552; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_rPort_0_en_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire [31:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_rPort_0_output_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_sEn_1; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_sDone_1; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire [1:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_ofs_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_en_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire [31:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_output_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire [1:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_ofs_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire [31:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_data_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_en_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_sEn_5; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_sDone_5; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire [1:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_ofs_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire [31:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_data_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_en_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_sEn_5; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_sDone_5; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_b543; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire [63:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_instrctrs_15_cycs; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire [63:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_instrctrs_15_iters; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_done; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_iiIssue; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire [31:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_rr; // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
  wire  x652_inr_Foreach_sm_clock; // @[sm_x652_inr_Foreach.scala 35:18:@69143.4]
  wire  x652_inr_Foreach_sm_reset; // @[sm_x652_inr_Foreach.scala 35:18:@69143.4]
  wire  x652_inr_Foreach_sm_io_enable; // @[sm_x652_inr_Foreach.scala 35:18:@69143.4]
  wire  x652_inr_Foreach_sm_io_done; // @[sm_x652_inr_Foreach.scala 35:18:@69143.4]
  wire  x652_inr_Foreach_sm_io_doneLatch; // @[sm_x652_inr_Foreach.scala 35:18:@69143.4]
  wire  x652_inr_Foreach_sm_io_ctrDone; // @[sm_x652_inr_Foreach.scala 35:18:@69143.4]
  wire  x652_inr_Foreach_sm_io_datapathEn; // @[sm_x652_inr_Foreach.scala 35:18:@69143.4]
  wire  x652_inr_Foreach_sm_io_ctrInc; // @[sm_x652_inr_Foreach.scala 35:18:@69143.4]
  wire  x652_inr_Foreach_sm_io_ctrRst; // @[sm_x652_inr_Foreach.scala 35:18:@69143.4]
  wire  x652_inr_Foreach_sm_io_parentAck; // @[sm_x652_inr_Foreach.scala 35:18:@69143.4]
  wire  x652_inr_Foreach_sm_io_backpressure; // @[sm_x652_inr_Foreach.scala 35:18:@69143.4]
  wire  x652_inr_Foreach_sm_io_break; // @[sm_x652_inr_Foreach.scala 35:18:@69143.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@69172.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@69172.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@69172.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@69172.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@69172.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@69181.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@69181.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@69181.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@69181.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@69181.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@69191.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@69191.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@69191.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@69191.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@69191.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@69232.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@69232.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@69232.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@69232.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@69232.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@69240.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@69240.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@69240.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@69240.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@69240.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_clock; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_reset; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire [31:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_b550_number; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire [1:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_ofs_0; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_en_0; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire [31:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_output_0; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_6; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_6; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire [1:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_ofs_0; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire [31:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_data_0; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_en_0; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire [1:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_ofs_0; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_en_0; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire [31:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_output_0; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire [1:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_ofs_0; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire [31:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_data_0; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_en_0; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_b543; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire [63:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_instrctrs_16_cycs; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire [63:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_instrctrs_16_iters; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_done; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire [31:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_rr; // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@69577.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@69577.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@69577.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@69577.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@69577.4]
  wire  _T_786; // @[package.scala 100:49:@64030.4]
  reg  _T_789; // @[package.scala 48:56:@64031.4]
  reg [31:0] _RAND_0;
  wire  b552; // @[sm_x653_outr_Reduce.scala 100:18:@64190.4]
  wire  b552_chain_read_1; // @[sm_x653_outr_Reduce.scala 103:61:@64264.4]
  wire  b552_chain_read_2; // @[sm_x653_outr_Reduce.scala 104:61:@64265.4]
  wire  b552_chain_read_4; // @[sm_x653_outr_Reduce.scala 106:61:@64267.4]
  wire  b552_chain_read_5; // @[sm_x653_outr_Reduce.scala 107:61:@64268.4]
  wire  _T_911; // @[package.scala 96:25:@64594.4 package.scala 96:25:@64595.4]
  wire  _T_915; // @[package.scala 96:25:@64603.4 package.scala 96:25:@64604.4]
  wire  _T_919; // @[package.scala 96:25:@64613.4 package.scala 96:25:@64614.4]
  wire  x579_inr_Foreach_mySignalsIn_mask; // @[sm_x653_outr_Reduce.scala 126:81:@64627.4]
  wire  _T_936; // @[package.scala 96:25:@64655.4 package.scala 96:25:@64656.4]
  wire  _T_942; // @[package.scala 96:25:@64663.4 package.scala 96:25:@64664.4]
  wire  _T_945; // @[SpatialBlocks.scala 137:99:@64666.4]
  wire  _T_947; // @[SpatialBlocks.scala 156:36:@64675.4]
  wire  _T_948; // @[SpatialBlocks.scala 156:78:@64676.4]
  wire  _T_1016; // @[package.scala 100:49:@65339.4]
  reg  _T_1019; // @[package.scala 48:56:@65340.4]
  reg [31:0] _RAND_1;
  wire  _T_1022; // @[package.scala 96:25:@65349.4 package.scala 96:25:@65350.4]
  wire  _T_1026; // @[package.scala 96:25:@65359.4 package.scala 96:25:@65360.4]
  wire  x593_inr_UnitPipe_mySignalsIn_mask; // @[sm_x653_outr_Reduce.scala 138:60:@65372.4]
  wire  _T_1043; // @[package.scala 96:25:@65395.4 package.scala 96:25:@65396.4]
  wire  _T_1049; // @[package.scala 96:25:@65403.4 package.scala 96:25:@65404.4]
  wire  _T_1052; // @[SpatialBlocks.scala 137:99:@65406.4]
  wire  _T_1123; // @[package.scala 100:49:@66132.4]
  reg  _T_1126; // @[package.scala 48:56:@66133.4]
  reg [31:0] _RAND_2;
  wire  _T_1129; // @[package.scala 96:25:@66142.4 package.scala 96:25:@66143.4]
  wire  _T_1133; // @[package.scala 96:25:@66152.4 package.scala 96:25:@66153.4]
  wire  x605_inr_UnitPipe_mySignalsIn_mask; // @[sm_x653_outr_Reduce.scala 152:60:@66165.4]
  wire  _T_1150; // @[package.scala 96:25:@66188.4 package.scala 96:25:@66189.4]
  wire  _T_1156; // @[package.scala 96:25:@66196.4 package.scala 96:25:@66197.4]
  wire  _T_1159; // @[SpatialBlocks.scala 137:99:@66199.4]
  wire  _T_1257; // @[package.scala 96:25:@66965.4 package.scala 96:25:@66966.4]
  wire  _T_1261; // @[package.scala 96:25:@66975.4 package.scala 96:25:@66976.4]
  wire  _T_1279; // @[package.scala 96:25:@67017.4 package.scala 96:25:@67018.4]
  wire  _T_1285; // @[package.scala 96:25:@67025.4 package.scala 96:25:@67026.4]
  wire  _T_1288; // @[SpatialBlocks.scala 137:99:@67028.4]
  wire  _T_1356; // @[package.scala 100:49:@67758.4]
  reg  _T_1359; // @[package.scala 48:56:@67759.4]
  reg [31:0] _RAND_3;
  wire  _T_1362; // @[package.scala 96:25:@67768.4 package.scala 96:25:@67769.4]
  wire  _T_1366; // @[package.scala 96:25:@67778.4 package.scala 96:25:@67779.4]
  wire  x623_inr_UnitPipe_mySignalsIn_mask; // @[sm_x653_outr_Reduce.scala 188:60:@67791.4]
  wire  _T_1383; // @[package.scala 96:25:@67814.4 package.scala 96:25:@67815.4]
  wire  _T_1389; // @[package.scala 96:25:@67822.4 package.scala 96:25:@67823.4]
  wire  _T_1392; // @[SpatialBlocks.scala 137:99:@67825.4]
  wire  _T_1464; // @[package.scala 96:25:@68453.4 package.scala 96:25:@68454.4]
  wire  _T_1468; // @[package.scala 96:25:@68462.4 package.scala 96:25:@68463.4]
  wire  _T_1472; // @[package.scala 96:25:@68472.4 package.scala 96:25:@68473.4]
  wire  x639_inr_Foreach_mySignalsIn_mask; // @[sm_x653_outr_Reduce.scala 203:94:@68486.4]
  wire  _T_1489; // @[package.scala 96:25:@68514.4 package.scala 96:25:@68515.4]
  wire  _T_1495; // @[package.scala 96:25:@68522.4 package.scala 96:25:@68523.4]
  wire  _T_1498; // @[SpatialBlocks.scala 137:99:@68525.4]
  wire  _T_1500; // @[SpatialBlocks.scala 156:36:@68534.4]
  wire  _T_1501; // @[SpatialBlocks.scala 156:78:@68535.4]
  wire  _T_1504; // @[SpatialBlocks.scala 157:128:@68541.4]
  wire  x639_inr_Foreach_mySignalsIn_iiDone; // @[SpatialBlocks.scala 157:126:@68542.4]
  wire  _T_1570; // @[package.scala 96:25:@69177.4 package.scala 96:25:@69178.4]
  wire  _T_1574; // @[package.scala 96:25:@69186.4 package.scala 96:25:@69187.4]
  wire  _T_1578; // @[package.scala 96:25:@69196.4 package.scala 96:25:@69197.4]
  wire  _T_1595; // @[package.scala 96:25:@69237.4 package.scala 96:25:@69238.4]
  wire  _T_1601; // @[package.scala 96:25:@69245.4 package.scala 96:25:@69246.4]
  wire  _T_1604; // @[SpatialBlocks.scala 137:99:@69248.4]
  wire  _T_1606; // @[SpatialBlocks.scala 156:36:@69257.4]
  wire  _T_1607; // @[SpatialBlocks.scala 156:78:@69258.4]
  wire  _T_1619; // @[package.scala 96:25:@69582.4 package.scala 96:25:@69583.4]
  InstrumentationCounter cycles_x653_outr_Reduce ( // @[sm_x653_outr_Reduce.scala 86:43:@64023.4]
    .clock(cycles_x653_outr_Reduce_clock),
    .reset(cycles_x653_outr_Reduce_reset),
    .io_enable(cycles_x653_outr_Reduce_io_enable),
    .io_count(cycles_x653_outr_Reduce_io_count)
  );
  InstrumentationCounter iters_x653_outr_Reduce ( // @[sm_x653_outr_Reduce.scala 87:42:@64026.4]
    .clock(iters_x653_outr_Reduce_clock),
    .reset(iters_x653_outr_Reduce_reset),
    .io_enable(iters_x653_outr_Reduce_io_enable),
    .io_count(iters_x653_outr_Reduce_io_count)
  );
  _ _ ( // @[Math.scala 720:24:@64043.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  b550_chain b550_chain ( // @[sm_x653_outr_Reduce.scala 92:30:@64051.4]
    .clock(b550_chain_clock),
    .reset(b550_chain_reset),
    .io_rPort_5_output_0(b550_chain_io_rPort_5_output_0),
    .io_rPort_4_output_0(b550_chain_io_rPort_4_output_0),
    .io_rPort_3_output_0(b550_chain_io_rPort_3_output_0),
    .io_rPort_2_output_0(b550_chain_io_rPort_2_output_0),
    .io_rPort_1_output_0(b550_chain_io_rPort_1_output_0),
    .io_rPort_0_output_0(b550_chain_io_rPort_0_output_0),
    .io_wPort_0_data_0(b550_chain_io_wPort_0_data_0),
    .io_wPort_0_reset(b550_chain_io_wPort_0_reset),
    .io_wPort_0_en_0(b550_chain_io_wPort_0_en_0),
    .io_sEn_0(b550_chain_io_sEn_0),
    .io_sEn_1(b550_chain_io_sEn_1),
    .io_sEn_2(b550_chain_io_sEn_2),
    .io_sEn_3(b550_chain_io_sEn_3),
    .io_sEn_4(b550_chain_io_sEn_4),
    .io_sEn_5(b550_chain_io_sEn_5),
    .io_sEn_6(b550_chain_io_sEn_6),
    .io_sDone_0(b550_chain_io_sDone_0),
    .io_sDone_1(b550_chain_io_sDone_1),
    .io_sDone_2(b550_chain_io_sDone_2),
    .io_sDone_3(b550_chain_io_sDone_3),
    .io_sDone_4(b550_chain_io_sDone_4),
    .io_sDone_5(b550_chain_io_sDone_5),
    .io_sDone_6(b550_chain_io_sDone_6)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@64115.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  _ __1 ( // @[Math.scala 720:24:@64127.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  _ __2 ( // @[Math.scala 720:24:@64138.4]
    .io_b(__2_io_b),
    .io_result(__2_io_result)
  );
  _ __3 ( // @[Math.scala 720:24:@64149.4]
    .io_b(__3_io_b),
    .io_result(__3_io_result)
  );
  _ __4 ( // @[Math.scala 720:24:@64160.4]
    .io_b(__4_io_b),
    .io_result(__4_io_result)
  );
  _ __5 ( // @[Math.scala 720:24:@64171.4]
    .io_b(__5_io_b),
    .io_result(__5_io_result)
  );
  _ __6 ( // @[Math.scala 720:24:@64182.4]
    .io_b(__6_io_b),
    .io_result(__6_io_result)
  );
  b552_chain b552_chain ( // @[sm_x653_outr_Reduce.scala 101:30:@64191.4]
    .clock(b552_chain_clock),
    .reset(b552_chain_reset),
    .io_rPort_4_output_0(b552_chain_io_rPort_4_output_0),
    .io_rPort_3_output_0(b552_chain_io_rPort_3_output_0),
    .io_rPort_1_output_0(b552_chain_io_rPort_1_output_0),
    .io_rPort_0_output_0(b552_chain_io_rPort_0_output_0),
    .io_wPort_0_data_0(b552_chain_io_wPort_0_data_0),
    .io_wPort_0_reset(b552_chain_io_wPort_0_reset),
    .io_wPort_0_en_0(b552_chain_io_wPort_0_en_0),
    .io_sEn_0(b552_chain_io_sEn_0),
    .io_sEn_1(b552_chain_io_sEn_1),
    .io_sEn_2(b552_chain_io_sEn_2),
    .io_sEn_3(b552_chain_io_sEn_3),
    .io_sEn_4(b552_chain_io_sEn_4),
    .io_sEn_5(b552_chain_io_sEn_5),
    .io_sEn_6(b552_chain_io_sEn_6),
    .io_sDone_0(b552_chain_io_sDone_0),
    .io_sDone_1(b552_chain_io_sDone_1),
    .io_sDone_2(b552_chain_io_sDone_2),
    .io_sDone_3(b552_chain_io_sDone_3),
    .io_sDone_4(b552_chain_io_sDone_4),
    .io_sDone_5(b552_chain_io_sDone_5),
    .io_sDone_6(b552_chain_io_sDone_6)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@64255.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x554_tmp_0 x554_tmp_0 ( // @[m_x554_tmp_0.scala 28:22:@64270.4]
    .clock(x554_tmp_0_clock),
    .reset(x554_tmp_0_reset),
    .io_rPort_0_ofs_0(x554_tmp_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x554_tmp_0_io_rPort_0_en_0),
    .io_rPort_0_output_0(x554_tmp_0_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(x554_tmp_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x554_tmp_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x554_tmp_0_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(x554_tmp_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x554_tmp_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x554_tmp_0_io_wPort_0_en_0),
    .io_sEn_0(x554_tmp_0_io_sEn_0),
    .io_sEn_1(x554_tmp_0_io_sEn_1),
    .io_sEn_2(x554_tmp_0_io_sEn_2),
    .io_sEn_3(x554_tmp_0_io_sEn_3),
    .io_sEn_4(x554_tmp_0_io_sEn_4),
    .io_sEn_5(x554_tmp_0_io_sEn_5),
    .io_sDone_0(x554_tmp_0_io_sDone_0),
    .io_sDone_1(x554_tmp_0_io_sDone_1),
    .io_sDone_2(x554_tmp_0_io_sDone_2),
    .io_sDone_3(x554_tmp_0_io_sDone_3),
    .io_sDone_4(x554_tmp_0_io_sDone_4),
    .io_sDone_5(x554_tmp_0_io_sDone_5)
  );
  x554_tmp_0 x555_tmp_1 ( // @[m_x555_tmp_1.scala 28:22:@64317.4]
    .clock(x555_tmp_1_clock),
    .reset(x555_tmp_1_reset),
    .io_rPort_0_ofs_0(x555_tmp_1_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x555_tmp_1_io_rPort_0_en_0),
    .io_rPort_0_output_0(x555_tmp_1_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(x555_tmp_1_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x555_tmp_1_io_wPort_1_data_0),
    .io_wPort_1_en_0(x555_tmp_1_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(x555_tmp_1_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x555_tmp_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(x555_tmp_1_io_wPort_0_en_0),
    .io_sEn_0(x555_tmp_1_io_sEn_0),
    .io_sEn_1(x555_tmp_1_io_sEn_1),
    .io_sEn_2(x555_tmp_1_io_sEn_2),
    .io_sEn_3(x555_tmp_1_io_sEn_3),
    .io_sEn_4(x555_tmp_1_io_sEn_4),
    .io_sEn_5(x555_tmp_1_io_sEn_5),
    .io_sDone_0(x555_tmp_1_io_sDone_0),
    .io_sDone_1(x555_tmp_1_io_sDone_1),
    .io_sDone_2(x555_tmp_1_io_sDone_2),
    .io_sDone_3(x555_tmp_1_io_sDone_3),
    .io_sDone_4(x555_tmp_1_io_sDone_4),
    .io_sDone_5(x555_tmp_1_io_sDone_5)
  );
  x554_tmp_0 x556_tmp_2 ( // @[m_x556_tmp_2.scala 28:22:@64364.4]
    .clock(x556_tmp_2_clock),
    .reset(x556_tmp_2_reset),
    .io_rPort_0_ofs_0(x556_tmp_2_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x556_tmp_2_io_rPort_0_en_0),
    .io_rPort_0_output_0(x556_tmp_2_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(x556_tmp_2_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x556_tmp_2_io_wPort_1_data_0),
    .io_wPort_1_en_0(x556_tmp_2_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(x556_tmp_2_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x556_tmp_2_io_wPort_0_data_0),
    .io_wPort_0_en_0(x556_tmp_2_io_wPort_0_en_0),
    .io_sEn_0(x556_tmp_2_io_sEn_0),
    .io_sEn_1(x556_tmp_2_io_sEn_1),
    .io_sEn_2(x556_tmp_2_io_sEn_2),
    .io_sEn_3(x556_tmp_2_io_sEn_3),
    .io_sEn_4(x556_tmp_2_io_sEn_4),
    .io_sEn_5(x556_tmp_2_io_sEn_5),
    .io_sDone_0(x556_tmp_2_io_sDone_0),
    .io_sDone_1(x556_tmp_2_io_sDone_1),
    .io_sDone_2(x556_tmp_2_io_sDone_2),
    .io_sDone_3(x556_tmp_2_io_sDone_3),
    .io_sDone_4(x556_tmp_2_io_sDone_4),
    .io_sDone_5(x556_tmp_2_io_sDone_5)
  );
  x557_tmp_3 x557_tmp_3 ( // @[m_x557_tmp_3.scala 28:22:@64411.4]
    .clock(x557_tmp_3_clock),
    .reset(x557_tmp_3_reset),
    .io_rPort_0_ofs_0(x557_tmp_3_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x557_tmp_3_io_rPort_0_en_0),
    .io_rPort_0_output_0(x557_tmp_3_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(x557_tmp_3_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x557_tmp_3_io_wPort_1_data_0),
    .io_wPort_1_en_0(x557_tmp_3_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(x557_tmp_3_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x557_tmp_3_io_wPort_0_data_0),
    .io_wPort_0_en_0(x557_tmp_3_io_wPort_0_en_0),
    .io_sEn_0(x557_tmp_3_io_sEn_0),
    .io_sEn_1(x557_tmp_3_io_sEn_1),
    .io_sEn_2(x557_tmp_3_io_sEn_2),
    .io_sEn_3(x557_tmp_3_io_sEn_3),
    .io_sEn_4(x557_tmp_3_io_sEn_4),
    .io_sEn_5(x557_tmp_3_io_sEn_5),
    .io_sDone_0(x557_tmp_3_io_sDone_0),
    .io_sDone_1(x557_tmp_3_io_sDone_1),
    .io_sDone_2(x557_tmp_3_io_sDone_2),
    .io_sDone_3(x557_tmp_3_io_sDone_3),
    .io_sDone_4(x557_tmp_3_io_sDone_4),
    .io_sDone_5(x557_tmp_3_io_sDone_5)
  );
  x558_tmp_4 x558_tmp_4 ( // @[m_x558_tmp_4.scala 28:22:@64458.4]
    .clock(x558_tmp_4_clock),
    .reset(x558_tmp_4_reset),
    .io_rPort_0_ofs_0(x558_tmp_4_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x558_tmp_4_io_rPort_0_en_0),
    .io_rPort_0_output_0(x558_tmp_4_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(x558_tmp_4_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x558_tmp_4_io_wPort_1_data_0),
    .io_wPort_1_en_0(x558_tmp_4_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(x558_tmp_4_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x558_tmp_4_io_wPort_0_data_0),
    .io_wPort_0_en_0(x558_tmp_4_io_wPort_0_en_0),
    .io_sEn_0(x558_tmp_4_io_sEn_0),
    .io_sEn_1(x558_tmp_4_io_sEn_1),
    .io_sEn_2(x558_tmp_4_io_sEn_2),
    .io_sEn_3(x558_tmp_4_io_sEn_3),
    .io_sEn_4(x558_tmp_4_io_sEn_4),
    .io_sEn_5(x558_tmp_4_io_sEn_5),
    .io_sEn_6(x558_tmp_4_io_sEn_6),
    .io_sDone_0(x558_tmp_4_io_sDone_0),
    .io_sDone_1(x558_tmp_4_io_sDone_1),
    .io_sDone_2(x558_tmp_4_io_sDone_2),
    .io_sDone_3(x558_tmp_4_io_sDone_3),
    .io_sDone_4(x558_tmp_4_io_sDone_4),
    .io_sDone_5(x558_tmp_4_io_sDone_5),
    .io_sDone_6(x558_tmp_4_io_sDone_6)
  );
  x549_ctrchain x560_ctrchain ( // @[SpatialBlocks.scala 37:22:@64507.4]
    .clock(x560_ctrchain_clock),
    .reset(x560_ctrchain_reset),
    .io_input_reset(x560_ctrchain_io_input_reset),
    .io_input_enable(x560_ctrchain_io_input_enable),
    .io_output_counts_0(x560_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x560_ctrchain_io_output_oobs_0),
    .io_output_done(x560_ctrchain_io_output_done)
  );
  x579_inr_Foreach_sm x579_inr_Foreach_sm ( // @[sm_x579_inr_Foreach.scala 35:18:@64560.4]
    .clock(x579_inr_Foreach_sm_clock),
    .reset(x579_inr_Foreach_sm_reset),
    .io_enable(x579_inr_Foreach_sm_io_enable),
    .io_done(x579_inr_Foreach_sm_io_done),
    .io_ctrDone(x579_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x579_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x579_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x579_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x579_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x579_inr_Foreach_sm_io_backpressure),
    .io_break(x579_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@64589.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@64598.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@64608.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@64650.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@64658.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1 x579_inr_Foreach_kernelx579_inr_Foreach_concrete1 ( // @[sm_x579_inr_Foreach.scala 187:24:@64692.4]
    .clock(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_clock),
    .reset(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_reset),
    .io_in_x555_tmp_1_wPort_0_ofs_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_ofs_0),
    .io_in_x555_tmp_1_wPort_0_data_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_data_0),
    .io_in_x555_tmp_1_wPort_0_en_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_en_0),
    .io_in_x555_tmp_1_sEn_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_sEn_0),
    .io_in_x555_tmp_1_sDone_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_sDone_0),
    .io_in_b550_number(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b550_number),
    .io_in_x472_A_sram_1_rPort_0_ofs_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0),
    .io_in_x472_A_sram_1_rPort_0_en_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_en_0),
    .io_in_x472_A_sram_1_rPort_0_output_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_output_0),
    .io_in_b542_number(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b542_number),
    .io_in_x471_A_sram_0_rPort_0_ofs_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0),
    .io_in_x471_A_sram_0_rPort_0_en_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_en_0),
    .io_in_x471_A_sram_0_rPort_0_output_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_output_0),
    .io_in_x554_tmp_0_wPort_0_ofs_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_ofs_0),
    .io_in_x554_tmp_0_wPort_0_data_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_data_0),
    .io_in_x554_tmp_0_wPort_0_en_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_en_0),
    .io_in_x554_tmp_0_sEn_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_sEn_0),
    .io_in_x554_tmp_0_sDone_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_sDone_0),
    .io_in_x558_tmp_4_wPort_0_ofs_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_ofs_0),
    .io_in_x558_tmp_4_wPort_0_data_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_data_0),
    .io_in_x558_tmp_4_wPort_0_en_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_en_0),
    .io_in_x558_tmp_4_sEn_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_0),
    .io_in_x558_tmp_4_sDone_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_0),
    .io_in_b552(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b552),
    .io_in_x557_tmp_3_wPort_0_ofs_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_ofs_0),
    .io_in_x557_tmp_3_wPort_0_data_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_data_0),
    .io_in_x557_tmp_3_wPort_0_en_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_en_0),
    .io_in_x557_tmp_3_sEn_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_sEn_0),
    .io_in_x557_tmp_3_sDone_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_sDone_0),
    .io_in_x556_tmp_2_wPort_0_ofs_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_ofs_0),
    .io_in_x556_tmp_2_wPort_0_data_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_data_0),
    .io_in_x556_tmp_2_wPort_0_en_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_en_0),
    .io_in_x556_tmp_2_sEn_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_sEn_0),
    .io_in_x556_tmp_2_sDone_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_sDone_0),
    .io_in_b543(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b543),
    .io_in_instrctrs_8_cycs(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_instrctrs_8_cycs),
    .io_in_instrctrs_8_iters(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_instrctrs_8_iters),
    .io_sigsIn_done(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_datapathEn(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_rr)
  );
  x580_r_0 x580_r_0 ( // @[m_x580_r_0.scala 28:22:@65236.4]
    .clock(x580_r_0_clock),
    .reset(x580_r_0_reset),
    .io_rPort_1_en_0(x580_r_0_io_rPort_1_en_0),
    .io_rPort_1_output_0(x580_r_0_io_rPort_1_output_0),
    .io_rPort_0_en_0(x580_r_0_io_rPort_0_en_0),
    .io_rPort_0_output_0(x580_r_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(x580_r_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x580_r_0_io_wPort_0_en_0),
    .io_sEn_0(x580_r_0_io_sEn_0),
    .io_sEn_1(x580_r_0_io_sEn_1),
    .io_sEn_2(x580_r_0_io_sEn_2),
    .io_sDone_0(x580_r_0_io_sDone_0),
    .io_sDone_1(x580_r_0_io_sDone_1),
    .io_sDone_2(x580_r_0_io_sDone_2)
  );
  x593_inr_UnitPipe_sm x593_inr_UnitPipe_sm ( // @[sm_x593_inr_UnitPipe.scala 33:18:@65311.4]
    .clock(x593_inr_UnitPipe_sm_clock),
    .reset(x593_inr_UnitPipe_sm_reset),
    .io_enable(x593_inr_UnitPipe_sm_io_enable),
    .io_done(x593_inr_UnitPipe_sm_io_done),
    .io_ctrDone(x593_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x593_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x593_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x593_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x593_inr_UnitPipe_sm_io_backpressure),
    .io_break(x593_inr_UnitPipe_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@65344.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@65354.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@65390.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@65398.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1 x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1 ( // @[sm_x593_inr_UnitPipe.scala 141:24:@65427.4]
    .clock(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_clock),
    .reset(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_reset),
    .io_in_x555_tmp_1_rPort_0_en_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_rPort_0_en_0),
    .io_in_x555_tmp_1_rPort_0_output_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_rPort_0_output_0),
    .io_in_x555_tmp_1_sEn_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_1),
    .io_in_x555_tmp_1_sDone_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_1),
    .io_in_x554_tmp_0_rPort_0_en_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_rPort_0_en_0),
    .io_in_x554_tmp_0_rPort_0_output_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_rPort_0_output_0),
    .io_in_x554_tmp_0_sEn_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_1),
    .io_in_x554_tmp_0_sDone_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_1),
    .io_in_x558_tmp_4_sEn_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_1),
    .io_in_x558_tmp_4_sDone_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_1),
    .io_in_x557_tmp_3_sEn_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_1),
    .io_in_x557_tmp_3_sDone_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_1),
    .io_in_x580_r_0_wPort_0_data_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_wPort_0_data_0),
    .io_in_x580_r_0_wPort_0_en_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_wPort_0_en_0),
    .io_in_x580_r_0_sEn_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_sEn_0),
    .io_in_x580_r_0_sDone_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_sDone_0),
    .io_in_x556_tmp_2_rPort_0_en_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_rPort_0_en_0),
    .io_in_x556_tmp_2_rPort_0_output_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_rPort_0_output_0),
    .io_in_x556_tmp_2_sEn_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_1),
    .io_in_x556_tmp_2_sDone_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_1),
    .io_in_instrctrs_9_cycs(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_instrctrs_9_cycs),
    .io_in_instrctrs_9_iters(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_instrctrs_9_iters),
    .io_sigsIn_done(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_done),
    .io_sigsIn_datapathEn(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_break),
    .io_rr(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_rr)
  );
  x594_force_0 x594_force_0 ( // @[m_x594_force_0.scala 27:22:@65971.4]
    .clock(x594_force_0_clock),
    .reset(x594_force_0_reset),
    .io_rPort_0_en_0(x594_force_0_io_rPort_0_en_0),
    .io_rPort_0_output_0(x594_force_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(x594_force_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x594_force_0_io_wPort_0_en_0),
    .io_sEn_0(x594_force_0_io_sEn_0),
    .io_sEn_1(x594_force_0_io_sEn_1),
    .io_sDone_0(x594_force_0_io_sDone_0),
    .io_sDone_1(x594_force_0_io_sDone_1)
  );
  x595_reg x595_reg ( // @[m_x595_reg.scala 28:22:@66001.4]
    .clock(x595_reg_clock),
    .reset(x595_reg_reset),
    .io_rPort_1_output_0(x595_reg_io_rPort_1_output_0),
    .io_rPort_0_output_0(x595_reg_io_rPort_0_output_0),
    .io_wPort_0_data_0(x595_reg_io_wPort_0_data_0),
    .io_wPort_0_reset(x595_reg_io_wPort_0_reset),
    .io_wPort_0_en_0(x595_reg_io_wPort_0_en_0),
    .io_sEn_0(x595_reg_io_sEn_0),
    .io_sEn_1(x595_reg_io_sEn_1),
    .io_sDone_0(x595_reg_io_sDone_0),
    .io_sDone_1(x595_reg_io_sDone_1)
  );
  x596_reg x596_reg ( // @[m_x596_reg.scala 27:22:@66038.4]
    .clock(x596_reg_clock),
    .reset(x596_reg_reset),
    .io_rPort_0_output_0(x596_reg_io_rPort_0_output_0),
    .io_wPort_0_data_0(x596_reg_io_wPort_0_data_0),
    .io_wPort_0_reset(x596_reg_io_wPort_0_reset),
    .io_wPort_0_en_0(x596_reg_io_wPort_0_en_0),
    .io_sEn_0(x596_reg_io_sEn_0),
    .io_sEn_1(x596_reg_io_sEn_1),
    .io_sDone_0(x596_reg_io_sDone_0),
    .io_sDone_1(x596_reg_io_sDone_1)
  );
  x536_inr_Foreach_sm x605_inr_UnitPipe_sm ( // @[sm_x605_inr_UnitPipe.scala 33:18:@66104.4]
    .clock(x605_inr_UnitPipe_sm_clock),
    .reset(x605_inr_UnitPipe_sm_reset),
    .io_enable(x605_inr_UnitPipe_sm_io_enable),
    .io_done(x605_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x605_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x605_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x605_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x605_inr_UnitPipe_sm_io_ctrInc),
    .io_ctrRst(x605_inr_UnitPipe_sm_io_ctrRst),
    .io_parentAck(x605_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x605_inr_UnitPipe_sm_io_backpressure),
    .io_break(x605_inr_UnitPipe_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_11 ( // @[package.scala 93:22:@66137.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper RetimeWrapper_12 ( // @[package.scala 93:22:@66147.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 ( // @[package.scala 93:22:@66183.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@66191.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1 x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1 ( // @[sm_x605_inr_UnitPipe.scala 136:24:@66220.4]
    .clock(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_clock),
    .reset(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_reset),
    .io_in_x555_tmp_1_sEn_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_2),
    .io_in_x555_tmp_1_sDone_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_2),
    .io_in_x554_tmp_0_sEn_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_2),
    .io_in_x554_tmp_0_sDone_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_2),
    .io_in_x558_tmp_4_sEn_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_2),
    .io_in_x558_tmp_4_sDone_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_2),
    .io_in_x557_tmp_3_sEn_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_2),
    .io_in_x557_tmp_3_sDone_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_2),
    .io_in_x580_r_0_rPort_0_en_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_rPort_0_en_0),
    .io_in_x580_r_0_rPort_0_output_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_rPort_0_output_0),
    .io_in_x580_r_0_sEn_1(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_sEn_1),
    .io_in_x580_r_0_sDone_1(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_sDone_1),
    .io_in_x595_reg_wPort_0_data_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_data_0),
    .io_in_x595_reg_wPort_0_reset(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_reset),
    .io_in_x595_reg_wPort_0_en_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_en_0),
    .io_in_x595_reg_reset(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_reset),
    .io_in_x595_reg_sEn_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_sEn_0),
    .io_in_x595_reg_sDone_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_sDone_0),
    .io_in_x556_tmp_2_sEn_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_2),
    .io_in_x556_tmp_2_sDone_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_2),
    .io_in_x596_reg_wPort_0_data_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_data_0),
    .io_in_x596_reg_wPort_0_reset(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_reset),
    .io_in_x596_reg_wPort_0_en_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_en_0),
    .io_in_x596_reg_reset(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_reset),
    .io_in_x596_reg_sEn_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_sEn_0),
    .io_in_x596_reg_sDone_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_sDone_0),
    .io_in_instrctrs_10_cycs(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_instrctrs_10_cycs),
    .io_in_instrctrs_10_iters(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_instrctrs_10_iters),
    .io_sigsIn_done(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_done),
    .io_sigsIn_datapathEn(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_break),
    .io_rr(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_rr)
  );
  x621_inr_Switch_sm x621_inr_Switch_sm ( // @[sm_x621_inr_Switch.scala 33:18:@66923.4]
    .clock(x621_inr_Switch_sm_clock),
    .reset(x621_inr_Switch_sm_reset),
    .io_enable(x621_inr_Switch_sm_io_enable),
    .io_done(x621_inr_Switch_sm_io_done),
    .io_parentAck(x621_inr_Switch_sm_io_parentAck),
    .io_backpressure(x621_inr_Switch_sm_io_backpressure),
    .io_doneIn_0(x621_inr_Switch_sm_io_doneIn_0),
    .io_doneIn_1(x621_inr_Switch_sm_io_doneIn_1),
    .io_childAck_0(x621_inr_Switch_sm_io_childAck_0),
    .io_childAck_1(x621_inr_Switch_sm_io_childAck_1),
    .io_selectsIn_0(x621_inr_Switch_sm_io_selectsIn_0),
    .io_selectsIn_1(x621_inr_Switch_sm_io_selectsIn_1),
    .io_selectsOut_0(x621_inr_Switch_sm_io_selectsOut_0),
    .io_selectsOut_1(x621_inr_Switch_sm_io_selectsOut_1)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@66960.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 ( // @[package.scala 93:22:@66970.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper RetimeWrapper_17 ( // @[package.scala 93:22:@67012.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 ( // @[package.scala 93:22:@67020.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  x621_inr_Switch_kernelx621_inr_Switch_concrete1 x621_inr_Switch_kernelx621_inr_Switch_concrete1 ( // @[sm_x621_inr_Switch.scala 139:24:@67049.4]
    .clock(x621_inr_Switch_kernelx621_inr_Switch_concrete1_clock),
    .reset(x621_inr_Switch_kernelx621_inr_Switch_concrete1_reset),
    .io_in_x555_tmp_1_sEn_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x555_tmp_1_sEn_3),
    .io_in_x555_tmp_1_sDone_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x555_tmp_1_sDone_3),
    .io_in_x554_tmp_0_sEn_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x554_tmp_0_sEn_3),
    .io_in_x554_tmp_0_sDone_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x554_tmp_0_sDone_3),
    .io_in_x558_tmp_4_sEn_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x558_tmp_4_sEn_3),
    .io_in_x558_tmp_4_sDone_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x558_tmp_4_sDone_3),
    .io_in_x736_rd_x596(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x736_rd_x596),
    .io_in_x557_tmp_3_sEn_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x557_tmp_3_sEn_3),
    .io_in_x557_tmp_3_sDone_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x557_tmp_3_sDone_3),
    .io_in_x580_r_0_rPort_1_en_0(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_rPort_1_en_0),
    .io_in_x580_r_0_rPort_1_output_0(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_rPort_1_output_0),
    .io_in_x580_r_0_sEn_2(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_sEn_2),
    .io_in_x580_r_0_sDone_2(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_sDone_2),
    .io_in_x595_reg_rPort_1_output_0(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_rPort_1_output_0),
    .io_in_x595_reg_sEn_1(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_sEn_1),
    .io_in_x595_reg_sDone_1(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_sDone_1),
    .io_in_x556_tmp_2_sEn_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x556_tmp_2_sEn_3),
    .io_in_x556_tmp_2_sDone_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x556_tmp_2_sDone_3),
    .io_in_x735_rd_x595(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x735_rd_x595),
    .io_in_x596_reg_sEn_1(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x596_reg_sEn_1),
    .io_in_x596_reg_sDone_1(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x596_reg_sDone_1),
    .io_in_instrctrs_11_cycs(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_11_cycs),
    .io_in_instrctrs_11_iters(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_11_iters),
    .io_in_instrctrs_12_cycs(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_12_cycs),
    .io_in_instrctrs_12_iters(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_12_iters),
    .io_in_instrctrs_13_cycs(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_13_cycs),
    .io_in_instrctrs_13_iters(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_13_iters),
    .io_sigsIn_done(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smSelectsOut_0(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smSelectsOut_0),
    .io_sigsIn_smSelectsOut_1(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smSelectsOut_1),
    .io_sigsIn_smChildAcks_0(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_rr),
    .io_ret_number(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_ret_number)
  );
  x516_inr_UnitPipe_sm x623_inr_UnitPipe_sm ( // @[sm_x623_inr_UnitPipe.scala 34:18:@67730.4]
    .clock(x623_inr_UnitPipe_sm_clock),
    .reset(x623_inr_UnitPipe_sm_reset),
    .io_enable(x623_inr_UnitPipe_sm_io_enable),
    .io_done(x623_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x623_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x623_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x623_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x623_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x623_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x623_inr_UnitPipe_sm_io_backpressure),
    .io_break(x623_inr_UnitPipe_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_19 ( // @[package.scala 93:22:@67763.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper RetimeWrapper_20 ( // @[package.scala 93:22:@67773.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper RetimeWrapper_21 ( // @[package.scala 93:22:@67809.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper RetimeWrapper_22 ( // @[package.scala 93:22:@67817.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1 x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1 ( // @[sm_x623_inr_UnitPipe.scala 109:24:@67846.4]
    .clock(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_clock),
    .reset(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_reset),
    .io_in_x555_tmp_1_sEn_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_4),
    .io_in_x555_tmp_1_sDone_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_4),
    .io_in_x554_tmp_0_sEn_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_4),
    .io_in_x554_tmp_0_sDone_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_4),
    .io_in_x558_tmp_4_sEn_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_4),
    .io_in_x558_tmp_4_sDone_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_4),
    .io_in_x594_force_0_wPort_0_data_0(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_wPort_0_data_0),
    .io_in_x594_force_0_wPort_0_en_0(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_wPort_0_en_0),
    .io_in_x594_force_0_sEn_0(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_sEn_0),
    .io_in_x594_force_0_sDone_0(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_sDone_0),
    .io_in_x621_inr_Switch_number(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x621_inr_Switch_number),
    .io_in_x557_tmp_3_sEn_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_4),
    .io_in_x557_tmp_3_sDone_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_4),
    .io_in_x556_tmp_2_sEn_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_4),
    .io_in_x556_tmp_2_sDone_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_4),
    .io_in_instrctrs_14_cycs(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_instrctrs_14_cycs),
    .io_in_instrctrs_14_iters(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_instrctrs_14_iters),
    .io_sigsIn_done(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_done),
    .io_sigsIn_datapathEn(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_break),
    .io_rr(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_rr)
  );
  x549_ctrchain x625_ctrchain ( // @[SpatialBlocks.scala 37:22:@68366.4]
    .clock(x625_ctrchain_clock),
    .reset(x625_ctrchain_reset),
    .io_input_reset(x625_ctrchain_io_input_reset),
    .io_input_enable(x625_ctrchain_io_input_enable),
    .io_output_counts_0(x625_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x625_ctrchain_io_output_oobs_0),
    .io_output_done(x625_ctrchain_io_output_done)
  );
  x639_inr_Foreach_sm x639_inr_Foreach_sm ( // @[sm_x639_inr_Foreach.scala 33:18:@68419.4]
    .clock(x639_inr_Foreach_sm_clock),
    .reset(x639_inr_Foreach_sm_reset),
    .io_enable(x639_inr_Foreach_sm_io_enable),
    .io_done(x639_inr_Foreach_sm_io_done),
    .io_rst(x639_inr_Foreach_sm_io_rst),
    .io_ctrDone(x639_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x639_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x639_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x639_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x639_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x639_inr_Foreach_sm_io_backpressure),
    .io_break(x639_inr_Foreach_sm_io_break)
  );
  x639_inr_Foreach_iiCtr x639_inr_Foreach_iiCtr ( // @[sm_x639_inr_Foreach.scala 34:21:@68444.4]
    .clock(x639_inr_Foreach_iiCtr_clock),
    .reset(x639_inr_Foreach_iiCtr_reset),
    .io_input_enable(x639_inr_Foreach_iiCtr_io_input_enable),
    .io_input_reset(x639_inr_Foreach_iiCtr_io_input_reset),
    .io_output_issue(x639_inr_Foreach_iiCtr_io_output_issue),
    .io_output_done(x639_inr_Foreach_iiCtr_io_output_done)
  );
  RetimeWrapper RetimeWrapper_23 ( // @[package.scala 93:22:@68448.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper RetimeWrapper_24 ( // @[package.scala 93:22:@68457.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@68467.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper RetimeWrapper_26 ( // @[package.scala 93:22:@68509.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper RetimeWrapper_27 ( // @[package.scala 93:22:@68517.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1 x639_inr_Foreach_kernelx639_inr_Foreach_concrete1 ( // @[sm_x639_inr_Foreach.scala 158:24:@68551.4]
    .clock(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_clock),
    .reset(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_reset),
    .io_in_x555_tmp_1_wPort_1_ofs_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_ofs_0),
    .io_in_x555_tmp_1_wPort_1_data_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_data_0),
    .io_in_x555_tmp_1_wPort_1_en_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_en_0),
    .io_in_x555_tmp_1_sEn_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_sEn_5),
    .io_in_x555_tmp_1_sDone_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_sDone_5),
    .io_in_x554_tmp_0_wPort_1_ofs_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_ofs_0),
    .io_in_x554_tmp_0_wPort_1_data_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_data_0),
    .io_in_x554_tmp_0_wPort_1_en_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_en_0),
    .io_in_x554_tmp_0_sEn_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_sEn_5),
    .io_in_x554_tmp_0_sDone_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_sDone_5),
    .io_in_x558_tmp_4_wPort_1_ofs_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_ofs_0),
    .io_in_x558_tmp_4_wPort_1_data_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_data_0),
    .io_in_x558_tmp_4_wPort_1_en_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_en_0),
    .io_in_x558_tmp_4_sEn_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_5),
    .io_in_x558_tmp_4_sDone_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_5),
    .io_in_b552(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_b552),
    .io_in_x594_force_0_rPort_0_en_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_rPort_0_en_0),
    .io_in_x594_force_0_rPort_0_output_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_rPort_0_output_0),
    .io_in_x594_force_0_sEn_1(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_sEn_1),
    .io_in_x594_force_0_sDone_1(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_sDone_1),
    .io_in_x557_tmp_3_rPort_0_ofs_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_ofs_0),
    .io_in_x557_tmp_3_rPort_0_en_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_en_0),
    .io_in_x557_tmp_3_rPort_0_output_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_output_0),
    .io_in_x557_tmp_3_wPort_1_ofs_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_ofs_0),
    .io_in_x557_tmp_3_wPort_1_data_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_data_0),
    .io_in_x557_tmp_3_wPort_1_en_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_en_0),
    .io_in_x557_tmp_3_sEn_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_sEn_5),
    .io_in_x557_tmp_3_sDone_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_sDone_5),
    .io_in_x556_tmp_2_wPort_1_ofs_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_ofs_0),
    .io_in_x556_tmp_2_wPort_1_data_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_data_0),
    .io_in_x556_tmp_2_wPort_1_en_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_en_0),
    .io_in_x556_tmp_2_sEn_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_sEn_5),
    .io_in_x556_tmp_2_sDone_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_sDone_5),
    .io_in_b543(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_b543),
    .io_in_instrctrs_15_cycs(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_instrctrs_15_cycs),
    .io_in_instrctrs_15_iters(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_instrctrs_15_iters),
    .io_sigsIn_done(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_iiIssue(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_iiIssue),
    .io_sigsIn_datapathEn(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_rr)
  );
  x652_inr_Foreach_sm x652_inr_Foreach_sm ( // @[sm_x652_inr_Foreach.scala 35:18:@69143.4]
    .clock(x652_inr_Foreach_sm_clock),
    .reset(x652_inr_Foreach_sm_reset),
    .io_enable(x652_inr_Foreach_sm_io_enable),
    .io_done(x652_inr_Foreach_sm_io_done),
    .io_doneLatch(x652_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x652_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x652_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x652_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x652_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x652_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x652_inr_Foreach_sm_io_backpressure),
    .io_break(x652_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_28 ( // @[package.scala 93:22:@69172.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper RetimeWrapper_29 ( // @[package.scala 93:22:@69181.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper RetimeWrapper_30 ( // @[package.scala 93:22:@69191.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper RetimeWrapper_31 ( // @[package.scala 93:22:@69232.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper RetimeWrapper_32 ( // @[package.scala 93:22:@69240.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1 x652_inr_Foreach_kernelx652_inr_Foreach_concrete1 ( // @[sm_x652_inr_Foreach.scala 130:24:@69274.4]
    .clock(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_clock),
    .reset(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_reset),
    .io_in_b550_number(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_b550_number),
    .io_in_x558_tmp_4_rPort_0_ofs_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_ofs_0),
    .io_in_x558_tmp_4_rPort_0_en_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_en_0),
    .io_in_x558_tmp_4_rPort_0_output_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_output_0),
    .io_in_x558_tmp_4_sEn_6(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_6),
    .io_in_x558_tmp_4_sDone_6(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_6),
    .io_in_x545_accum_1_wPort_0_ofs_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_ofs_0),
    .io_in_x545_accum_1_wPort_0_data_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_data_0),
    .io_in_x545_accum_1_wPort_0_en_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_en_0),
    .io_in_x544_accum_0_rPort_0_ofs_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_ofs_0),
    .io_in_x544_accum_0_rPort_0_en_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_en_0),
    .io_in_x544_accum_0_rPort_0_output_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_output_0),
    .io_in_x544_accum_0_wPort_0_ofs_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_ofs_0),
    .io_in_x544_accum_0_wPort_0_data_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_data_0),
    .io_in_x544_accum_0_wPort_0_en_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_en_0),
    .io_in_b543(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_b543),
    .io_in_instrctrs_16_cycs(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_instrctrs_16_cycs),
    .io_in_instrctrs_16_iters(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_instrctrs_16_iters),
    .io_sigsIn_done(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_datapathEn(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_rr)
  );
  RetimeWrapper RetimeWrapper_33 ( // @[package.scala 93:22:@69577.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  assign _T_786 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@64030.4]
  assign b552 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x653_outr_Reduce.scala 100:18:@64190.4]
  assign b552_chain_read_1 = b552_chain_io_rPort_0_output_0; // @[sm_x653_outr_Reduce.scala 103:61:@64264.4]
  assign b552_chain_read_2 = b552_chain_io_rPort_1_output_0; // @[sm_x653_outr_Reduce.scala 104:61:@64265.4]
  assign b552_chain_read_4 = b552_chain_io_rPort_3_output_0; // @[sm_x653_outr_Reduce.scala 106:61:@64267.4]
  assign b552_chain_read_5 = b552_chain_io_rPort_4_output_0; // @[sm_x653_outr_Reduce.scala 107:61:@64268.4]
  assign _T_911 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@64594.4 package.scala 96:25:@64595.4]
  assign _T_915 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@64603.4 package.scala 96:25:@64604.4]
  assign _T_919 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@64613.4 package.scala 96:25:@64614.4]
  assign x579_inr_Foreach_mySignalsIn_mask = b552 & io_in_b543; // @[sm_x653_outr_Reduce.scala 126:81:@64627.4]
  assign _T_936 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@64655.4 package.scala 96:25:@64656.4]
  assign _T_942 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@64663.4 package.scala 96:25:@64664.4]
  assign _T_945 = ~ _T_942; // @[SpatialBlocks.scala 137:99:@64666.4]
  assign _T_947 = x579_inr_Foreach_sm_io_datapathEn & x579_inr_Foreach_mySignalsIn_mask; // @[SpatialBlocks.scala 156:36:@64675.4]
  assign _T_948 = ~ x579_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 156:78:@64676.4]
  assign _T_1016 = x593_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@65339.4]
  assign _T_1022 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@65349.4 package.scala 96:25:@65350.4]
  assign _T_1026 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@65359.4 package.scala 96:25:@65360.4]
  assign x593_inr_UnitPipe_mySignalsIn_mask = b552_chain_read_1 & io_in_b543; // @[sm_x653_outr_Reduce.scala 138:60:@65372.4]
  assign _T_1043 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@65395.4 package.scala 96:25:@65396.4]
  assign _T_1049 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@65403.4 package.scala 96:25:@65404.4]
  assign _T_1052 = ~ _T_1049; // @[SpatialBlocks.scala 137:99:@65406.4]
  assign _T_1123 = x605_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@66132.4]
  assign _T_1129 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@66142.4 package.scala 96:25:@66143.4]
  assign _T_1133 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@66152.4 package.scala 96:25:@66153.4]
  assign x605_inr_UnitPipe_mySignalsIn_mask = b552_chain_read_2 & io_in_b543; // @[sm_x653_outr_Reduce.scala 152:60:@66165.4]
  assign _T_1150 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@66188.4 package.scala 96:25:@66189.4]
  assign _T_1156 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@66196.4 package.scala 96:25:@66197.4]
  assign _T_1159 = ~ _T_1156; // @[SpatialBlocks.scala 137:99:@66199.4]
  assign _T_1257 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@66965.4 package.scala 96:25:@66966.4]
  assign _T_1261 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@66975.4 package.scala 96:25:@66976.4]
  assign _T_1279 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@67017.4 package.scala 96:25:@67018.4]
  assign _T_1285 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@67025.4 package.scala 96:25:@67026.4]
  assign _T_1288 = ~ _T_1285; // @[SpatialBlocks.scala 137:99:@67028.4]
  assign _T_1356 = x623_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@67758.4]
  assign _T_1362 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@67768.4 package.scala 96:25:@67769.4]
  assign _T_1366 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@67778.4 package.scala 96:25:@67779.4]
  assign x623_inr_UnitPipe_mySignalsIn_mask = b552_chain_read_4 & io_in_b543; // @[sm_x653_outr_Reduce.scala 188:60:@67791.4]
  assign _T_1383 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@67814.4 package.scala 96:25:@67815.4]
  assign _T_1389 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@67822.4 package.scala 96:25:@67823.4]
  assign _T_1392 = ~ _T_1389; // @[SpatialBlocks.scala 137:99:@67825.4]
  assign _T_1464 = RetimeWrapper_23_io_out; // @[package.scala 96:25:@68453.4 package.scala 96:25:@68454.4]
  assign _T_1468 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@68462.4 package.scala 96:25:@68463.4]
  assign _T_1472 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@68472.4 package.scala 96:25:@68473.4]
  assign x639_inr_Foreach_mySignalsIn_mask = b552_chain_read_5 & io_in_b543; // @[sm_x653_outr_Reduce.scala 203:94:@68486.4]
  assign _T_1489 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@68514.4 package.scala 96:25:@68515.4]
  assign _T_1495 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@68522.4 package.scala 96:25:@68523.4]
  assign _T_1498 = ~ _T_1495; // @[SpatialBlocks.scala 137:99:@68525.4]
  assign _T_1500 = x639_inr_Foreach_sm_io_datapathEn & x639_inr_Foreach_mySignalsIn_mask; // @[SpatialBlocks.scala 156:36:@68534.4]
  assign _T_1501 = ~ x639_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 156:78:@68535.4]
  assign _T_1504 = ~ x639_inr_Foreach_mySignalsIn_mask; // @[SpatialBlocks.scala 157:128:@68541.4]
  assign x639_inr_Foreach_mySignalsIn_iiDone = x639_inr_Foreach_iiCtr_io_output_done | _T_1504; // @[SpatialBlocks.scala 157:126:@68542.4]
  assign _T_1570 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@69177.4 package.scala 96:25:@69178.4]
  assign _T_1574 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@69186.4 package.scala 96:25:@69187.4]
  assign _T_1578 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@69196.4 package.scala 96:25:@69197.4]
  assign _T_1595 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@69237.4 package.scala 96:25:@69238.4]
  assign _T_1601 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@69245.4 package.scala 96:25:@69246.4]
  assign _T_1604 = ~ _T_1601; // @[SpatialBlocks.scala 137:99:@69248.4]
  assign _T_1606 = x652_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 156:36:@69257.4]
  assign _T_1607 = ~ x652_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 156:78:@69258.4]
  assign _T_1619 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@69582.4 package.scala 96:25:@69583.4]
  assign io_in_x472_A_sram_1_rPort_0_ofs_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@65095.4]
  assign io_in_x472_A_sram_1_rPort_0_en_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@65094.4]
  assign io_in_x471_A_sram_0_rPort_0_ofs_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@65101.4]
  assign io_in_x471_A_sram_0_rPort_0_en_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@65100.4]
  assign io_in_x545_accum_1_wPort_0_ofs_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@69530.4]
  assign io_in_x545_accum_1_wPort_0_data_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@69529.4]
  assign io_in_x545_accum_1_wPort_0_en_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@69525.4]
  assign io_in_x545_accum_1_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@69585.4]
  assign io_in_x545_accum_1_sDone_0 = io_rr ? _T_1619 : 1'h0; // @[MemInterfaceType.scala 197:17:@69586.4]
  assign io_in_x544_accum_0_rPort_0_ofs_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@69535.4]
  assign io_in_x544_accum_0_rPort_0_en_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@69534.4]
  assign io_in_x544_accum_0_wPort_0_ofs_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@69542.4]
  assign io_in_x544_accum_0_wPort_0_data_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@69541.4]
  assign io_in_x544_accum_0_wPort_0_en_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@69537.4]
  assign io_in_x549_ctrchain_input_reset = x652_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@69273.4]
  assign io_in_x549_ctrchain_input_enable = x652_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 158:42:@69272.4]
  assign io_in_instrctrs_7_cycs = cycles_x653_outr_Reduce_io_count; // @[Ledger.scala 293:21:@64035.4]
  assign io_in_instrctrs_7_iters = iters_x653_outr_Reduce_io_count; // @[Ledger.scala 294:22:@64036.4]
  assign io_in_instrctrs_8_cycs = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_instrctrs_8_cycs; // @[Ledger.scala 302:78:@65208.4]
  assign io_in_instrctrs_8_iters = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_instrctrs_8_iters; // @[Ledger.scala 302:78:@65207.4]
  assign io_in_instrctrs_9_cycs = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_instrctrs_9_cycs; // @[Ledger.scala 302:78:@65943.4]
  assign io_in_instrctrs_9_iters = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_instrctrs_9_iters; // @[Ledger.scala 302:78:@65942.4]
  assign io_in_instrctrs_10_cycs = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_instrctrs_10_cycs; // @[Ledger.scala 302:78:@66826.4]
  assign io_in_instrctrs_10_iters = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_instrctrs_10_iters; // @[Ledger.scala 302:78:@66825.4]
  assign io_in_instrctrs_11_cycs = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_11_cycs; // @[Ledger.scala 302:78:@67652.4]
  assign io_in_instrctrs_11_iters = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_11_iters; // @[Ledger.scala 302:78:@67651.4]
  assign io_in_instrctrs_12_cycs = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_12_cycs; // @[Ledger.scala 302:78:@67656.4]
  assign io_in_instrctrs_12_iters = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_12_iters; // @[Ledger.scala 302:78:@67655.4]
  assign io_in_instrctrs_13_cycs = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_13_cycs; // @[Ledger.scala 302:78:@67660.4]
  assign io_in_instrctrs_13_iters = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_instrctrs_13_iters; // @[Ledger.scala 302:78:@67659.4]
  assign io_in_instrctrs_14_cycs = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_instrctrs_14_cycs; // @[Ledger.scala 302:78:@68338.4]
  assign io_in_instrctrs_14_iters = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_instrctrs_14_iters; // @[Ledger.scala 302:78:@68337.4]
  assign io_in_instrctrs_15_cycs = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_instrctrs_15_cycs; // @[Ledger.scala 302:78:@69079.4]
  assign io_in_instrctrs_15_iters = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_instrctrs_15_iters; // @[Ledger.scala 302:78:@69078.4]
  assign io_in_instrctrs_16_cycs = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_instrctrs_16_cycs; // @[Ledger.scala 302:78:@69548.4]
  assign io_in_instrctrs_16_iters = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_instrctrs_16_iters; // @[Ledger.scala 302:78:@69547.4]
  assign io_sigsOut_smDoneIn_0 = x579_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@64673.4]
  assign io_sigsOut_smDoneIn_1 = x593_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 155:56:@65413.4]
  assign io_sigsOut_smDoneIn_2 = x605_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 155:56:@66206.4]
  assign io_sigsOut_smDoneIn_3 = x621_inr_Switch_sm_io_done; // @[SpatialBlocks.scala 155:56:@67035.4]
  assign io_sigsOut_smDoneIn_4 = x623_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 155:56:@67832.4]
  assign io_sigsOut_smDoneIn_5 = x639_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@68532.4]
  assign io_sigsOut_smDoneIn_6 = x652_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@69255.4]
  assign io_sigsOut_smMaskIn_0 = b552 & io_in_b543; // @[SpatialBlocks.scala 155:86:@64674.4]
  assign io_sigsOut_smMaskIn_1 = b552_chain_read_1 & io_in_b543; // @[SpatialBlocks.scala 155:86:@65414.4]
  assign io_sigsOut_smMaskIn_2 = b552_chain_read_2 & io_in_b543; // @[SpatialBlocks.scala 155:86:@66207.4]
  assign io_sigsOut_smMaskIn_4 = b552_chain_read_4 & io_in_b543; // @[SpatialBlocks.scala 155:86:@67833.4]
  assign io_sigsOut_smMaskIn_5 = b552_chain_read_5 & io_in_b543; // @[SpatialBlocks.scala 155:86:@68533.4]
  assign cycles_x653_outr_Reduce_clock = clock; // @[:@64024.4]
  assign cycles_x653_outr_Reduce_reset = reset; // @[:@64025.4]
  assign cycles_x653_outr_Reduce_io_enable = io_sigsIn_baseEn; // @[sm_x653_outr_Reduce.scala 88:41:@64029.4]
  assign iters_x653_outr_Reduce_clock = clock; // @[:@64027.4]
  assign iters_x653_outr_Reduce_reset = reset; // @[:@64028.4]
  assign iters_x653_outr_Reduce_io_enable = io_sigsIn_done & _T_789; // @[sm_x653_outr_Reduce.scala 89:40:@64034.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@64046.4]
  assign b550_chain_clock = clock; // @[:@64052.4]
  assign b550_chain_reset = reset; // @[:@64053.4]
  assign b550_chain_io_wPort_0_data_0 = __io_result; // @[NBuffers.scala 309:54:@64113.4]
  assign b550_chain_io_wPort_0_reset = RetimeWrapper_io_out; // @[NBuffers.scala 312:23:@64122.4]
  assign b550_chain_io_wPort_0_en_0 = io_sigsOut_smDoneIn_0; // @[NBuffers.scala 311:25:@64114.4]
  assign b550_chain_io_sEn_0 = _T_936 & _T_945; // @[NBuffers.scala 302:18:@64606.4]
  assign b550_chain_io_sEn_1 = _T_1043 & _T_1052; // @[NBuffers.scala 302:18:@65352.4]
  assign b550_chain_io_sEn_2 = _T_1150 & _T_1159; // @[NBuffers.scala 302:18:@66145.4]
  assign b550_chain_io_sEn_3 = _T_1279 & _T_1288; // @[NBuffers.scala 302:18:@66968.4]
  assign b550_chain_io_sEn_4 = _T_1383 & _T_1392; // @[NBuffers.scala 302:18:@67771.4]
  assign b550_chain_io_sEn_5 = _T_1489 & _T_1498; // @[NBuffers.scala 302:18:@68465.4]
  assign b550_chain_io_sEn_6 = _T_1595 & _T_1604; // @[NBuffers.scala 302:18:@69189.4]
  assign b550_chain_io_sDone_0 = io_rr ? _T_915 : 1'h0; // @[NBuffers.scala 303:20:@64607.4]
  assign b550_chain_io_sDone_1 = io_rr ? _T_1022 : 1'h0; // @[NBuffers.scala 303:20:@65353.4]
  assign b550_chain_io_sDone_2 = io_rr ? _T_1129 : 1'h0; // @[NBuffers.scala 303:20:@66146.4]
  assign b550_chain_io_sDone_3 = io_rr ? _T_1257 : 1'h0; // @[NBuffers.scala 303:20:@66969.4]
  assign b550_chain_io_sDone_4 = io_rr ? _T_1362 : 1'h0; // @[NBuffers.scala 303:20:@67772.4]
  assign b550_chain_io_sDone_5 = io_rr ? _T_1468 : 1'h0; // @[NBuffers.scala 303:20:@68466.4]
  assign b550_chain_io_sDone_6 = io_rr ? _T_1574 : 1'h0; // @[NBuffers.scala 303:20:@69190.4]
  assign RetimeWrapper_clock = clock; // @[:@64116.4]
  assign RetimeWrapper_reset = reset; // @[:@64117.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@64119.4]
  assign RetimeWrapper_io_in = b550_chain_reset; // @[package.scala 94:16:@64118.4]
  assign __1_io_b = b550_chain_io_rPort_0_output_0; // @[Math.scala 721:17:@64130.4]
  assign __2_io_b = b550_chain_io_rPort_1_output_0; // @[Math.scala 721:17:@64141.4]
  assign __3_io_b = b550_chain_io_rPort_2_output_0; // @[Math.scala 721:17:@64152.4]
  assign __4_io_b = b550_chain_io_rPort_3_output_0; // @[Math.scala 721:17:@64163.4]
  assign __5_io_b = b550_chain_io_rPort_4_output_0; // @[Math.scala 721:17:@64174.4]
  assign __6_io_b = b550_chain_io_rPort_5_output_0; // @[Math.scala 721:17:@64185.4]
  assign b552_chain_clock = clock; // @[:@64192.4]
  assign b552_chain_reset = reset; // @[:@64193.4]
  assign b552_chain_io_wPort_0_data_0 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[NBuffers.scala 308:54:@64253.4]
  assign b552_chain_io_wPort_0_reset = RetimeWrapper_1_io_out; // @[NBuffers.scala 312:23:@64262.4]
  assign b552_chain_io_wPort_0_en_0 = io_sigsOut_smDoneIn_0; // @[NBuffers.scala 311:25:@64254.4]
  assign b552_chain_io_sEn_0 = _T_936 & _T_945; // @[NBuffers.scala 302:18:@64616.4]
  assign b552_chain_io_sEn_1 = _T_1043 & _T_1052; // @[NBuffers.scala 302:18:@65362.4]
  assign b552_chain_io_sEn_2 = _T_1150 & _T_1159; // @[NBuffers.scala 302:18:@66155.4]
  assign b552_chain_io_sEn_3 = _T_1279 & _T_1288; // @[NBuffers.scala 302:18:@66978.4]
  assign b552_chain_io_sEn_4 = _T_1383 & _T_1392; // @[NBuffers.scala 302:18:@67781.4]
  assign b552_chain_io_sEn_5 = _T_1489 & _T_1498; // @[NBuffers.scala 302:18:@68475.4]
  assign b552_chain_io_sEn_6 = _T_1595 & _T_1604; // @[NBuffers.scala 302:18:@69199.4]
  assign b552_chain_io_sDone_0 = io_rr ? _T_919 : 1'h0; // @[NBuffers.scala 303:20:@64617.4]
  assign b552_chain_io_sDone_1 = io_rr ? _T_1026 : 1'h0; // @[NBuffers.scala 303:20:@65363.4]
  assign b552_chain_io_sDone_2 = io_rr ? _T_1133 : 1'h0; // @[NBuffers.scala 303:20:@66156.4]
  assign b552_chain_io_sDone_3 = io_rr ? _T_1261 : 1'h0; // @[NBuffers.scala 303:20:@66979.4]
  assign b552_chain_io_sDone_4 = io_rr ? _T_1366 : 1'h0; // @[NBuffers.scala 303:20:@67782.4]
  assign b552_chain_io_sDone_5 = io_rr ? _T_1472 : 1'h0; // @[NBuffers.scala 303:20:@68476.4]
  assign b552_chain_io_sDone_6 = io_rr ? _T_1578 : 1'h0; // @[NBuffers.scala 303:20:@69200.4]
  assign RetimeWrapper_1_clock = clock; // @[:@64256.4]
  assign RetimeWrapper_1_reset = reset; // @[:@64257.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@64259.4]
  assign RetimeWrapper_1_io_in = b552_chain_reset; // @[package.scala 94:16:@64258.4]
  assign x554_tmp_0_clock = clock; // @[:@64271.4]
  assign x554_tmp_0_reset = reset; // @[:@64272.4]
  assign x554_tmp_0_io_rPort_0_ofs_0 = 2'h0; // @[MemInterfaceType.scala 66:44:@65852.4]
  assign x554_tmp_0_io_rPort_0_en_0 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@65851.4]
  assign x554_tmp_0_io_wPort_1_ofs_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_ofs_0; // @[MemInterfaceType.scala 67:44:@68971.4]
  assign x554_tmp_0_io_wPort_1_data_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_data_0; // @[MemInterfaceType.scala 67:44:@68970.4]
  assign x554_tmp_0_io_wPort_1_en_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_en_0; // @[MemInterfaceType.scala 67:44:@68966.4]
  assign x554_tmp_0_io_wPort_0_ofs_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@65126.4]
  assign x554_tmp_0_io_wPort_0_data_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@65125.4]
  assign x554_tmp_0_io_wPort_0_en_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@65121.4]
  assign x554_tmp_0_io_sEn_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_sEn_0; // @[MemInterfaceType.scala 189:41:@65111.4]
  assign x554_tmp_0_io_sEn_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_1; // @[MemInterfaceType.scala 189:41:@65839.4]
  assign x554_tmp_0_io_sEn_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_2; // @[MemInterfaceType.scala 189:41:@66686.4]
  assign x554_tmp_0_io_sEn_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x554_tmp_0_sEn_3; // @[MemInterfaceType.scala 189:41:@67521.4]
  assign x554_tmp_0_io_sEn_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_4; // @[MemInterfaceType.scala 189:41:@68245.4]
  assign x554_tmp_0_io_sEn_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_sEn_5; // @[MemInterfaceType.scala 189:41:@68956.4]
  assign x554_tmp_0_io_sDone_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_sDone_0; // @[MemInterfaceType.scala 189:64:@65112.4]
  assign x554_tmp_0_io_sDone_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_1; // @[MemInterfaceType.scala 189:64:@65840.4]
  assign x554_tmp_0_io_sDone_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_2; // @[MemInterfaceType.scala 189:64:@66687.4]
  assign x554_tmp_0_io_sDone_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x554_tmp_0_sDone_3; // @[MemInterfaceType.scala 189:64:@67522.4]
  assign x554_tmp_0_io_sDone_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_4; // @[MemInterfaceType.scala 189:64:@68246.4]
  assign x554_tmp_0_io_sDone_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_sDone_5; // @[MemInterfaceType.scala 189:64:@68957.4]
  assign x555_tmp_1_clock = clock; // @[:@64318.4]
  assign x555_tmp_1_reset = reset; // @[:@64319.4]
  assign x555_tmp_1_io_rPort_0_ofs_0 = 2'h1; // @[MemInterfaceType.scala 66:44:@65829.4]
  assign x555_tmp_1_io_rPort_0_en_0 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@65828.4]
  assign x555_tmp_1_io_wPort_1_ofs_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_ofs_0; // @[MemInterfaceType.scala 67:44:@68946.4]
  assign x555_tmp_1_io_wPort_1_data_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_data_0; // @[MemInterfaceType.scala 67:44:@68945.4]
  assign x555_tmp_1_io_wPort_1_en_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_en_0; // @[MemInterfaceType.scala 67:44:@68941.4]
  assign x555_tmp_1_io_wPort_0_ofs_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@65089.4]
  assign x555_tmp_1_io_wPort_0_data_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@65088.4]
  assign x555_tmp_1_io_wPort_0_en_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@65084.4]
  assign x555_tmp_1_io_sEn_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_sEn_0; // @[MemInterfaceType.scala 189:41:@65074.4]
  assign x555_tmp_1_io_sEn_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_1; // @[MemInterfaceType.scala 189:41:@65816.4]
  assign x555_tmp_1_io_sEn_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_2; // @[MemInterfaceType.scala 189:41:@66668.4]
  assign x555_tmp_1_io_sEn_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x555_tmp_1_sEn_3; // @[MemInterfaceType.scala 189:41:@67503.4]
  assign x555_tmp_1_io_sEn_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_4; // @[MemInterfaceType.scala 189:41:@68227.4]
  assign x555_tmp_1_io_sEn_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_sEn_5; // @[MemInterfaceType.scala 189:41:@68931.4]
  assign x555_tmp_1_io_sDone_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_sDone_0; // @[MemInterfaceType.scala 189:64:@65075.4]
  assign x555_tmp_1_io_sDone_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_1; // @[MemInterfaceType.scala 189:64:@65817.4]
  assign x555_tmp_1_io_sDone_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_2; // @[MemInterfaceType.scala 189:64:@66669.4]
  assign x555_tmp_1_io_sDone_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x555_tmp_1_sDone_3; // @[MemInterfaceType.scala 189:64:@67504.4]
  assign x555_tmp_1_io_sDone_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_4; // @[MemInterfaceType.scala 189:64:@68228.4]
  assign x555_tmp_1_io_sDone_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_sDone_5; // @[MemInterfaceType.scala 189:64:@68932.4]
  assign x556_tmp_2_clock = clock; // @[:@64365.4]
  assign x556_tmp_2_reset = reset; // @[:@64366.4]
  assign x556_tmp_2_io_rPort_0_ofs_0 = 2'h2; // @[MemInterfaceType.scala 66:44:@65937.4]
  assign x556_tmp_2_io_rPort_0_en_0 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@65936.4]
  assign x556_tmp_2_io_wPort_1_ofs_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_ofs_0; // @[MemInterfaceType.scala 67:44:@69073.4]
  assign x556_tmp_2_io_wPort_1_data_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_data_0; // @[MemInterfaceType.scala 67:44:@69072.4]
  assign x556_tmp_2_io_wPort_1_en_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_en_0; // @[MemInterfaceType.scala 67:44:@69068.4]
  assign x556_tmp_2_io_wPort_0_ofs_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@65202.4]
  assign x556_tmp_2_io_wPort_0_data_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@65201.4]
  assign x556_tmp_2_io_wPort_0_en_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@65197.4]
  assign x556_tmp_2_io_sEn_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_sEn_0; // @[MemInterfaceType.scala 189:41:@65187.4]
  assign x556_tmp_2_io_sEn_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_1; // @[MemInterfaceType.scala 189:41:@65924.4]
  assign x556_tmp_2_io_sEn_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_2; // @[MemInterfaceType.scala 189:41:@66789.4]
  assign x556_tmp_2_io_sEn_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x556_tmp_2_sEn_3; // @[MemInterfaceType.scala 189:41:@67622.4]
  assign x556_tmp_2_io_sEn_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_4; // @[MemInterfaceType.scala 189:41:@68324.4]
  assign x556_tmp_2_io_sEn_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_sEn_5; // @[MemInterfaceType.scala 189:41:@69058.4]
  assign x556_tmp_2_io_sDone_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_sDone_0; // @[MemInterfaceType.scala 189:64:@65188.4]
  assign x556_tmp_2_io_sDone_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_1; // @[MemInterfaceType.scala 189:64:@65925.4]
  assign x556_tmp_2_io_sDone_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_2; // @[MemInterfaceType.scala 189:64:@66790.4]
  assign x556_tmp_2_io_sDone_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x556_tmp_2_sDone_3; // @[MemInterfaceType.scala 189:64:@67623.4]
  assign x556_tmp_2_io_sDone_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_4; // @[MemInterfaceType.scala 189:64:@68325.4]
  assign x556_tmp_2_io_sDone_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_sDone_5; // @[MemInterfaceType.scala 189:64:@69059.4]
  assign x557_tmp_3_clock = clock; // @[:@64412.4]
  assign x557_tmp_3_reset = reset; // @[:@64413.4]
  assign x557_tmp_3_io_rPort_0_ofs_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@69041.4]
  assign x557_tmp_3_io_rPort_0_en_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@69040.4]
  assign x557_tmp_3_io_wPort_1_ofs_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_ofs_0; // @[MemInterfaceType.scala 67:44:@69048.4]
  assign x557_tmp_3_io_wPort_1_data_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_data_0; // @[MemInterfaceType.scala 67:44:@69047.4]
  assign x557_tmp_3_io_wPort_1_en_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_en_0; // @[MemInterfaceType.scala 67:44:@69043.4]
  assign x557_tmp_3_io_wPort_0_ofs_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@65177.4]
  assign x557_tmp_3_io_wPort_0_data_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@65176.4]
  assign x557_tmp_3_io_wPort_0_en_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@65172.4]
  assign x557_tmp_3_io_sEn_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_sEn_0; // @[MemInterfaceType.scala 189:41:@65162.4]
  assign x557_tmp_3_io_sEn_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_1; // @[MemInterfaceType.scala 189:41:@65881.4]
  assign x557_tmp_3_io_sEn_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_2; // @[MemInterfaceType.scala 189:41:@66723.4]
  assign x557_tmp_3_io_sEn_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x557_tmp_3_sEn_3; // @[MemInterfaceType.scala 189:41:@67558.4]
  assign x557_tmp_3_io_sEn_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_4; // @[MemInterfaceType.scala 189:41:@68306.4]
  assign x557_tmp_3_io_sEn_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_sEn_5; // @[MemInterfaceType.scala 189:41:@69028.4]
  assign x557_tmp_3_io_sDone_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_sDone_0; // @[MemInterfaceType.scala 189:64:@65163.4]
  assign x557_tmp_3_io_sDone_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_1; // @[MemInterfaceType.scala 189:64:@65882.4]
  assign x557_tmp_3_io_sDone_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_2; // @[MemInterfaceType.scala 189:64:@66724.4]
  assign x557_tmp_3_io_sDone_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x557_tmp_3_sDone_3; // @[MemInterfaceType.scala 189:64:@67559.4]
  assign x557_tmp_3_io_sDone_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_4; // @[MemInterfaceType.scala 189:64:@68307.4]
  assign x557_tmp_3_io_sDone_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_sDone_5; // @[MemInterfaceType.scala 189:64:@69029.4]
  assign x558_tmp_4_clock = clock; // @[:@64459.4]
  assign x558_tmp_4_reset = reset; // @[:@64460.4]
  assign x558_tmp_4_io_rPort_0_ofs_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@69509.4]
  assign x558_tmp_4_io_rPort_0_en_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@69508.4]
  assign x558_tmp_4_io_wPort_1_ofs_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_ofs_0; // @[MemInterfaceType.scala 67:44:@68996.4]
  assign x558_tmp_4_io_wPort_1_data_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_data_0; // @[MemInterfaceType.scala 67:44:@68995.4]
  assign x558_tmp_4_io_wPort_1_en_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_en_0; // @[MemInterfaceType.scala 67:44:@68991.4]
  assign x558_tmp_4_io_wPort_0_ofs_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@65151.4]
  assign x558_tmp_4_io_wPort_0_data_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@65150.4]
  assign x558_tmp_4_io_wPort_0_en_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@65146.4]
  assign x558_tmp_4_io_sEn_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_0; // @[MemInterfaceType.scala 189:41:@65136.4]
  assign x558_tmp_4_io_sEn_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_1; // @[MemInterfaceType.scala 189:41:@65862.4]
  assign x558_tmp_4_io_sEn_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_2; // @[MemInterfaceType.scala 189:41:@66704.4]
  assign x558_tmp_4_io_sEn_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x558_tmp_4_sEn_3; // @[MemInterfaceType.scala 189:41:@67539.4]
  assign x558_tmp_4_io_sEn_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_4; // @[MemInterfaceType.scala 189:41:@68263.4]
  assign x558_tmp_4_io_sEn_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_5; // @[MemInterfaceType.scala 189:41:@68981.4]
  assign x558_tmp_4_io_sEn_6 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_6; // @[MemInterfaceType.scala 189:41:@69496.4]
  assign x558_tmp_4_io_sDone_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_0; // @[MemInterfaceType.scala 189:64:@65137.4]
  assign x558_tmp_4_io_sDone_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_1; // @[MemInterfaceType.scala 189:64:@65863.4]
  assign x558_tmp_4_io_sDone_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_2; // @[MemInterfaceType.scala 189:64:@66705.4]
  assign x558_tmp_4_io_sDone_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x558_tmp_4_sDone_3; // @[MemInterfaceType.scala 189:64:@67540.4]
  assign x558_tmp_4_io_sDone_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_4; // @[MemInterfaceType.scala 189:64:@68264.4]
  assign x558_tmp_4_io_sDone_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_5; // @[MemInterfaceType.scala 189:64:@68982.4]
  assign x558_tmp_4_io_sDone_6 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_6; // @[MemInterfaceType.scala 189:64:@69497.4]
  assign x560_ctrchain_clock = clock; // @[:@64508.4]
  assign x560_ctrchain_reset = reset; // @[:@64509.4]
  assign x560_ctrchain_io_input_reset = x579_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@64691.4]
  assign x560_ctrchain_io_input_enable = x579_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 158:42:@64690.4]
  assign x579_inr_Foreach_sm_clock = clock; // @[:@64561.4]
  assign x579_inr_Foreach_sm_reset = reset; // @[:@64562.4]
  assign x579_inr_Foreach_sm_io_enable = _T_936 & _T_945; // @[SpatialBlocks.scala 139:18:@64670.4]
  assign x579_inr_Foreach_sm_io_ctrDone = io_rr ? _T_911 : 1'h0; // @[sm_x653_outr_Reduce.scala 119:38:@64597.4]
  assign x579_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@64672.4]
  assign x579_inr_Foreach_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@64644.4]
  assign x579_inr_Foreach_sm_io_break = 1'h0; // @[sm_x653_outr_Reduce.scala 125:36:@64624.4]
  assign RetimeWrapper_2_clock = clock; // @[:@64590.4]
  assign RetimeWrapper_2_reset = reset; // @[:@64591.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@64593.4]
  assign RetimeWrapper_2_io_in = x560_ctrchain_io_output_done; // @[package.scala 94:16:@64592.4]
  assign RetimeWrapper_3_clock = clock; // @[:@64599.4]
  assign RetimeWrapper_3_reset = reset; // @[:@64600.4]
  assign RetimeWrapper_3_io_flow = x579_inr_Foreach_sm_io_backpressure; // @[package.scala 95:18:@64602.4]
  assign RetimeWrapper_3_io_in = x579_inr_Foreach_sm_io_done; // @[package.scala 94:16:@64601.4]
  assign RetimeWrapper_4_clock = clock; // @[:@64609.4]
  assign RetimeWrapper_4_reset = reset; // @[:@64610.4]
  assign RetimeWrapper_4_io_flow = x579_inr_Foreach_sm_io_backpressure; // @[package.scala 95:18:@64612.4]
  assign RetimeWrapper_4_io_in = x579_inr_Foreach_sm_io_done; // @[package.scala 94:16:@64611.4]
  assign RetimeWrapper_5_clock = clock; // @[:@64651.4]
  assign RetimeWrapper_5_reset = reset; // @[:@64652.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@64654.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@64653.4]
  assign RetimeWrapper_6_clock = clock; // @[:@64659.4]
  assign RetimeWrapper_6_reset = reset; // @[:@64660.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@64662.4]
  assign RetimeWrapper_6_io_in = x579_inr_Foreach_sm_io_done; // @[package.scala 94:16:@64661.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_clock = clock; // @[:@64693.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_reset = reset; // @[:@64694.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b550_number = __io_result; // @[sm_x579_inr_Foreach.scala 71:23:@65091.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_output_0 = io_in_x472_A_sram_1_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@65092.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b542_number = io_in_b542_number; // @[sm_x579_inr_Foreach.scala 73:23:@65097.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_output_0 = io_in_x471_A_sram_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@65098.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b552 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x579_inr_Foreach.scala 77:23:@65153.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b543 = io_in_b543; // @[sm_x579_inr_Foreach.scala 80:23:@65204.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_done = x579_inr_Foreach_sm_io_done; // @[sm_x579_inr_Foreach.scala 193:22:@65228.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_947 & _T_948; // @[sm_x579_inr_Foreach.scala 193:22:@65221.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_baseEn = _T_936 & _T_945; // @[sm_x579_inr_Foreach.scala 193:22:@65220.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_break = x579_inr_Foreach_sm_io_break; // @[sm_x579_inr_Foreach.scala 193:22:@65219.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{28{x560_ctrchain_io_output_counts_0[3]}},x560_ctrchain_io_output_counts_0}; // @[sm_x579_inr_Foreach.scala 193:22:@65214.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x560_ctrchain_io_output_oobs_0; // @[sm_x579_inr_Foreach.scala 193:22:@65213.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x579_inr_Foreach.scala 192:18:@65209.4]
  assign x580_r_0_clock = clock; // @[:@65237.4]
  assign x580_r_0_reset = reset; // @[:@65238.4]
  assign x580_r_0_io_rPort_1_en_0 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_rPort_1_en_0; // @[MemInterfaceType.scala 66:44:@67588.4]
  assign x580_r_0_io_rPort_0_en_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@66753.4]
  assign x580_r_0_io_wPort_0_data_0 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@65913.4]
  assign x580_r_0_io_wPort_0_en_0 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@65909.4]
  assign x580_r_0_io_sEn_0 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_sEn_0; // @[MemInterfaceType.scala 189:41:@65899.4]
  assign x580_r_0_io_sEn_1 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_sEn_1; // @[MemInterfaceType.scala 189:41:@66741.4]
  assign x580_r_0_io_sEn_2 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_sEn_2; // @[MemInterfaceType.scala 189:41:@67576.4]
  assign x580_r_0_io_sDone_0 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_sDone_0; // @[MemInterfaceType.scala 189:64:@65900.4]
  assign x580_r_0_io_sDone_1 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_sDone_1; // @[MemInterfaceType.scala 189:64:@66742.4]
  assign x580_r_0_io_sDone_2 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_sDone_2; // @[MemInterfaceType.scala 189:64:@67577.4]
  assign x593_inr_UnitPipe_sm_clock = clock; // @[:@65312.4]
  assign x593_inr_UnitPipe_sm_reset = reset; // @[:@65313.4]
  assign x593_inr_UnitPipe_sm_io_enable = _T_1043 & _T_1052; // @[SpatialBlocks.scala 139:18:@65410.4]
  assign x593_inr_UnitPipe_sm_io_ctrDone = x593_inr_UnitPipe_sm_io_ctrInc & _T_1019; // @[sm_x653_outr_Reduce.scala 131:39:@65343.4]
  assign x593_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 141:21:@65412.4]
  assign x593_inr_UnitPipe_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@65384.4]
  assign x593_inr_UnitPipe_sm_io_break = 1'h0; // @[sm_x653_outr_Reduce.scala 137:37:@65370.4]
  assign RetimeWrapper_7_clock = clock; // @[:@65345.4]
  assign RetimeWrapper_7_reset = reset; // @[:@65346.4]
  assign RetimeWrapper_7_io_flow = x593_inr_UnitPipe_sm_io_backpressure; // @[package.scala 95:18:@65348.4]
  assign RetimeWrapper_7_io_in = x593_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@65347.4]
  assign RetimeWrapper_8_clock = clock; // @[:@65355.4]
  assign RetimeWrapper_8_reset = reset; // @[:@65356.4]
  assign RetimeWrapper_8_io_flow = x593_inr_UnitPipe_sm_io_backpressure; // @[package.scala 95:18:@65358.4]
  assign RetimeWrapper_8_io_in = x593_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@65357.4]
  assign RetimeWrapper_9_clock = clock; // @[:@65391.4]
  assign RetimeWrapper_9_reset = reset; // @[:@65392.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@65394.4]
  assign RetimeWrapper_9_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@65393.4]
  assign RetimeWrapper_10_clock = clock; // @[:@65399.4]
  assign RetimeWrapper_10_reset = reset; // @[:@65400.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@65402.4]
  assign RetimeWrapper_10_io_in = x593_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@65401.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_clock = clock; // @[:@65428.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_reset = reset; // @[:@65429.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_rPort_0_output_0 = x555_tmp_1_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@65826.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_rPort_0_output_0 = x554_tmp_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@65849.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_rPort_0_output_0 = x556_tmp_2_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@65934.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_done = x593_inr_UnitPipe_sm_io_done; // @[sm_x593_inr_UnitPipe.scala 147:22:@65963.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x593_inr_UnitPipe_sm_io_datapathEn & x593_inr_UnitPipe_mySignalsIn_mask; // @[sm_x593_inr_UnitPipe.scala 147:22:@65956.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_baseEn = _T_1043 & _T_1052; // @[sm_x593_inr_UnitPipe.scala 147:22:@65955.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_break = x593_inr_UnitPipe_sm_io_break; // @[sm_x593_inr_UnitPipe.scala 147:22:@65954.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x593_inr_UnitPipe.scala 146:18:@65944.4]
  assign x594_force_0_clock = clock; // @[:@65972.4]
  assign x594_force_0_reset = reset; // @[:@65973.4]
  assign x594_force_0_io_rPort_0_en_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@69017.4]
  assign x594_force_0_io_wPort_0_data_0 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@68294.4]
  assign x594_force_0_io_wPort_0_en_0 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@68290.4]
  assign x594_force_0_io_sEn_0 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_sEn_0; // @[MemInterfaceType.scala 189:41:@68281.4]
  assign x594_force_0_io_sEn_1 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_sEn_1; // @[MemInterfaceType.scala 189:41:@69006.4]
  assign x594_force_0_io_sDone_0 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_sDone_0; // @[MemInterfaceType.scala 189:64:@68282.4]
  assign x594_force_0_io_sDone_1 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_sDone_1; // @[MemInterfaceType.scala 189:64:@69007.4]
  assign x595_reg_clock = clock; // @[:@66002.4]
  assign x595_reg_reset = reset; // @[:@66003.4]
  assign x595_reg_io_wPort_0_data_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@66778.4]
  assign x595_reg_io_wPort_0_reset = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_reset; // @[MemInterfaceType.scala 67:44:@66777.4]
  assign x595_reg_io_wPort_0_en_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@66774.4]
  assign x595_reg_io_sEn_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_sEn_0; // @[MemInterfaceType.scala 189:41:@66764.4]
  assign x595_reg_io_sEn_1 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_sEn_1; // @[MemInterfaceType.scala 189:41:@67599.4]
  assign x595_reg_io_sDone_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_sDone_0; // @[MemInterfaceType.scala 189:64:@66765.4]
  assign x595_reg_io_sDone_1 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_sDone_1; // @[MemInterfaceType.scala 189:64:@67600.4]
  assign x596_reg_clock = clock; // @[:@66039.4]
  assign x596_reg_reset = reset; // @[:@66040.4]
  assign x596_reg_io_wPort_0_data_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@66819.4]
  assign x596_reg_io_wPort_0_reset = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_reset; // @[MemInterfaceType.scala 67:44:@66818.4]
  assign x596_reg_io_wPort_0_en_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@66815.4]
  assign x596_reg_io_sEn_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_sEn_0; // @[MemInterfaceType.scala 189:41:@66806.4]
  assign x596_reg_io_sEn_1 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x596_reg_sEn_1; // @[MemInterfaceType.scala 189:41:@67640.4]
  assign x596_reg_io_sDone_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_sDone_0; // @[MemInterfaceType.scala 189:64:@66807.4]
  assign x596_reg_io_sDone_1 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x596_reg_sDone_1; // @[MemInterfaceType.scala 189:64:@67641.4]
  assign x605_inr_UnitPipe_sm_clock = clock; // @[:@66105.4]
  assign x605_inr_UnitPipe_sm_reset = reset; // @[:@66106.4]
  assign x605_inr_UnitPipe_sm_io_enable = _T_1150 & _T_1159; // @[SpatialBlocks.scala 139:18:@66203.4]
  assign x605_inr_UnitPipe_sm_io_ctrDone = x605_inr_UnitPipe_sm_io_ctrInc & _T_1126; // @[sm_x653_outr_Reduce.scala 145:39:@66136.4]
  assign x605_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 141:21:@66205.4]
  assign x605_inr_UnitPipe_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@66177.4]
  assign x605_inr_UnitPipe_sm_io_break = 1'h0; // @[sm_x653_outr_Reduce.scala 151:37:@66163.4]
  assign RetimeWrapper_11_clock = clock; // @[:@66138.4]
  assign RetimeWrapper_11_reset = reset; // @[:@66139.4]
  assign RetimeWrapper_11_io_flow = x605_inr_UnitPipe_sm_io_backpressure; // @[package.scala 95:18:@66141.4]
  assign RetimeWrapper_11_io_in = x605_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@66140.4]
  assign RetimeWrapper_12_clock = clock; // @[:@66148.4]
  assign RetimeWrapper_12_reset = reset; // @[:@66149.4]
  assign RetimeWrapper_12_io_flow = x605_inr_UnitPipe_sm_io_backpressure; // @[package.scala 95:18:@66151.4]
  assign RetimeWrapper_12_io_in = x605_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@66150.4]
  assign RetimeWrapper_13_clock = clock; // @[:@66184.4]
  assign RetimeWrapper_13_reset = reset; // @[:@66185.4]
  assign RetimeWrapper_13_io_flow = 1'h1; // @[package.scala 95:18:@66187.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@66186.4]
  assign RetimeWrapper_14_clock = clock; // @[:@66192.4]
  assign RetimeWrapper_14_reset = reset; // @[:@66193.4]
  assign RetimeWrapper_14_io_flow = 1'h1; // @[package.scala 95:18:@66195.4]
  assign RetimeWrapper_14_io_in = x605_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@66194.4]
  assign x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_clock = clock; // @[:@66221.4]
  assign x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_reset = reset; // @[:@66222.4]
  assign x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_rPort_0_output_0 = x580_r_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@66751.4]
  assign x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_done = x605_inr_UnitPipe_sm_io_done; // @[sm_x605_inr_UnitPipe.scala 142:22:@66846.4]
  assign x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x605_inr_UnitPipe_sm_io_datapathEn & x605_inr_UnitPipe_mySignalsIn_mask; // @[sm_x605_inr_UnitPipe.scala 142:22:@66839.4]
  assign x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_baseEn = _T_1150 & _T_1159; // @[sm_x605_inr_UnitPipe.scala 142:22:@66838.4]
  assign x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_break = x605_inr_UnitPipe_sm_io_break; // @[sm_x605_inr_UnitPipe.scala 142:22:@66837.4]
  assign x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x605_inr_UnitPipe.scala 141:18:@66827.4]
  assign x621_inr_Switch_sm_clock = clock; // @[:@66924.4]
  assign x621_inr_Switch_sm_reset = reset; // @[:@66925.4]
  assign x621_inr_Switch_sm_io_enable = _T_1279 & _T_1288; // @[SpatialBlocks.scala 139:18:@67032.4]
  assign x621_inr_Switch_sm_io_parentAck = io_sigsIn_smChildAcks_3; // @[SpatialBlocks.scala 141:21:@67034.4]
  assign x621_inr_Switch_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@67006.4]
  assign x621_inr_Switch_sm_io_doneIn_0 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@67002.4]
  assign x621_inr_Switch_sm_io_doneIn_1 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:72:@67003.4]
  assign x621_inr_Switch_sm_io_selectsIn_0 = x595_reg_io_rPort_0_output_0; // @[sm_x653_outr_Reduce.scala 168:46:@66958.4]
  assign x621_inr_Switch_sm_io_selectsIn_1 = x596_reg_io_rPort_0_output_0; // @[sm_x653_outr_Reduce.scala 169:46:@66959.4]
  assign RetimeWrapper_15_clock = clock; // @[:@66961.4]
  assign RetimeWrapper_15_reset = reset; // @[:@66962.4]
  assign RetimeWrapper_15_io_flow = x621_inr_Switch_sm_io_backpressure; // @[package.scala 95:18:@66964.4]
  assign RetimeWrapper_15_io_in = x621_inr_Switch_sm_io_done; // @[package.scala 94:16:@66963.4]
  assign RetimeWrapper_16_clock = clock; // @[:@66971.4]
  assign RetimeWrapper_16_reset = reset; // @[:@66972.4]
  assign RetimeWrapper_16_io_flow = x621_inr_Switch_sm_io_backpressure; // @[package.scala 95:18:@66974.4]
  assign RetimeWrapper_16_io_in = x621_inr_Switch_sm_io_done; // @[package.scala 94:16:@66973.4]
  assign RetimeWrapper_17_clock = clock; // @[:@67013.4]
  assign RetimeWrapper_17_reset = reset; // @[:@67014.4]
  assign RetimeWrapper_17_io_flow = 1'h1; // @[package.scala 95:18:@67016.4]
  assign RetimeWrapper_17_io_in = io_sigsIn_smEnableOuts_3; // @[package.scala 94:16:@67015.4]
  assign RetimeWrapper_18_clock = clock; // @[:@67021.4]
  assign RetimeWrapper_18_reset = reset; // @[:@67022.4]
  assign RetimeWrapper_18_io_flow = 1'h1; // @[package.scala 95:18:@67024.4]
  assign RetimeWrapper_18_io_in = x621_inr_Switch_sm_io_done; // @[package.scala 94:16:@67023.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_clock = clock; // @[:@67050.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_reset = reset; // @[:@67051.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x736_rd_x596 = x596_reg_io_rPort_0_output_0; // @[sm_x621_inr_Switch.scala 70:31:@67549.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_rPort_1_output_0 = x580_r_0_io_rPort_1_output_0; // @[MemInterfaceType.scala 66:44:@67586.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_rPort_1_output_0 = x595_reg_io_rPort_1_output_0; // @[MemInterfaceType.scala 66:44:@67609.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x735_rd_x595 = x595_reg_io_rPort_0_output_0; // @[sm_x621_inr_Switch.scala 75:31:@67632.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_done = x621_inr_Switch_sm_io_done; // @[sm_x621_inr_Switch.scala 145:22:@67683.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_baseEn = _T_1279 & _T_1288; // @[sm_x621_inr_Switch.scala 145:22:@67675.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smSelectsOut_0 = x621_inr_Switch_sm_io_selectsOut_0; // @[sm_x621_inr_Switch.scala 145:22:@67669.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smSelectsOut_1 = x621_inr_Switch_sm_io_selectsOut_1; // @[sm_x621_inr_Switch.scala 145:22:@67670.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smChildAcks_0 = x621_inr_Switch_sm_io_childAck_0; // @[sm_x621_inr_Switch.scala 145:22:@67667.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smChildAcks_1 = x621_inr_Switch_sm_io_childAck_1; // @[sm_x621_inr_Switch.scala 145:22:@67668.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_rr = io_rr; // @[sm_x621_inr_Switch.scala 144:18:@67661.4]
  assign x623_inr_UnitPipe_sm_clock = clock; // @[:@67731.4]
  assign x623_inr_UnitPipe_sm_reset = reset; // @[:@67732.4]
  assign x623_inr_UnitPipe_sm_io_enable = _T_1383 & _T_1392; // @[SpatialBlocks.scala 139:18:@67829.4]
  assign x623_inr_UnitPipe_sm_io_ctrDone = x623_inr_UnitPipe_sm_io_ctrInc & _T_1359; // @[sm_x653_outr_Reduce.scala 181:39:@67762.4]
  assign x623_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_4; // @[SpatialBlocks.scala 141:21:@67831.4]
  assign x623_inr_UnitPipe_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@67803.4]
  assign x623_inr_UnitPipe_sm_io_break = 1'h0; // @[sm_x653_outr_Reduce.scala 187:37:@67789.4]
  assign RetimeWrapper_19_clock = clock; // @[:@67764.4]
  assign RetimeWrapper_19_reset = reset; // @[:@67765.4]
  assign RetimeWrapper_19_io_flow = x623_inr_UnitPipe_sm_io_backpressure; // @[package.scala 95:18:@67767.4]
  assign RetimeWrapper_19_io_in = x623_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@67766.4]
  assign RetimeWrapper_20_clock = clock; // @[:@67774.4]
  assign RetimeWrapper_20_reset = reset; // @[:@67775.4]
  assign RetimeWrapper_20_io_flow = x623_inr_UnitPipe_sm_io_backpressure; // @[package.scala 95:18:@67777.4]
  assign RetimeWrapper_20_io_in = x623_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@67776.4]
  assign RetimeWrapper_21_clock = clock; // @[:@67810.4]
  assign RetimeWrapper_21_reset = reset; // @[:@67811.4]
  assign RetimeWrapper_21_io_flow = 1'h1; // @[package.scala 95:18:@67813.4]
  assign RetimeWrapper_21_io_in = io_sigsIn_smEnableOuts_4; // @[package.scala 94:16:@67812.4]
  assign RetimeWrapper_22_clock = clock; // @[:@67818.4]
  assign RetimeWrapper_22_reset = reset; // @[:@67819.4]
  assign RetimeWrapper_22_io_flow = 1'h1; // @[package.scala 95:18:@67821.4]
  assign RetimeWrapper_22_io_in = x623_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@67820.4]
  assign x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_clock = clock; // @[:@67847.4]
  assign x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_reset = reset; // @[:@67848.4]
  assign x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x621_inr_Switch_number = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_ret_number; // @[sm_x623_inr_UnitPipe.scala 70:34:@68297.4]
  assign x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_done = x623_inr_UnitPipe_sm_io_done; // @[sm_x623_inr_UnitPipe.scala 115:22:@68358.4]
  assign x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x623_inr_UnitPipe_sm_io_datapathEn & x623_inr_UnitPipe_mySignalsIn_mask; // @[sm_x623_inr_UnitPipe.scala 115:22:@68351.4]
  assign x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_baseEn = _T_1383 & _T_1392; // @[sm_x623_inr_UnitPipe.scala 115:22:@68350.4]
  assign x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_break = x623_inr_UnitPipe_sm_io_break; // @[sm_x623_inr_UnitPipe.scala 115:22:@68349.4]
  assign x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x623_inr_UnitPipe.scala 114:18:@68339.4]
  assign x625_ctrchain_clock = clock; // @[:@68367.4]
  assign x625_ctrchain_reset = reset; // @[:@68368.4]
  assign x625_ctrchain_io_input_reset = x639_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@68550.4]
  assign x625_ctrchain_io_input_enable = x639_inr_Foreach_sm_io_ctrInc & x639_inr_Foreach_mySignalsIn_iiDone; // @[SpatialBlocks.scala 158:42:@68549.4]
  assign x639_inr_Foreach_sm_clock = clock; // @[:@68420.4]
  assign x639_inr_Foreach_sm_reset = reset; // @[:@68421.4]
  assign x639_inr_Foreach_sm_io_enable = _T_1489 & _T_1498; // @[SpatialBlocks.scala 139:18:@68529.4]
  assign x639_inr_Foreach_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 133:15:@68504.4]
  assign x639_inr_Foreach_sm_io_ctrDone = io_rr ? _T_1464 : 1'h0; // @[sm_x653_outr_Reduce.scala 196:38:@68456.4]
  assign x639_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_5; // @[SpatialBlocks.scala 141:21:@68531.4]
  assign x639_inr_Foreach_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@68503.4]
  assign x639_inr_Foreach_sm_io_break = 1'h0; // @[sm_x653_outr_Reduce.scala 202:36:@68483.4]
  assign x639_inr_Foreach_iiCtr_clock = clock; // @[:@68445.4]
  assign x639_inr_Foreach_iiCtr_reset = reset; // @[:@68446.4]
  assign x639_inr_Foreach_iiCtr_io_input_enable = _T_1500 & _T_1501; // @[SpatialBlocks.scala 157:27:@68538.4]
  assign x639_inr_Foreach_iiCtr_io_input_reset = x639_inr_Foreach_sm_io_rst | x639_inr_Foreach_sm_io_parentAck; // @[SpatialBlocks.scala 157:63:@68540.4]
  assign RetimeWrapper_23_clock = clock; // @[:@68449.4]
  assign RetimeWrapper_23_reset = reset; // @[:@68450.4]
  assign RetimeWrapper_23_io_flow = 1'h1; // @[package.scala 95:18:@68452.4]
  assign RetimeWrapper_23_io_in = x625_ctrchain_io_output_done; // @[package.scala 94:16:@68451.4]
  assign RetimeWrapper_24_clock = clock; // @[:@68458.4]
  assign RetimeWrapper_24_reset = reset; // @[:@68459.4]
  assign RetimeWrapper_24_io_flow = x639_inr_Foreach_sm_io_backpressure; // @[package.scala 95:18:@68461.4]
  assign RetimeWrapper_24_io_in = x639_inr_Foreach_sm_io_done; // @[package.scala 94:16:@68460.4]
  assign RetimeWrapper_25_clock = clock; // @[:@68468.4]
  assign RetimeWrapper_25_reset = reset; // @[:@68469.4]
  assign RetimeWrapper_25_io_flow = x639_inr_Foreach_sm_io_backpressure; // @[package.scala 95:18:@68471.4]
  assign RetimeWrapper_25_io_in = x639_inr_Foreach_sm_io_done; // @[package.scala 94:16:@68470.4]
  assign RetimeWrapper_26_clock = clock; // @[:@68510.4]
  assign RetimeWrapper_26_reset = reset; // @[:@68511.4]
  assign RetimeWrapper_26_io_flow = 1'h1; // @[package.scala 95:18:@68513.4]
  assign RetimeWrapper_26_io_in = io_sigsIn_smEnableOuts_5; // @[package.scala 94:16:@68512.4]
  assign RetimeWrapper_27_clock = clock; // @[:@68518.4]
  assign RetimeWrapper_27_reset = reset; // @[:@68519.4]
  assign RetimeWrapper_27_io_flow = 1'h1; // @[package.scala 95:18:@68521.4]
  assign RetimeWrapper_27_io_in = x639_inr_Foreach_sm_io_done; // @[package.scala 94:16:@68520.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_clock = clock; // @[:@68552.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_reset = reset; // @[:@68553.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_b552 = b552_chain_io_rPort_4_output_0; // @[sm_x639_inr_Foreach.scala 65:23:@68998.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_rPort_0_output_0 = x594_force_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@69015.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_output_0 = x557_tmp_3_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@69038.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_b543 = io_in_b543; // @[sm_x639_inr_Foreach.scala 69:23:@69075.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_done = x639_inr_Foreach_sm_io_done; // @[sm_x639_inr_Foreach.scala 164:22:@69099.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_iiIssue = x639_inr_Foreach_iiCtr_io_output_issue | _T_1504; // @[sm_x639_inr_Foreach.scala 164:22:@69096.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_1500 & _T_1501; // @[sm_x639_inr_Foreach.scala 164:22:@69092.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_baseEn = _T_1489 & _T_1498; // @[sm_x639_inr_Foreach.scala 164:22:@69091.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_break = x639_inr_Foreach_sm_io_break; // @[sm_x639_inr_Foreach.scala 164:22:@69090.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{28{x625_ctrchain_io_output_counts_0[3]}},x625_ctrchain_io_output_counts_0}; // @[sm_x639_inr_Foreach.scala 164:22:@69085.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x625_ctrchain_io_output_oobs_0; // @[sm_x639_inr_Foreach.scala 164:22:@69084.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x639_inr_Foreach.scala 163:18:@69080.4]
  assign x652_inr_Foreach_sm_clock = clock; // @[:@69144.4]
  assign x652_inr_Foreach_sm_reset = reset; // @[:@69145.4]
  assign x652_inr_Foreach_sm_io_enable = _T_1595 & _T_1604; // @[SpatialBlocks.scala 139:18:@69252.4]
  assign x652_inr_Foreach_sm_io_ctrDone = io_rr ? _T_1570 : 1'h0; // @[sm_x653_outr_Reduce.scala 207:38:@69180.4]
  assign x652_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_6; // @[SpatialBlocks.scala 141:21:@69254.4]
  assign x652_inr_Foreach_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@69226.4]
  assign x652_inr_Foreach_sm_io_break = 1'h0; // @[sm_x653_outr_Reduce.scala 213:36:@69207.4]
  assign RetimeWrapper_28_clock = clock; // @[:@69173.4]
  assign RetimeWrapper_28_reset = reset; // @[:@69174.4]
  assign RetimeWrapper_28_io_flow = 1'h1; // @[package.scala 95:18:@69176.4]
  assign RetimeWrapper_28_io_in = io_in_x549_ctrchain_output_done; // @[package.scala 94:16:@69175.4]
  assign RetimeWrapper_29_clock = clock; // @[:@69182.4]
  assign RetimeWrapper_29_reset = reset; // @[:@69183.4]
  assign RetimeWrapper_29_io_flow = x652_inr_Foreach_sm_io_backpressure; // @[package.scala 95:18:@69185.4]
  assign RetimeWrapper_29_io_in = x652_inr_Foreach_sm_io_done; // @[package.scala 94:16:@69184.4]
  assign RetimeWrapper_30_clock = clock; // @[:@69192.4]
  assign RetimeWrapper_30_reset = reset; // @[:@69193.4]
  assign RetimeWrapper_30_io_flow = x652_inr_Foreach_sm_io_backpressure; // @[package.scala 95:18:@69195.4]
  assign RetimeWrapper_30_io_in = x652_inr_Foreach_sm_io_done; // @[package.scala 94:16:@69194.4]
  assign RetimeWrapper_31_clock = clock; // @[:@69233.4]
  assign RetimeWrapper_31_reset = reset; // @[:@69234.4]
  assign RetimeWrapper_31_io_flow = 1'h1; // @[package.scala 95:18:@69236.4]
  assign RetimeWrapper_31_io_in = io_sigsIn_smEnableOuts_6; // @[package.scala 94:16:@69235.4]
  assign RetimeWrapper_32_clock = clock; // @[:@69241.4]
  assign RetimeWrapper_32_reset = reset; // @[:@69242.4]
  assign RetimeWrapper_32_io_flow = 1'h1; // @[package.scala 95:18:@69244.4]
  assign RetimeWrapper_32_io_in = x652_inr_Foreach_sm_io_done; // @[package.scala 94:16:@69243.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_clock = clock; // @[:@69275.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_reset = reset; // @[:@69276.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_b550_number = __6_io_result; // @[sm_x652_inr_Foreach.scala 58:23:@69487.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_output_0 = x558_tmp_4_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@69506.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_output_0 = io_in_x544_accum_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@69532.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_b543 = io_in_b543; // @[sm_x652_inr_Foreach.scala 62:23:@69544.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_done = x652_inr_Foreach_sm_io_done; // @[sm_x652_inr_Foreach.scala 136:22:@69568.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_1606 & _T_1607; // @[sm_x652_inr_Foreach.scala 136:22:@69561.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_baseEn = _T_1595 & _T_1604; // @[sm_x652_inr_Foreach.scala 136:22:@69560.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_break = x652_inr_Foreach_sm_io_break; // @[sm_x652_inr_Foreach.scala 136:22:@69559.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{28{io_in_x549_ctrchain_output_counts_0[3]}},io_in_x549_ctrchain_output_counts_0}; // @[sm_x652_inr_Foreach.scala 136:22:@69554.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = io_in_x549_ctrchain_output_oobs_0; // @[sm_x652_inr_Foreach.scala 136:22:@69553.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x652_inr_Foreach.scala 135:18:@69549.4]
  assign RetimeWrapper_33_clock = clock; // @[:@69578.4]
  assign RetimeWrapper_33_reset = reset; // @[:@69579.4]
  assign RetimeWrapper_33_io_flow = 1'h1; // @[package.scala 95:18:@69581.4]
  assign RetimeWrapper_33_io_in = io_sigsIn_done; // @[package.scala 94:16:@69580.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_789 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1019 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1126 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1359 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_789 <= 1'h0;
    end else begin
      _T_789 <= _T_786;
    end
    if (reset) begin
      _T_1019 <= 1'h0;
    end else begin
      _T_1019 <= _T_1016;
    end
    if (reset) begin
      _T_1126 <= 1'h0;
    end else begin
      _T_1126 <= _T_1123;
    end
    if (reset) begin
      _T_1359 <= 1'h0;
    end else begin
      _T_1359 <= _T_1356;
    end
  end
endmodule
module x667_inr_Foreach_kernelx667_inr_Foreach_concrete1( // @[:@71205.2]
  input         clock, // @[:@71206.4]
  input         reset, // @[:@71207.4]
  input  [31:0] io_in_b542_number, // @[:@71208.4]
  output [1:0]  io_in_x545_accum_1_rPort_0_ofs_0, // @[:@71208.4]
  output        io_in_x545_accum_1_rPort_0_en_0, // @[:@71208.4]
  input  [31:0] io_in_x545_accum_1_rPort_0_output_0, // @[:@71208.4]
  output        io_in_x545_accum_1_sEn_1, // @[:@71208.4]
  output        io_in_x545_accum_1_sDone_1, // @[:@71208.4]
  output [8:0]  io_in_x473_A_sram_2_rPort_0_ofs_0, // @[:@71208.4]
  output        io_in_x473_A_sram_2_rPort_0_en_0, // @[:@71208.4]
  input  [31:0] io_in_x473_A_sram_2_rPort_0_output_0, // @[:@71208.4]
  output [8:0]  io_in_x539_out_sram_0_wPort_0_ofs_0, // @[:@71208.4]
  output [31:0] io_in_x539_out_sram_0_wPort_0_data_0, // @[:@71208.4]
  output        io_in_x539_out_sram_0_wPort_0_en_0, // @[:@71208.4]
  input         io_in_b543, // @[:@71208.4]
  output [63:0] io_in_instrctrs_17_cycs, // @[:@71208.4]
  output [63:0] io_in_instrctrs_17_iters, // @[:@71208.4]
  input         io_sigsIn_done, // @[:@71208.4]
  input         io_sigsIn_datapathEn, // @[:@71208.4]
  input         io_sigsIn_baseEn, // @[:@71208.4]
  input         io_sigsIn_break, // @[:@71208.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@71208.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@71208.4]
  input         io_rr // @[:@71208.4]
);
  wire  cycles_x667_inr_Foreach_clock; // @[sm_x667_inr_Foreach.scala 77:43:@71366.4]
  wire  cycles_x667_inr_Foreach_reset; // @[sm_x667_inr_Foreach.scala 77:43:@71366.4]
  wire  cycles_x667_inr_Foreach_io_enable; // @[sm_x667_inr_Foreach.scala 77:43:@71366.4]
  wire [63:0] cycles_x667_inr_Foreach_io_count; // @[sm_x667_inr_Foreach.scala 77:43:@71366.4]
  wire  iters_x667_inr_Foreach_clock; // @[sm_x667_inr_Foreach.scala 78:42:@71369.4]
  wire  iters_x667_inr_Foreach_reset; // @[sm_x667_inr_Foreach.scala 78:42:@71369.4]
  wire  iters_x667_inr_Foreach_io_enable; // @[sm_x667_inr_Foreach.scala 78:42:@71369.4]
  wire [63:0] iters_x667_inr_Foreach_io_count; // @[sm_x667_inr_Foreach.scala 78:42:@71369.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@71386.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@71386.4]
  wire  x751_sum_1_clock; // @[Math.scala 150:24:@71422.4]
  wire  x751_sum_1_reset; // @[Math.scala 150:24:@71422.4]
  wire [31:0] x751_sum_1_io_a; // @[Math.scala 150:24:@71422.4]
  wire [31:0] x751_sum_1_io_b; // @[Math.scala 150:24:@71422.4]
  wire  x751_sum_1_io_flow; // @[Math.scala 150:24:@71422.4]
  wire [31:0] x751_sum_1_io_result; // @[Math.scala 150:24:@71422.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@71433.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@71433.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@71433.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@71433.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@71433.4]
  wire  x662_sum_1_clock; // @[Math.scala 150:24:@71442.4]
  wire  x662_sum_1_reset; // @[Math.scala 150:24:@71442.4]
  wire [31:0] x662_sum_1_io_a; // @[Math.scala 150:24:@71442.4]
  wire [31:0] x662_sum_1_io_b; // @[Math.scala 150:24:@71442.4]
  wire  x662_sum_1_io_flow; // @[Math.scala 150:24:@71442.4]
  wire [31:0] x662_sum_1_io_result; // @[Math.scala 150:24:@71442.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@71453.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@71453.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@71453.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@71453.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@71453.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@71463.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@71463.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@71463.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@71463.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@71463.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@71475.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@71475.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@71475.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@71475.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@71475.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@71487.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@71487.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@71487.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@71487.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@71487.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@71508.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@71508.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@71508.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@71508.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@71508.4]
  wire  x665_sum_1_clock; // @[Math.scala 150:24:@71517.4]
  wire  x665_sum_1_reset; // @[Math.scala 150:24:@71517.4]
  wire [31:0] x665_sum_1_io_a; // @[Math.scala 150:24:@71517.4]
  wire [31:0] x665_sum_1_io_b; // @[Math.scala 150:24:@71517.4]
  wire [31:0] x665_sum_1_io_result; // @[Math.scala 150:24:@71517.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@71528.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@71528.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@71528.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@71528.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@71528.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@71538.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@71538.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@71538.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@71538.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@71548.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@71548.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@71548.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@71548.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@71548.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@71562.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@71562.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@71562.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@71562.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@71562.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@71582.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@71582.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@71582.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@71582.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@71582.4]
  wire  _T_590; // @[package.scala 100:49:@71373.4]
  reg  _T_593; // @[package.scala 48:56:@71374.4]
  reg [31:0] _RAND_0;
  wire  b657; // @[sm_x667_inr_Foreach.scala 83:18:@71394.4]
  wire  _T_618; // @[sm_x667_inr_Foreach.scala 88:114:@71400.4]
  wire  _T_619; // @[sm_x667_inr_Foreach.scala 88:111:@71401.4]
  wire  _T_624; // @[implicits.scala 56:10:@71404.4]
  wire  _T_625; // @[sm_x667_inr_Foreach.scala 88:131:@71405.4]
  wire  _T_626; // @[sm_x667_inr_Foreach.scala 88:228:@71406.4]
  wire [32:0] _GEN_0; // @[Math.scala 461:32:@71418.4]
  wire [32:0] _T_632; // @[Math.scala 461:32:@71418.4]
  wire  _T_669; // @[package.scala 96:25:@71480.4 package.scala 96:25:@71481.4]
  wire  _T_671; // @[implicits.scala 56:10:@71482.4]
  wire  _T_673; // @[sm_x667_inr_Foreach.scala 109:111:@71484.4]
  wire  _T_678; // @[package.scala 96:25:@71492.4 package.scala 96:25:@71493.4]
  wire  _T_680; // @[implicits.scala 56:10:@71494.4]
  wire  _T_681; // @[sm_x667_inr_Foreach.scala 109:131:@71495.4]
  wire  x796_b657_D2; // @[package.scala 96:25:@71468.4 package.scala 96:25:@71469.4]
  wire  _T_682; // @[sm_x667_inr_Foreach.scala 109:228:@71496.4]
  wire  x795_b543_D2; // @[package.scala 96:25:@71458.4 package.scala 96:25:@71459.4]
  wire  _T_719; // @[package.scala 96:25:@71567.4 package.scala 96:25:@71568.4]
  wire  _T_721; // @[implicits.scala 56:10:@71569.4]
  wire  _T_722; // @[sm_x667_inr_Foreach.scala 128:120:@71570.4]
  wire  _T_724; // @[sm_x667_inr_Foreach.scala 128:217:@71572.4]
  wire  x800_b657_D5; // @[package.scala 96:25:@71553.4 package.scala 96:25:@71554.4]
  wire  _T_726; // @[sm_x667_inr_Foreach.scala 128:262:@71574.4]
  wire  x798_b543_D5; // @[package.scala 96:25:@71533.4 package.scala 96:25:@71534.4]
  wire  _T_731; // @[package.scala 96:25:@71587.4 package.scala 96:25:@71588.4]
  wire [31:0] b656_number; // @[Math.scala 723:22:@71391.4 Math.scala 724:14:@71392.4]
  wire [31:0] x662_sum_number; // @[Math.scala 154:22:@71448.4 Math.scala 155:14:@71449.4]
  wire [31:0] x799_x662_sum_D3_number; // @[package.scala 96:25:@71543.4 package.scala 96:25:@71544.4]
  InstrumentationCounter cycles_x667_inr_Foreach ( // @[sm_x667_inr_Foreach.scala 77:43:@71366.4]
    .clock(cycles_x667_inr_Foreach_clock),
    .reset(cycles_x667_inr_Foreach_reset),
    .io_enable(cycles_x667_inr_Foreach_io_enable),
    .io_count(cycles_x667_inr_Foreach_io_count)
  );
  InstrumentationCounter iters_x667_inr_Foreach ( // @[sm_x667_inr_Foreach.scala 78:42:@71369.4]
    .clock(iters_x667_inr_Foreach_clock),
    .reset(iters_x667_inr_Foreach_reset),
    .io_enable(iters_x667_inr_Foreach_io_enable),
    .io_count(iters_x667_inr_Foreach_io_count)
  );
  _ _ ( // @[Math.scala 720:24:@71386.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x739_sum x751_sum_1 ( // @[Math.scala 150:24:@71422.4]
    .clock(x751_sum_1_clock),
    .reset(x751_sum_1_reset),
    .io_a(x751_sum_1_io_a),
    .io_b(x751_sum_1_io_b),
    .io_flow(x751_sum_1_io_flow),
    .io_result(x751_sum_1_io_result)
  );
  RetimeWrapper_32 RetimeWrapper ( // @[package.scala 93:22:@71433.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x739_sum x662_sum_1 ( // @[Math.scala 150:24:@71442.4]
    .clock(x662_sum_1_clock),
    .reset(x662_sum_1_reset),
    .io_a(x662_sum_1_io_a),
    .io_b(x662_sum_1_io_b),
    .io_flow(x662_sum_1_io_flow),
    .io_result(x662_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@71453.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@71463.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@71475.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@71487.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_45 RetimeWrapper_5 ( // @[package.scala 93:22:@71508.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  x648_sum x665_sum_1 ( // @[Math.scala 150:24:@71517.4]
    .clock(x665_sum_1_clock),
    .reset(x665_sum_1_reset),
    .io_a(x665_sum_1_io_a),
    .io_b(x665_sum_1_io_b),
    .io_result(x665_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_6 ( // @[package.scala 93:22:@71528.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_718 RetimeWrapper_7 ( // @[package.scala 93:22:@71538.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_8 ( // @[package.scala 93:22:@71548.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_9 ( // @[package.scala 93:22:@71562.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@71582.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_590 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@71373.4]
  assign b657 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x667_inr_Foreach.scala 83:18:@71394.4]
  assign _T_618 = ~ io_sigsIn_break; // @[sm_x667_inr_Foreach.scala 88:114:@71400.4]
  assign _T_619 = io_rr & _T_618; // @[sm_x667_inr_Foreach.scala 88:111:@71401.4]
  assign _T_624 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 56:10:@71404.4]
  assign _T_625 = _T_619 & _T_624; // @[sm_x667_inr_Foreach.scala 88:131:@71405.4]
  assign _T_626 = _T_625 & b657; // @[sm_x667_inr_Foreach.scala 88:228:@71406.4]
  assign _GEN_0 = {{1'd0}, io_in_b542_number}; // @[Math.scala 461:32:@71418.4]
  assign _T_632 = _GEN_0 << 1; // @[Math.scala 461:32:@71418.4]
  assign _T_669 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@71480.4 package.scala 96:25:@71481.4]
  assign _T_671 = io_rr ? _T_669 : 1'h0; // @[implicits.scala 56:10:@71482.4]
  assign _T_673 = _T_671 & _T_618; // @[sm_x667_inr_Foreach.scala 109:111:@71484.4]
  assign _T_678 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@71492.4 package.scala 96:25:@71493.4]
  assign _T_680 = io_rr ? _T_678 : 1'h0; // @[implicits.scala 56:10:@71494.4]
  assign _T_681 = _T_673 & _T_680; // @[sm_x667_inr_Foreach.scala 109:131:@71495.4]
  assign x796_b657_D2 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@71468.4 package.scala 96:25:@71469.4]
  assign _T_682 = _T_681 & x796_b657_D2; // @[sm_x667_inr_Foreach.scala 109:228:@71496.4]
  assign x795_b543_D2 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@71458.4 package.scala 96:25:@71459.4]
  assign _T_719 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@71567.4 package.scala 96:25:@71568.4]
  assign _T_721 = io_rr ? _T_719 : 1'h0; // @[implicits.scala 56:10:@71569.4]
  assign _T_722 = _T_618 & _T_721; // @[sm_x667_inr_Foreach.scala 128:120:@71570.4]
  assign _T_724 = _T_722 & _T_618; // @[sm_x667_inr_Foreach.scala 128:217:@71572.4]
  assign x800_b657_D5 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@71553.4 package.scala 96:25:@71554.4]
  assign _T_726 = _T_724 & x800_b657_D5; // @[sm_x667_inr_Foreach.scala 128:262:@71574.4]
  assign x798_b543_D5 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@71533.4 package.scala 96:25:@71534.4]
  assign _T_731 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@71587.4 package.scala 96:25:@71588.4]
  assign b656_number = __io_result; // @[Math.scala 723:22:@71391.4 Math.scala 724:14:@71392.4]
  assign x662_sum_number = x662_sum_1_io_result; // @[Math.scala 154:22:@71448.4 Math.scala 155:14:@71449.4]
  assign x799_x662_sum_D3_number = RetimeWrapper_7_io_out; // @[package.scala 96:25:@71543.4 package.scala 96:25:@71544.4]
  assign io_in_x545_accum_1_rPort_0_ofs_0 = b656_number[1:0]; // @[MemInterfaceType.scala 107:54:@71410.4]
  assign io_in_x545_accum_1_rPort_0_en_0 = _T_626 & io_in_b543; // @[MemInterfaceType.scala 110:79:@71412.4]
  assign io_in_x545_accum_1_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@71590.4]
  assign io_in_x545_accum_1_sDone_1 = io_rr ? _T_731 : 1'h0; // @[MemInterfaceType.scala 197:17:@71591.4]
  assign io_in_x473_A_sram_2_rPort_0_ofs_0 = x662_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@71500.4]
  assign io_in_x473_A_sram_2_rPort_0_en_0 = _T_682 & x795_b543_D2; // @[MemInterfaceType.scala 110:79:@71502.4]
  assign io_in_x539_out_sram_0_wPort_0_ofs_0 = x799_x662_sum_D3_number[8:0]; // @[MemInterfaceType.scala 89:54:@71577.4]
  assign io_in_x539_out_sram_0_wPort_0_data_0 = x665_sum_1_io_result; // @[MemInterfaceType.scala 90:56:@71578.4]
  assign io_in_x539_out_sram_0_wPort_0_en_0 = _T_726 & x798_b543_D5; // @[MemInterfaceType.scala 93:57:@71580.4]
  assign io_in_instrctrs_17_cycs = cycles_x667_inr_Foreach_io_count; // @[Ledger.scala 293:21:@71378.4]
  assign io_in_instrctrs_17_iters = iters_x667_inr_Foreach_io_count; // @[Ledger.scala 294:22:@71379.4]
  assign cycles_x667_inr_Foreach_clock = clock; // @[:@71367.4]
  assign cycles_x667_inr_Foreach_reset = reset; // @[:@71368.4]
  assign cycles_x667_inr_Foreach_io_enable = io_sigsIn_baseEn; // @[sm_x667_inr_Foreach.scala 79:41:@71372.4]
  assign iters_x667_inr_Foreach_clock = clock; // @[:@71370.4]
  assign iters_x667_inr_Foreach_reset = reset; // @[:@71371.4]
  assign iters_x667_inr_Foreach_io_enable = io_sigsIn_done & _T_593; // @[sm_x667_inr_Foreach.scala 80:40:@71377.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@71389.4]
  assign x751_sum_1_clock = clock; // @[:@71423.4]
  assign x751_sum_1_reset = reset; // @[:@71424.4]
  assign x751_sum_1_io_a = _T_632[31:0]; // @[Math.scala 151:17:@71425.4]
  assign x751_sum_1_io_b = io_in_b542_number; // @[Math.scala 152:17:@71426.4]
  assign x751_sum_1_io_flow = 1'h1; // @[Math.scala 153:20:@71427.4]
  assign RetimeWrapper_clock = clock; // @[:@71434.4]
  assign RetimeWrapper_reset = reset; // @[:@71435.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@71437.4]
  assign RetimeWrapper_io_in = __io_result; // @[package.scala 94:16:@71436.4]
  assign x662_sum_1_clock = clock; // @[:@71443.4]
  assign x662_sum_1_reset = reset; // @[:@71444.4]
  assign x662_sum_1_io_a = x751_sum_1_io_result; // @[Math.scala 151:17:@71445.4]
  assign x662_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@71446.4]
  assign x662_sum_1_io_flow = 1'h1; // @[Math.scala 153:20:@71447.4]
  assign RetimeWrapper_1_clock = clock; // @[:@71454.4]
  assign RetimeWrapper_1_reset = reset; // @[:@71455.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@71457.4]
  assign RetimeWrapper_1_io_in = io_in_b543; // @[package.scala 94:16:@71456.4]
  assign RetimeWrapper_2_clock = clock; // @[:@71464.4]
  assign RetimeWrapper_2_reset = reset; // @[:@71465.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@71467.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@71466.4]
  assign RetimeWrapper_3_clock = clock; // @[:@71476.4]
  assign RetimeWrapper_3_reset = reset; // @[:@71477.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@71479.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@71478.4]
  assign RetimeWrapper_4_clock = clock; // @[:@71488.4]
  assign RetimeWrapper_4_reset = reset; // @[:@71489.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@71491.4]
  assign RetimeWrapper_4_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@71490.4]
  assign RetimeWrapper_5_clock = clock; // @[:@71509.4]
  assign RetimeWrapper_5_reset = reset; // @[:@71510.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@71512.4]
  assign RetimeWrapper_5_io_in = io_in_x545_accum_1_rPort_0_output_0; // @[package.scala 94:16:@71511.4]
  assign x665_sum_1_clock = clock; // @[:@71518.4]
  assign x665_sum_1_reset = reset; // @[:@71519.4]
  assign x665_sum_1_io_a = RetimeWrapper_5_io_out; // @[Math.scala 151:17:@71520.4]
  assign x665_sum_1_io_b = io_in_x473_A_sram_2_rPort_0_output_0; // @[Math.scala 152:17:@71521.4]
  assign RetimeWrapper_6_clock = clock; // @[:@71529.4]
  assign RetimeWrapper_6_reset = reset; // @[:@71530.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@71532.4]
  assign RetimeWrapper_6_io_in = io_in_b543; // @[package.scala 94:16:@71531.4]
  assign RetimeWrapper_7_clock = clock; // @[:@71539.4]
  assign RetimeWrapper_7_reset = reset; // @[:@71540.4]
  assign RetimeWrapper_7_io_in = x662_sum_1_io_result; // @[package.scala 94:16:@71541.4]
  assign RetimeWrapper_8_clock = clock; // @[:@71549.4]
  assign RetimeWrapper_8_reset = reset; // @[:@71550.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@71552.4]
  assign RetimeWrapper_8_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@71551.4]
  assign RetimeWrapper_9_clock = clock; // @[:@71563.4]
  assign RetimeWrapper_9_reset = reset; // @[:@71564.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@71566.4]
  assign RetimeWrapper_9_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@71565.4]
  assign RetimeWrapper_10_clock = clock; // @[:@71583.4]
  assign RetimeWrapper_10_reset = reset; // @[:@71584.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@71586.4]
  assign RetimeWrapper_10_io_in = io_sigsIn_done; // @[package.scala 94:16:@71585.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_593 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_593 <= 1'h0;
    end else begin
      _T_593 <= _T_590;
    end
  end
endmodule
module x668_outr_Foreach_kernelx668_outr_Foreach_concrete1( // @[:@71593.2]
  input         clock, // @[:@71594.4]
  input         reset, // @[:@71595.4]
  output [8:0]  io_in_x472_A_sram_1_rPort_0_ofs_0, // @[:@71596.4]
  output        io_in_x472_A_sram_1_rPort_0_en_0, // @[:@71596.4]
  input  [31:0] io_in_x472_A_sram_1_rPort_0_output_0, // @[:@71596.4]
  output [8:0]  io_in_x471_A_sram_0_rPort_0_ofs_0, // @[:@71596.4]
  output        io_in_x471_A_sram_0_rPort_0_en_0, // @[:@71596.4]
  input  [31:0] io_in_x471_A_sram_0_rPort_0_output_0, // @[:@71596.4]
  output [8:0]  io_in_x473_A_sram_2_rPort_0_ofs_0, // @[:@71596.4]
  output        io_in_x473_A_sram_2_rPort_0_en_0, // @[:@71596.4]
  input  [31:0] io_in_x473_A_sram_2_rPort_0_output_0, // @[:@71596.4]
  output [8:0]  io_in_x539_out_sram_0_wPort_0_ofs_0, // @[:@71596.4]
  output [31:0] io_in_x539_out_sram_0_wPort_0_data_0, // @[:@71596.4]
  output        io_in_x539_out_sram_0_wPort_0_en_0, // @[:@71596.4]
  output [63:0] io_in_instrctrs_6_cycs, // @[:@71596.4]
  output [63:0] io_in_instrctrs_6_iters, // @[:@71596.4]
  output [63:0] io_in_instrctrs_7_cycs, // @[:@71596.4]
  output [63:0] io_in_instrctrs_7_iters, // @[:@71596.4]
  output [63:0] io_in_instrctrs_8_cycs, // @[:@71596.4]
  output [63:0] io_in_instrctrs_8_iters, // @[:@71596.4]
  output [63:0] io_in_instrctrs_9_cycs, // @[:@71596.4]
  output [63:0] io_in_instrctrs_9_iters, // @[:@71596.4]
  output [63:0] io_in_instrctrs_10_cycs, // @[:@71596.4]
  output [63:0] io_in_instrctrs_10_iters, // @[:@71596.4]
  output [63:0] io_in_instrctrs_11_cycs, // @[:@71596.4]
  output [63:0] io_in_instrctrs_11_iters, // @[:@71596.4]
  output [63:0] io_in_instrctrs_12_cycs, // @[:@71596.4]
  output [63:0] io_in_instrctrs_12_iters, // @[:@71596.4]
  output [63:0] io_in_instrctrs_13_cycs, // @[:@71596.4]
  output [63:0] io_in_instrctrs_13_iters, // @[:@71596.4]
  output [63:0] io_in_instrctrs_14_cycs, // @[:@71596.4]
  output [63:0] io_in_instrctrs_14_iters, // @[:@71596.4]
  output [63:0] io_in_instrctrs_15_cycs, // @[:@71596.4]
  output [63:0] io_in_instrctrs_15_iters, // @[:@71596.4]
  output [63:0] io_in_instrctrs_16_cycs, // @[:@71596.4]
  output [63:0] io_in_instrctrs_16_iters, // @[:@71596.4]
  output [63:0] io_in_instrctrs_17_cycs, // @[:@71596.4]
  output [63:0] io_in_instrctrs_17_iters, // @[:@71596.4]
  input         io_sigsIn_done, // @[:@71596.4]
  input         io_sigsIn_baseEn, // @[:@71596.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@71596.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@71596.4]
  input         io_sigsIn_smChildAcks_0, // @[:@71596.4]
  input         io_sigsIn_smChildAcks_1, // @[:@71596.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@71596.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@71596.4]
  output        io_sigsOut_smDoneIn_0, // @[:@71596.4]
  output        io_sigsOut_smDoneIn_1, // @[:@71596.4]
  output        io_sigsOut_smMaskIn_0, // @[:@71596.4]
  output        io_sigsOut_smMaskIn_1, // @[:@71596.4]
  input         io_rr // @[:@71596.4]
);
  wire  cycles_x668_outr_Foreach_clock; // @[sm_x668_outr_Foreach.scala 70:44:@71756.4]
  wire  cycles_x668_outr_Foreach_reset; // @[sm_x668_outr_Foreach.scala 70:44:@71756.4]
  wire  cycles_x668_outr_Foreach_io_enable; // @[sm_x668_outr_Foreach.scala 70:44:@71756.4]
  wire [63:0] cycles_x668_outr_Foreach_io_count; // @[sm_x668_outr_Foreach.scala 70:44:@71756.4]
  wire  iters_x668_outr_Foreach_clock; // @[sm_x668_outr_Foreach.scala 71:43:@71759.4]
  wire  iters_x668_outr_Foreach_reset; // @[sm_x668_outr_Foreach.scala 71:43:@71759.4]
  wire  iters_x668_outr_Foreach_io_enable; // @[sm_x668_outr_Foreach.scala 71:43:@71759.4]
  wire [63:0] iters_x668_outr_Foreach_io_count; // @[sm_x668_outr_Foreach.scala 71:43:@71759.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@71776.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@71776.4]
  wire  b542_chain_clock; // @[sm_x668_outr_Foreach.scala 76:30:@71784.4]
  wire  b542_chain_reset; // @[sm_x668_outr_Foreach.scala 76:30:@71784.4]
  wire [31:0] b542_chain_io_rPort_0_output_0; // @[sm_x668_outr_Foreach.scala 76:30:@71784.4]
  wire [31:0] b542_chain_io_wPort_0_data_0; // @[sm_x668_outr_Foreach.scala 76:30:@71784.4]
  wire  b542_chain_io_wPort_0_reset; // @[sm_x668_outr_Foreach.scala 76:30:@71784.4]
  wire  b542_chain_io_wPort_0_en_0; // @[sm_x668_outr_Foreach.scala 76:30:@71784.4]
  wire  b542_chain_io_sEn_0; // @[sm_x668_outr_Foreach.scala 76:30:@71784.4]
  wire  b542_chain_io_sEn_1; // @[sm_x668_outr_Foreach.scala 76:30:@71784.4]
  wire  b542_chain_io_sDone_0; // @[sm_x668_outr_Foreach.scala 76:30:@71784.4]
  wire  b542_chain_io_sDone_1; // @[sm_x668_outr_Foreach.scala 76:30:@71784.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@71813.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@71813.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@71813.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@71813.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@71813.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@71825.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@71825.4]
  wire  b543_chain_clock; // @[sm_x668_outr_Foreach.scala 80:30:@71834.4]
  wire  b543_chain_reset; // @[sm_x668_outr_Foreach.scala 80:30:@71834.4]
  wire  b543_chain_io_rPort_0_output_0; // @[sm_x668_outr_Foreach.scala 80:30:@71834.4]
  wire  b543_chain_io_wPort_0_data_0; // @[sm_x668_outr_Foreach.scala 80:30:@71834.4]
  wire  b543_chain_io_wPort_0_reset; // @[sm_x668_outr_Foreach.scala 80:30:@71834.4]
  wire  b543_chain_io_wPort_0_en_0; // @[sm_x668_outr_Foreach.scala 80:30:@71834.4]
  wire  b543_chain_io_sEn_0; // @[sm_x668_outr_Foreach.scala 80:30:@71834.4]
  wire  b543_chain_io_sEn_1; // @[sm_x668_outr_Foreach.scala 80:30:@71834.4]
  wire  b543_chain_io_sDone_0; // @[sm_x668_outr_Foreach.scala 80:30:@71834.4]
  wire  b543_chain_io_sDone_1; // @[sm_x668_outr_Foreach.scala 80:30:@71834.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@71863.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@71863.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@71863.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@71863.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@71863.4]
  wire  x544_accum_0_clock; // @[m_x544_accum_0.scala 27:22:@71873.4]
  wire  x544_accum_0_reset; // @[m_x544_accum_0.scala 27:22:@71873.4]
  wire [1:0] x544_accum_0_io_rPort_0_ofs_0; // @[m_x544_accum_0.scala 27:22:@71873.4]
  wire  x544_accum_0_io_rPort_0_en_0; // @[m_x544_accum_0.scala 27:22:@71873.4]
  wire [31:0] x544_accum_0_io_rPort_0_output_0; // @[m_x544_accum_0.scala 27:22:@71873.4]
  wire [1:0] x544_accum_0_io_wPort_0_ofs_0; // @[m_x544_accum_0.scala 27:22:@71873.4]
  wire [31:0] x544_accum_0_io_wPort_0_data_0; // @[m_x544_accum_0.scala 27:22:@71873.4]
  wire  x544_accum_0_io_wPort_0_en_0; // @[m_x544_accum_0.scala 27:22:@71873.4]
  wire  x545_accum_1_clock; // @[m_x545_accum_1.scala 27:22:@71890.4]
  wire  x545_accum_1_reset; // @[m_x545_accum_1.scala 27:22:@71890.4]
  wire [1:0] x545_accum_1_io_rPort_0_ofs_0; // @[m_x545_accum_1.scala 27:22:@71890.4]
  wire  x545_accum_1_io_rPort_0_en_0; // @[m_x545_accum_1.scala 27:22:@71890.4]
  wire [31:0] x545_accum_1_io_rPort_0_output_0; // @[m_x545_accum_1.scala 27:22:@71890.4]
  wire [1:0] x545_accum_1_io_wPort_0_ofs_0; // @[m_x545_accum_1.scala 27:22:@71890.4]
  wire [31:0] x545_accum_1_io_wPort_0_data_0; // @[m_x545_accum_1.scala 27:22:@71890.4]
  wire  x545_accum_1_io_wPort_0_en_0; // @[m_x545_accum_1.scala 27:22:@71890.4]
  wire  x545_accum_1_io_sEn_0; // @[m_x545_accum_1.scala 27:22:@71890.4]
  wire  x545_accum_1_io_sEn_1; // @[m_x545_accum_1.scala 27:22:@71890.4]
  wire  x545_accum_1_io_sDone_0; // @[m_x545_accum_1.scala 27:22:@71890.4]
  wire  x545_accum_1_io_sDone_1; // @[m_x545_accum_1.scala 27:22:@71890.4]
  wire  x547_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@71920.4]
  wire  x547_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@71920.4]
  wire  x547_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@71920.4]
  wire  x547_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@71920.4]
  wire [8:0] x547_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@71920.4]
  wire  x547_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@71920.4]
  wire  x547_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@71920.4]
  wire  x549_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@71937.4]
  wire  x549_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@71937.4]
  wire  x549_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@71937.4]
  wire  x549_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@71937.4]
  wire [3:0] x549_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@71937.4]
  wire  x549_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@71937.4]
  wire  x549_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@71937.4]
  wire  x653_outr_Reduce_sm_clock; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_reset; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_enable; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_done; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_ctrDone; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_ctrInc; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_ctrRst; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_parentAck; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_backpressure; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_doneIn_0; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_doneIn_1; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_doneIn_2; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_doneIn_3; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_doneIn_4; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_doneIn_5; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_doneIn_6; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_maskIn_0; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_maskIn_1; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_maskIn_2; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_maskIn_4; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_maskIn_5; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_enableOut_0; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_enableOut_1; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_enableOut_2; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_enableOut_3; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_enableOut_4; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_enableOut_5; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_enableOut_6; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_childAck_0; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_childAck_1; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_childAck_2; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_childAck_3; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_childAck_4; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_childAck_5; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  x653_outr_Reduce_sm_io_childAck_6; // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@72079.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@72079.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@72079.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@72079.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@72079.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@72088.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@72088.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@72088.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@72088.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@72088.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@72098.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@72098.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@72098.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@72098.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@72098.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@72169.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@72169.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@72169.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@72169.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@72169.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@72177.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@72177.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@72177.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@72177.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@72177.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_clock; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_reset; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [8:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_en_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [31:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_output_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [31:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_b542_number; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [8:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_en_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [31:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_output_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [1:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_ofs_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [31:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_data_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_en_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_sEn_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_sDone_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [1:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_ofs_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_en_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [31:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_output_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [1:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_ofs_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [31:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_data_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_en_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_input_reset; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_input_enable; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [3:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_counts_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_oobs_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_done; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_b543; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_7_cycs; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_7_iters; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_8_cycs; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_8_iters; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_9_cycs; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_9_iters; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_10_cycs; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_10_iters; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_11_cycs; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_11_iters; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_12_cycs; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_12_iters; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_13_cycs; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_13_iters; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_14_cycs; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_14_iters; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_15_cycs; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_15_iters; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_16_cycs; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [63:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_16_iters; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_done; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_baseEn; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_3; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_4; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_5; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_6; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_3; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_4; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_5; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_6; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire [31:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_3; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_4; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_5; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_6; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_0; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_1; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_2; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_4; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_5; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_rr; // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
  wire  x655_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@72598.4]
  wire  x655_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@72598.4]
  wire  x655_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@72598.4]
  wire  x655_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@72598.4]
  wire [3:0] x655_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@72598.4]
  wire  x655_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@72598.4]
  wire  x655_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@72598.4]
  wire  x667_inr_Foreach_sm_clock; // @[sm_x667_inr_Foreach.scala 35:18:@72651.4]
  wire  x667_inr_Foreach_sm_reset; // @[sm_x667_inr_Foreach.scala 35:18:@72651.4]
  wire  x667_inr_Foreach_sm_io_enable; // @[sm_x667_inr_Foreach.scala 35:18:@72651.4]
  wire  x667_inr_Foreach_sm_io_done; // @[sm_x667_inr_Foreach.scala 35:18:@72651.4]
  wire  x667_inr_Foreach_sm_io_ctrDone; // @[sm_x667_inr_Foreach.scala 35:18:@72651.4]
  wire  x667_inr_Foreach_sm_io_datapathEn; // @[sm_x667_inr_Foreach.scala 35:18:@72651.4]
  wire  x667_inr_Foreach_sm_io_ctrInc; // @[sm_x667_inr_Foreach.scala 35:18:@72651.4]
  wire  x667_inr_Foreach_sm_io_ctrRst; // @[sm_x667_inr_Foreach.scala 35:18:@72651.4]
  wire  x667_inr_Foreach_sm_io_parentAck; // @[sm_x667_inr_Foreach.scala 35:18:@72651.4]
  wire  x667_inr_Foreach_sm_io_backpressure; // @[sm_x667_inr_Foreach.scala 35:18:@72651.4]
  wire  x667_inr_Foreach_sm_io_break; // @[sm_x667_inr_Foreach.scala 35:18:@72651.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@72680.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@72680.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@72680.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@72680.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@72680.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@72689.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@72689.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@72689.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@72689.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@72689.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@72699.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@72699.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@72699.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@72699.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@72699.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@72740.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@72740.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@72740.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@72740.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@72740.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@72748.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@72748.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@72748.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@72748.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@72748.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_clock; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_reset; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire [31:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_b542_number; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire [1:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_ofs_0; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_en_0; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire [31:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_output_0; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_sEn_1; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_sDone_1; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire [8:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_ofs_0; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_en_0; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire [31:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_output_0; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire [8:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_ofs_0; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire [31:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_data_0; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_en_0; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_b543; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire [63:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_instrctrs_17_cycs; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire [63:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_instrctrs_17_iters; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_done; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire [31:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_rr; // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
  wire  _T_628; // @[package.scala 100:49:@71763.4]
  reg  _T_631; // @[package.scala 48:56:@71764.4]
  reg [31:0] _RAND_0;
  wire  b543_chain_read_1; // @[sm_x668_outr_Foreach.scala 82:61:@71872.4]
  wire  _T_722; // @[package.scala 96:25:@72084.4 package.scala 96:25:@72085.4]
  wire  _T_726; // @[package.scala 96:25:@72093.4 package.scala 96:25:@72094.4]
  wire  _T_730; // @[package.scala 96:25:@72103.4 package.scala 96:25:@72104.4]
  wire  _T_746; // @[package.scala 96:25:@72174.4 package.scala 96:25:@72175.4]
  wire  _T_752; // @[package.scala 96:25:@72182.4 package.scala 96:25:@72183.4]
  wire  _T_755; // @[SpatialBlocks.scala 137:99:@72185.4]
  wire  _T_829; // @[package.scala 96:25:@72685.4 package.scala 96:25:@72686.4]
  wire  _T_833; // @[package.scala 96:25:@72694.4 package.scala 96:25:@72695.4]
  wire  _T_837; // @[package.scala 96:25:@72704.4 package.scala 96:25:@72705.4]
  wire  _T_853; // @[package.scala 96:25:@72745.4 package.scala 96:25:@72746.4]
  wire  _T_859; // @[package.scala 96:25:@72753.4 package.scala 96:25:@72754.4]
  wire  _T_862; // @[SpatialBlocks.scala 137:99:@72756.4]
  wire  _T_864; // @[SpatialBlocks.scala 156:36:@72765.4]
  wire  _T_865; // @[SpatialBlocks.scala 156:78:@72766.4]
  InstrumentationCounter cycles_x668_outr_Foreach ( // @[sm_x668_outr_Foreach.scala 70:44:@71756.4]
    .clock(cycles_x668_outr_Foreach_clock),
    .reset(cycles_x668_outr_Foreach_reset),
    .io_enable(cycles_x668_outr_Foreach_io_enable),
    .io_count(cycles_x668_outr_Foreach_io_count)
  );
  InstrumentationCounter iters_x668_outr_Foreach ( // @[sm_x668_outr_Foreach.scala 71:43:@71759.4]
    .clock(iters_x668_outr_Foreach_clock),
    .reset(iters_x668_outr_Foreach_reset),
    .io_enable(iters_x668_outr_Foreach_io_enable),
    .io_count(iters_x668_outr_Foreach_io_count)
  );
  _ _ ( // @[Math.scala 720:24:@71776.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  b542_chain b542_chain ( // @[sm_x668_outr_Foreach.scala 76:30:@71784.4]
    .clock(b542_chain_clock),
    .reset(b542_chain_reset),
    .io_rPort_0_output_0(b542_chain_io_rPort_0_output_0),
    .io_wPort_0_data_0(b542_chain_io_wPort_0_data_0),
    .io_wPort_0_reset(b542_chain_io_wPort_0_reset),
    .io_wPort_0_en_0(b542_chain_io_wPort_0_en_0),
    .io_sEn_0(b542_chain_io_sEn_0),
    .io_sEn_1(b542_chain_io_sEn_1),
    .io_sDone_0(b542_chain_io_sDone_0),
    .io_sDone_1(b542_chain_io_sDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@71813.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  _ __1 ( // @[Math.scala 720:24:@71825.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  b543_chain b543_chain ( // @[sm_x668_outr_Foreach.scala 80:30:@71834.4]
    .clock(b543_chain_clock),
    .reset(b543_chain_reset),
    .io_rPort_0_output_0(b543_chain_io_rPort_0_output_0),
    .io_wPort_0_data_0(b543_chain_io_wPort_0_data_0),
    .io_wPort_0_reset(b543_chain_io_wPort_0_reset),
    .io_wPort_0_en_0(b543_chain_io_wPort_0_en_0),
    .io_sEn_0(b543_chain_io_sEn_0),
    .io_sEn_1(b543_chain_io_sEn_1),
    .io_sDone_0(b543_chain_io_sDone_0),
    .io_sDone_1(b543_chain_io_sDone_1)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@71863.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x544_accum_0 x544_accum_0 ( // @[m_x544_accum_0.scala 27:22:@71873.4]
    .clock(x544_accum_0_clock),
    .reset(x544_accum_0_reset),
    .io_rPort_0_ofs_0(x544_accum_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x544_accum_0_io_rPort_0_en_0),
    .io_rPort_0_output_0(x544_accum_0_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(x544_accum_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x544_accum_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x544_accum_0_io_wPort_0_en_0)
  );
  x545_accum_1 x545_accum_1 ( // @[m_x545_accum_1.scala 27:22:@71890.4]
    .clock(x545_accum_1_clock),
    .reset(x545_accum_1_reset),
    .io_rPort_0_ofs_0(x545_accum_1_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x545_accum_1_io_rPort_0_en_0),
    .io_rPort_0_output_0(x545_accum_1_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(x545_accum_1_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x545_accum_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(x545_accum_1_io_wPort_0_en_0),
    .io_sEn_0(x545_accum_1_io_sEn_0),
    .io_sEn_1(x545_accum_1_io_sEn_1),
    .io_sDone_0(x545_accum_1_io_sDone_0),
    .io_sDone_1(x545_accum_1_io_sDone_1)
  );
  x478_ctrchain x547_ctrchain ( // @[SpatialBlocks.scala 37:22:@71920.4]
    .clock(x547_ctrchain_clock),
    .reset(x547_ctrchain_reset),
    .io_input_reset(x547_ctrchain_io_input_reset),
    .io_input_enable(x547_ctrchain_io_input_enable),
    .io_output_counts_0(x547_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x547_ctrchain_io_output_oobs_0),
    .io_output_done(x547_ctrchain_io_output_done)
  );
  x549_ctrchain x549_ctrchain ( // @[SpatialBlocks.scala 37:22:@71937.4]
    .clock(x549_ctrchain_clock),
    .reset(x549_ctrchain_reset),
    .io_input_reset(x549_ctrchain_io_input_reset),
    .io_input_enable(x549_ctrchain_io_input_enable),
    .io_output_counts_0(x549_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x549_ctrchain_io_output_oobs_0),
    .io_output_done(x549_ctrchain_io_output_done)
  );
  x653_outr_Reduce_sm x653_outr_Reduce_sm ( // @[sm_x653_outr_Reduce.scala 36:18:@72020.4]
    .clock(x653_outr_Reduce_sm_clock),
    .reset(x653_outr_Reduce_sm_reset),
    .io_enable(x653_outr_Reduce_sm_io_enable),
    .io_done(x653_outr_Reduce_sm_io_done),
    .io_ctrDone(x653_outr_Reduce_sm_io_ctrDone),
    .io_ctrInc(x653_outr_Reduce_sm_io_ctrInc),
    .io_ctrRst(x653_outr_Reduce_sm_io_ctrRst),
    .io_parentAck(x653_outr_Reduce_sm_io_parentAck),
    .io_backpressure(x653_outr_Reduce_sm_io_backpressure),
    .io_doneIn_0(x653_outr_Reduce_sm_io_doneIn_0),
    .io_doneIn_1(x653_outr_Reduce_sm_io_doneIn_1),
    .io_doneIn_2(x653_outr_Reduce_sm_io_doneIn_2),
    .io_doneIn_3(x653_outr_Reduce_sm_io_doneIn_3),
    .io_doneIn_4(x653_outr_Reduce_sm_io_doneIn_4),
    .io_doneIn_5(x653_outr_Reduce_sm_io_doneIn_5),
    .io_doneIn_6(x653_outr_Reduce_sm_io_doneIn_6),
    .io_maskIn_0(x653_outr_Reduce_sm_io_maskIn_0),
    .io_maskIn_1(x653_outr_Reduce_sm_io_maskIn_1),
    .io_maskIn_2(x653_outr_Reduce_sm_io_maskIn_2),
    .io_maskIn_4(x653_outr_Reduce_sm_io_maskIn_4),
    .io_maskIn_5(x653_outr_Reduce_sm_io_maskIn_5),
    .io_enableOut_0(x653_outr_Reduce_sm_io_enableOut_0),
    .io_enableOut_1(x653_outr_Reduce_sm_io_enableOut_1),
    .io_enableOut_2(x653_outr_Reduce_sm_io_enableOut_2),
    .io_enableOut_3(x653_outr_Reduce_sm_io_enableOut_3),
    .io_enableOut_4(x653_outr_Reduce_sm_io_enableOut_4),
    .io_enableOut_5(x653_outr_Reduce_sm_io_enableOut_5),
    .io_enableOut_6(x653_outr_Reduce_sm_io_enableOut_6),
    .io_childAck_0(x653_outr_Reduce_sm_io_childAck_0),
    .io_childAck_1(x653_outr_Reduce_sm_io_childAck_1),
    .io_childAck_2(x653_outr_Reduce_sm_io_childAck_2),
    .io_childAck_3(x653_outr_Reduce_sm_io_childAck_3),
    .io_childAck_4(x653_outr_Reduce_sm_io_childAck_4),
    .io_childAck_5(x653_outr_Reduce_sm_io_childAck_5),
    .io_childAck_6(x653_outr_Reduce_sm_io_childAck_6)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@72079.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@72088.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@72098.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@72169.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@72177.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1 x653_outr_Reduce_kernelx653_outr_Reduce_concrete1 ( // @[sm_x653_outr_Reduce.scala 219:24:@72211.4]
    .clock(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_clock),
    .reset(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_reset),
    .io_in_x472_A_sram_1_rPort_0_ofs_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0),
    .io_in_x472_A_sram_1_rPort_0_en_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_en_0),
    .io_in_x472_A_sram_1_rPort_0_output_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_output_0),
    .io_in_b542_number(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_b542_number),
    .io_in_x471_A_sram_0_rPort_0_ofs_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0),
    .io_in_x471_A_sram_0_rPort_0_en_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_en_0),
    .io_in_x471_A_sram_0_rPort_0_output_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_output_0),
    .io_in_x545_accum_1_wPort_0_ofs_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_ofs_0),
    .io_in_x545_accum_1_wPort_0_data_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_data_0),
    .io_in_x545_accum_1_wPort_0_en_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_en_0),
    .io_in_x545_accum_1_sEn_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_sEn_0),
    .io_in_x545_accum_1_sDone_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_sDone_0),
    .io_in_x544_accum_0_rPort_0_ofs_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_ofs_0),
    .io_in_x544_accum_0_rPort_0_en_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_en_0),
    .io_in_x544_accum_0_rPort_0_output_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_output_0),
    .io_in_x544_accum_0_wPort_0_ofs_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_ofs_0),
    .io_in_x544_accum_0_wPort_0_data_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_data_0),
    .io_in_x544_accum_0_wPort_0_en_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_en_0),
    .io_in_x549_ctrchain_input_reset(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_input_reset),
    .io_in_x549_ctrchain_input_enable(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_input_enable),
    .io_in_x549_ctrchain_output_counts_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_counts_0),
    .io_in_x549_ctrchain_output_oobs_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_oobs_0),
    .io_in_x549_ctrchain_output_done(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_done),
    .io_in_b543(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_b543),
    .io_in_instrctrs_7_cycs(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_7_cycs),
    .io_in_instrctrs_7_iters(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_7_iters),
    .io_in_instrctrs_8_cycs(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_8_cycs),
    .io_in_instrctrs_8_iters(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_8_iters),
    .io_in_instrctrs_9_cycs(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_9_cycs),
    .io_in_instrctrs_9_iters(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_9_iters),
    .io_in_instrctrs_10_cycs(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_10_cycs),
    .io_in_instrctrs_10_iters(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_10_iters),
    .io_in_instrctrs_11_cycs(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_11_cycs),
    .io_in_instrctrs_11_iters(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_11_iters),
    .io_in_instrctrs_12_cycs(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_12_cycs),
    .io_in_instrctrs_12_iters(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_12_iters),
    .io_in_instrctrs_13_cycs(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_13_cycs),
    .io_in_instrctrs_13_iters(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_13_iters),
    .io_in_instrctrs_14_cycs(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_14_cycs),
    .io_in_instrctrs_14_iters(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_14_iters),
    .io_in_instrctrs_15_cycs(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_15_cycs),
    .io_in_instrctrs_15_iters(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_15_iters),
    .io_in_instrctrs_16_cycs(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_16_cycs),
    .io_in_instrctrs_16_iters(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_16_iters),
    .io_sigsIn_done(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smEnableOuts_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smEnableOuts_3(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_3),
    .io_sigsIn_smEnableOuts_4(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_4),
    .io_sigsIn_smEnableOuts_5(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_5),
    .io_sigsIn_smEnableOuts_6(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_6),
    .io_sigsIn_smChildAcks_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsIn_smChildAcks_3(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_3),
    .io_sigsIn_smChildAcks_4(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_4),
    .io_sigsIn_smChildAcks_5(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_5),
    .io_sigsIn_smChildAcks_6(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_6),
    .io_sigsIn_cchainOutputs_0_counts_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsOut_smDoneIn_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smDoneIn_3(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_3),
    .io_sigsOut_smDoneIn_4(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_4),
    .io_sigsOut_smDoneIn_5(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_5),
    .io_sigsOut_smDoneIn_6(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_6),
    .io_sigsOut_smMaskIn_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_0),
    .io_sigsOut_smMaskIn_1(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_1),
    .io_sigsOut_smMaskIn_2(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_2),
    .io_sigsOut_smMaskIn_4(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_4),
    .io_sigsOut_smMaskIn_5(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_5),
    .io_rr(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_rr)
  );
  x549_ctrchain x655_ctrchain ( // @[SpatialBlocks.scala 37:22:@72598.4]
    .clock(x655_ctrchain_clock),
    .reset(x655_ctrchain_reset),
    .io_input_reset(x655_ctrchain_io_input_reset),
    .io_input_enable(x655_ctrchain_io_input_enable),
    .io_output_counts_0(x655_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x655_ctrchain_io_output_oobs_0),
    .io_output_done(x655_ctrchain_io_output_done)
  );
  x579_inr_Foreach_sm x667_inr_Foreach_sm ( // @[sm_x667_inr_Foreach.scala 35:18:@72651.4]
    .clock(x667_inr_Foreach_sm_clock),
    .reset(x667_inr_Foreach_sm_reset),
    .io_enable(x667_inr_Foreach_sm_io_enable),
    .io_done(x667_inr_Foreach_sm_io_done),
    .io_ctrDone(x667_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x667_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x667_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x667_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x667_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x667_inr_Foreach_sm_io_backpressure),
    .io_break(x667_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@72680.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@72689.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@72699.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@72740.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 ( // @[package.scala 93:22:@72748.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1 x667_inr_Foreach_kernelx667_inr_Foreach_concrete1 ( // @[sm_x667_inr_Foreach.scala 131:24:@72782.4]
    .clock(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_clock),
    .reset(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_reset),
    .io_in_b542_number(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_b542_number),
    .io_in_x545_accum_1_rPort_0_ofs_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_ofs_0),
    .io_in_x545_accum_1_rPort_0_en_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_en_0),
    .io_in_x545_accum_1_rPort_0_output_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_output_0),
    .io_in_x545_accum_1_sEn_1(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_sEn_1),
    .io_in_x545_accum_1_sDone_1(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_sDone_1),
    .io_in_x473_A_sram_2_rPort_0_ofs_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_ofs_0),
    .io_in_x473_A_sram_2_rPort_0_en_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_en_0),
    .io_in_x473_A_sram_2_rPort_0_output_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_output_0),
    .io_in_x539_out_sram_0_wPort_0_ofs_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_ofs_0),
    .io_in_x539_out_sram_0_wPort_0_data_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_data_0),
    .io_in_x539_out_sram_0_wPort_0_en_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_en_0),
    .io_in_b543(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_b543),
    .io_in_instrctrs_17_cycs(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_instrctrs_17_cycs),
    .io_in_instrctrs_17_iters(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_instrctrs_17_iters),
    .io_sigsIn_done(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_datapathEn(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_rr)
  );
  assign _T_628 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@71763.4]
  assign b543_chain_read_1 = b543_chain_io_rPort_0_output_0; // @[sm_x668_outr_Foreach.scala 82:61:@71872.4]
  assign _T_722 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@72084.4 package.scala 96:25:@72085.4]
  assign _T_726 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@72093.4 package.scala 96:25:@72094.4]
  assign _T_730 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@72103.4 package.scala 96:25:@72104.4]
  assign _T_746 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@72174.4 package.scala 96:25:@72175.4]
  assign _T_752 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@72182.4 package.scala 96:25:@72183.4]
  assign _T_755 = ~ _T_752; // @[SpatialBlocks.scala 137:99:@72185.4]
  assign _T_829 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@72685.4 package.scala 96:25:@72686.4]
  assign _T_833 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@72694.4 package.scala 96:25:@72695.4]
  assign _T_837 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@72704.4 package.scala 96:25:@72705.4]
  assign _T_853 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@72745.4 package.scala 96:25:@72746.4]
  assign _T_859 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@72753.4 package.scala 96:25:@72754.4]
  assign _T_862 = ~ _T_859; // @[SpatialBlocks.scala 137:99:@72756.4]
  assign _T_864 = x667_inr_Foreach_sm_io_datapathEn & b543_chain_read_1; // @[SpatialBlocks.scala 156:36:@72765.4]
  assign _T_865 = ~ x667_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 156:78:@72766.4]
  assign io_in_x472_A_sram_1_rPort_0_ofs_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@72450.4]
  assign io_in_x472_A_sram_1_rPort_0_en_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@72449.4]
  assign io_in_x471_A_sram_0_rPort_0_ofs_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@72456.4]
  assign io_in_x471_A_sram_0_rPort_0_en_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@72455.4]
  assign io_in_x473_A_sram_2_rPort_0_ofs_0 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@72988.4]
  assign io_in_x473_A_sram_2_rPort_0_en_0 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@72987.4]
  assign io_in_x539_out_sram_0_wPort_0_ofs_0 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@72995.4]
  assign io_in_x539_out_sram_0_wPort_0_data_0 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@72994.4]
  assign io_in_x539_out_sram_0_wPort_0_en_0 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@72990.4]
  assign io_in_instrctrs_6_cycs = cycles_x668_outr_Foreach_io_count; // @[Ledger.scala 293:21:@71768.4]
  assign io_in_instrctrs_6_iters = iters_x668_outr_Foreach_io_count; // @[Ledger.scala 294:22:@71769.4]
  assign io_in_instrctrs_7_cycs = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_7_cycs; // @[Ledger.scala 302:78:@72504.4]
  assign io_in_instrctrs_7_iters = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_7_iters; // @[Ledger.scala 302:78:@72503.4]
  assign io_in_instrctrs_8_cycs = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_8_cycs; // @[Ledger.scala 302:78:@72508.4]
  assign io_in_instrctrs_8_iters = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_8_iters; // @[Ledger.scala 302:78:@72507.4]
  assign io_in_instrctrs_9_cycs = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_9_cycs; // @[Ledger.scala 302:78:@72512.4]
  assign io_in_instrctrs_9_iters = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_9_iters; // @[Ledger.scala 302:78:@72511.4]
  assign io_in_instrctrs_10_cycs = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_10_cycs; // @[Ledger.scala 302:78:@72516.4]
  assign io_in_instrctrs_10_iters = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_10_iters; // @[Ledger.scala 302:78:@72515.4]
  assign io_in_instrctrs_11_cycs = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_11_cycs; // @[Ledger.scala 302:78:@72520.4]
  assign io_in_instrctrs_11_iters = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_11_iters; // @[Ledger.scala 302:78:@72519.4]
  assign io_in_instrctrs_12_cycs = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_12_cycs; // @[Ledger.scala 302:78:@72524.4]
  assign io_in_instrctrs_12_iters = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_12_iters; // @[Ledger.scala 302:78:@72523.4]
  assign io_in_instrctrs_13_cycs = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_13_cycs; // @[Ledger.scala 302:78:@72528.4]
  assign io_in_instrctrs_13_iters = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_13_iters; // @[Ledger.scala 302:78:@72527.4]
  assign io_in_instrctrs_14_cycs = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_14_cycs; // @[Ledger.scala 302:78:@72532.4]
  assign io_in_instrctrs_14_iters = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_14_iters; // @[Ledger.scala 302:78:@72531.4]
  assign io_in_instrctrs_15_cycs = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_15_cycs; // @[Ledger.scala 302:78:@72536.4]
  assign io_in_instrctrs_15_iters = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_15_iters; // @[Ledger.scala 302:78:@72535.4]
  assign io_in_instrctrs_16_cycs = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_16_cycs; // @[Ledger.scala 302:78:@72540.4]
  assign io_in_instrctrs_16_iters = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_instrctrs_16_iters; // @[Ledger.scala 302:78:@72539.4]
  assign io_in_instrctrs_17_cycs = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_instrctrs_17_cycs; // @[Ledger.scala 302:78:@73001.4]
  assign io_in_instrctrs_17_iters = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_instrctrs_17_iters; // @[Ledger.scala 302:78:@73000.4]
  assign io_sigsOut_smDoneIn_0 = x653_outr_Reduce_sm_io_done; // @[SpatialBlocks.scala 155:56:@72192.4]
  assign io_sigsOut_smDoneIn_1 = x667_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@72763.4]
  assign io_sigsOut_smMaskIn_0 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[SpatialBlocks.scala 155:86:@72193.4]
  assign io_sigsOut_smMaskIn_1 = b543_chain_io_rPort_0_output_0; // @[SpatialBlocks.scala 155:86:@72764.4]
  assign cycles_x668_outr_Foreach_clock = clock; // @[:@71757.4]
  assign cycles_x668_outr_Foreach_reset = reset; // @[:@71758.4]
  assign cycles_x668_outr_Foreach_io_enable = io_sigsIn_baseEn; // @[sm_x668_outr_Foreach.scala 72:42:@71762.4]
  assign iters_x668_outr_Foreach_clock = clock; // @[:@71760.4]
  assign iters_x668_outr_Foreach_reset = reset; // @[:@71761.4]
  assign iters_x668_outr_Foreach_io_enable = io_sigsIn_done & _T_631; // @[sm_x668_outr_Foreach.scala 73:41:@71767.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@71779.4]
  assign b542_chain_clock = clock; // @[:@71785.4]
  assign b542_chain_reset = reset; // @[:@71786.4]
  assign b542_chain_io_wPort_0_data_0 = __io_result; // @[NBuffers.scala 309:54:@71811.4]
  assign b542_chain_io_wPort_0_reset = RetimeWrapper_io_out; // @[NBuffers.scala 312:23:@71820.4]
  assign b542_chain_io_wPort_0_en_0 = io_sigsOut_smDoneIn_0; // @[NBuffers.scala 311:25:@71812.4]
  assign b542_chain_io_sEn_0 = _T_746 & _T_755; // @[NBuffers.scala 302:18:@72096.4]
  assign b542_chain_io_sEn_1 = _T_853 & _T_862; // @[NBuffers.scala 302:18:@72697.4]
  assign b542_chain_io_sDone_0 = io_rr ? _T_726 : 1'h0; // @[NBuffers.scala 303:20:@72097.4]
  assign b542_chain_io_sDone_1 = io_rr ? _T_833 : 1'h0; // @[NBuffers.scala 303:20:@72698.4]
  assign RetimeWrapper_clock = clock; // @[:@71814.4]
  assign RetimeWrapper_reset = reset; // @[:@71815.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@71817.4]
  assign RetimeWrapper_io_in = b542_chain_reset; // @[package.scala 94:16:@71816.4]
  assign __1_io_b = b542_chain_io_rPort_0_output_0; // @[Math.scala 721:17:@71828.4]
  assign b543_chain_clock = clock; // @[:@71835.4]
  assign b543_chain_reset = reset; // @[:@71836.4]
  assign b543_chain_io_wPort_0_data_0 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[NBuffers.scala 308:54:@71861.4]
  assign b543_chain_io_wPort_0_reset = RetimeWrapper_1_io_out; // @[NBuffers.scala 312:23:@71870.4]
  assign b543_chain_io_wPort_0_en_0 = io_sigsOut_smDoneIn_0; // @[NBuffers.scala 311:25:@71862.4]
  assign b543_chain_io_sEn_0 = _T_746 & _T_755; // @[NBuffers.scala 302:18:@72106.4]
  assign b543_chain_io_sEn_1 = _T_853 & _T_862; // @[NBuffers.scala 302:18:@72707.4]
  assign b543_chain_io_sDone_0 = io_rr ? _T_730 : 1'h0; // @[NBuffers.scala 303:20:@72107.4]
  assign b543_chain_io_sDone_1 = io_rr ? _T_837 : 1'h0; // @[NBuffers.scala 303:20:@72708.4]
  assign RetimeWrapper_1_clock = clock; // @[:@71864.4]
  assign RetimeWrapper_1_reset = reset; // @[:@71865.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@71867.4]
  assign RetimeWrapper_1_io_in = b543_chain_reset; // @[package.scala 94:16:@71866.4]
  assign x544_accum_0_clock = clock; // @[:@71874.4]
  assign x544_accum_0_reset = reset; // @[:@71875.4]
  assign x544_accum_0_io_rPort_0_ofs_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@72484.4]
  assign x544_accum_0_io_rPort_0_en_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@72483.4]
  assign x544_accum_0_io_wPort_0_ofs_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@72491.4]
  assign x544_accum_0_io_wPort_0_data_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@72490.4]
  assign x544_accum_0_io_wPort_0_en_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@72486.4]
  assign x545_accum_1_clock = clock; // @[:@71891.4]
  assign x545_accum_1_reset = reset; // @[:@71892.4]
  assign x545_accum_1_io_rPort_0_ofs_0 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@72983.4]
  assign x545_accum_1_io_rPort_0_en_0 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@72982.4]
  assign x545_accum_1_io_wPort_0_ofs_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@72479.4]
  assign x545_accum_1_io_wPort_0_data_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@72478.4]
  assign x545_accum_1_io_wPort_0_en_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@72474.4]
  assign x545_accum_1_io_sEn_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_sEn_0; // @[MemInterfaceType.scala 189:41:@72465.4]
  assign x545_accum_1_io_sEn_1 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_sEn_1; // @[MemInterfaceType.scala 189:41:@72971.4]
  assign x545_accum_1_io_sDone_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_sDone_0; // @[MemInterfaceType.scala 189:64:@72466.4]
  assign x545_accum_1_io_sDone_1 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_sDone_1; // @[MemInterfaceType.scala 189:64:@72972.4]
  assign x547_ctrchain_clock = clock; // @[:@71921.4]
  assign x547_ctrchain_reset = reset; // @[:@71922.4]
  assign x547_ctrchain_io_input_reset = x653_outr_Reduce_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@72210.4]
  assign x547_ctrchain_io_input_enable = x653_outr_Reduce_sm_io_ctrInc; // @[SpatialBlocks.scala 158:42:@72209.4]
  assign x549_ctrchain_clock = clock; // @[:@71938.4]
  assign x549_ctrchain_reset = reset; // @[:@71939.4]
  assign x549_ctrchain_io_input_reset = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_input_reset; // @[sm_x653_outr_Reduce.scala 68:38:@72494.4]
  assign x549_ctrchain_io_input_enable = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_input_enable; // @[sm_x653_outr_Reduce.scala 68:38:@72493.4]
  assign x653_outr_Reduce_sm_clock = clock; // @[:@72021.4]
  assign x653_outr_Reduce_sm_reset = reset; // @[:@72022.4]
  assign x653_outr_Reduce_sm_io_enable = _T_746 & _T_755; // @[SpatialBlocks.scala 139:18:@72189.4]
  assign x653_outr_Reduce_sm_io_ctrDone = io_rr ? _T_722 : 1'h0; // @[sm_x668_outr_Foreach.scala 94:38:@72087.4]
  assign x653_outr_Reduce_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@72191.4]
  assign x653_outr_Reduce_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@72163.4]
  assign x653_outr_Reduce_sm_io_doneIn_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@72149.4]
  assign x653_outr_Reduce_sm_io_doneIn_1 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:72:@72150.4]
  assign x653_outr_Reduce_sm_io_doneIn_2 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:72:@72151.4]
  assign x653_outr_Reduce_sm_io_doneIn_3 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_3; // @[SpatialBlocks.scala 130:72:@72152.4]
  assign x653_outr_Reduce_sm_io_doneIn_4 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_4; // @[SpatialBlocks.scala 130:72:@72153.4]
  assign x653_outr_Reduce_sm_io_doneIn_5 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_5; // @[SpatialBlocks.scala 130:72:@72154.4]
  assign x653_outr_Reduce_sm_io_doneIn_6 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_6; // @[SpatialBlocks.scala 130:72:@72155.4]
  assign x653_outr_Reduce_sm_io_maskIn_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_0; // @[SpatialBlocks.scala 131:72:@72156.4]
  assign x653_outr_Reduce_sm_io_maskIn_1 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_1; // @[SpatialBlocks.scala 131:72:@72157.4]
  assign x653_outr_Reduce_sm_io_maskIn_2 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_2; // @[SpatialBlocks.scala 131:72:@72158.4]
  assign x653_outr_Reduce_sm_io_maskIn_4 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_4; // @[SpatialBlocks.scala 131:72:@72160.4]
  assign x653_outr_Reduce_sm_io_maskIn_5 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_5; // @[SpatialBlocks.scala 131:72:@72161.4]
  assign RetimeWrapper_2_clock = clock; // @[:@72080.4]
  assign RetimeWrapper_2_reset = reset; // @[:@72081.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@72083.4]
  assign RetimeWrapper_2_io_in = x547_ctrchain_io_output_done; // @[package.scala 94:16:@72082.4]
  assign RetimeWrapper_3_clock = clock; // @[:@72089.4]
  assign RetimeWrapper_3_reset = reset; // @[:@72090.4]
  assign RetimeWrapper_3_io_flow = x653_outr_Reduce_sm_io_backpressure; // @[package.scala 95:18:@72092.4]
  assign RetimeWrapper_3_io_in = x653_outr_Reduce_sm_io_done; // @[package.scala 94:16:@72091.4]
  assign RetimeWrapper_4_clock = clock; // @[:@72099.4]
  assign RetimeWrapper_4_reset = reset; // @[:@72100.4]
  assign RetimeWrapper_4_io_flow = x653_outr_Reduce_sm_io_backpressure; // @[package.scala 95:18:@72102.4]
  assign RetimeWrapper_4_io_in = x653_outr_Reduce_sm_io_done; // @[package.scala 94:16:@72101.4]
  assign RetimeWrapper_5_clock = clock; // @[:@72170.4]
  assign RetimeWrapper_5_reset = reset; // @[:@72171.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@72173.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@72172.4]
  assign RetimeWrapper_6_clock = clock; // @[:@72178.4]
  assign RetimeWrapper_6_reset = reset; // @[:@72179.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@72181.4]
  assign RetimeWrapper_6_io_in = x653_outr_Reduce_sm_io_done; // @[package.scala 94:16:@72180.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_clock = clock; // @[:@72212.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_reset = reset; // @[:@72213.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_output_0 = io_in_x472_A_sram_1_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@72447.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_b542_number = __io_result; // @[sm_x653_outr_Reduce.scala 64:23:@72452.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_output_0 = io_in_x471_A_sram_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@72453.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_output_0 = x544_accum_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@72481.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_counts_0 = x549_ctrchain_io_output_counts_0; // @[sm_x653_outr_Reduce.scala 68:96:@72499.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_oobs_0 = x549_ctrchain_io_output_oobs_0; // @[sm_x653_outr_Reduce.scala 68:96:@72498.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_done = x549_ctrchain_io_output_done; // @[sm_x653_outr_Reduce.scala 68:96:@72496.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_b543 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x653_outr_Reduce.scala 69:23:@72500.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_done = x653_outr_Reduce_sm_io_done; // @[sm_x653_outr_Reduce.scala 225:22:@72578.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_baseEn = _T_746 & _T_755; // @[sm_x653_outr_Reduce.scala 225:22:@72570.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_0 = x653_outr_Reduce_sm_io_enableOut_0; // @[sm_x653_outr_Reduce.scala 225:22:@72561.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_1 = x653_outr_Reduce_sm_io_enableOut_1; // @[sm_x653_outr_Reduce.scala 225:22:@72562.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_2 = x653_outr_Reduce_sm_io_enableOut_2; // @[sm_x653_outr_Reduce.scala 225:22:@72563.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_3 = x653_outr_Reduce_sm_io_enableOut_3; // @[sm_x653_outr_Reduce.scala 225:22:@72564.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_4 = x653_outr_Reduce_sm_io_enableOut_4; // @[sm_x653_outr_Reduce.scala 225:22:@72565.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_5 = x653_outr_Reduce_sm_io_enableOut_5; // @[sm_x653_outr_Reduce.scala 225:22:@72566.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_6 = x653_outr_Reduce_sm_io_enableOut_6; // @[sm_x653_outr_Reduce.scala 225:22:@72567.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_0 = x653_outr_Reduce_sm_io_childAck_0; // @[sm_x653_outr_Reduce.scala 225:22:@72547.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_1 = x653_outr_Reduce_sm_io_childAck_1; // @[sm_x653_outr_Reduce.scala 225:22:@72548.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_2 = x653_outr_Reduce_sm_io_childAck_2; // @[sm_x653_outr_Reduce.scala 225:22:@72549.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_3 = x653_outr_Reduce_sm_io_childAck_3; // @[sm_x653_outr_Reduce.scala 225:22:@72550.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_4 = x653_outr_Reduce_sm_io_childAck_4; // @[sm_x653_outr_Reduce.scala 225:22:@72551.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_5 = x653_outr_Reduce_sm_io_childAck_5; // @[sm_x653_outr_Reduce.scala 225:22:@72552.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_6 = x653_outr_Reduce_sm_io_childAck_6; // @[sm_x653_outr_Reduce.scala 225:22:@72553.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{23{x547_ctrchain_io_output_counts_0[8]}},x547_ctrchain_io_output_counts_0}; // @[sm_x653_outr_Reduce.scala 225:22:@72546.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x547_ctrchain_io_output_oobs_0; // @[sm_x653_outr_Reduce.scala 225:22:@72545.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_rr = io_rr; // @[sm_x653_outr_Reduce.scala 224:18:@72541.4]
  assign x655_ctrchain_clock = clock; // @[:@72599.4]
  assign x655_ctrchain_reset = reset; // @[:@72600.4]
  assign x655_ctrchain_io_input_reset = x667_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@72781.4]
  assign x655_ctrchain_io_input_enable = x667_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 158:42:@72780.4]
  assign x667_inr_Foreach_sm_clock = clock; // @[:@72652.4]
  assign x667_inr_Foreach_sm_reset = reset; // @[:@72653.4]
  assign x667_inr_Foreach_sm_io_enable = _T_853 & _T_862; // @[SpatialBlocks.scala 139:18:@72760.4]
  assign x667_inr_Foreach_sm_io_ctrDone = io_rr ? _T_829 : 1'h0; // @[sm_x668_outr_Foreach.scala 109:38:@72688.4]
  assign x667_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 141:21:@72762.4]
  assign x667_inr_Foreach_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@72734.4]
  assign x667_inr_Foreach_sm_io_break = 1'h0; // @[sm_x668_outr_Foreach.scala 115:36:@72715.4]
  assign RetimeWrapper_7_clock = clock; // @[:@72681.4]
  assign RetimeWrapper_7_reset = reset; // @[:@72682.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@72684.4]
  assign RetimeWrapper_7_io_in = x655_ctrchain_io_output_done; // @[package.scala 94:16:@72683.4]
  assign RetimeWrapper_8_clock = clock; // @[:@72690.4]
  assign RetimeWrapper_8_reset = reset; // @[:@72691.4]
  assign RetimeWrapper_8_io_flow = x667_inr_Foreach_sm_io_backpressure; // @[package.scala 95:18:@72693.4]
  assign RetimeWrapper_8_io_in = x667_inr_Foreach_sm_io_done; // @[package.scala 94:16:@72692.4]
  assign RetimeWrapper_9_clock = clock; // @[:@72700.4]
  assign RetimeWrapper_9_reset = reset; // @[:@72701.4]
  assign RetimeWrapper_9_io_flow = x667_inr_Foreach_sm_io_backpressure; // @[package.scala 95:18:@72703.4]
  assign RetimeWrapper_9_io_in = x667_inr_Foreach_sm_io_done; // @[package.scala 94:16:@72702.4]
  assign RetimeWrapper_10_clock = clock; // @[:@72741.4]
  assign RetimeWrapper_10_reset = reset; // @[:@72742.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@72744.4]
  assign RetimeWrapper_10_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@72743.4]
  assign RetimeWrapper_11_clock = clock; // @[:@72749.4]
  assign RetimeWrapper_11_reset = reset; // @[:@72750.4]
  assign RetimeWrapper_11_io_flow = 1'h1; // @[package.scala 95:18:@72752.4]
  assign RetimeWrapper_11_io_in = x667_inr_Foreach_sm_io_done; // @[package.scala 94:16:@72751.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_clock = clock; // @[:@72783.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_reset = reset; // @[:@72784.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_b542_number = __1_io_result; // @[sm_x667_inr_Foreach.scala 58:23:@72963.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_output_0 = x545_accum_1_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@72980.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_output_0 = io_in_x473_A_sram_2_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@72985.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_b543 = b543_chain_io_rPort_0_output_0; // @[sm_x667_inr_Foreach.scala 62:23:@72997.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_done = x667_inr_Foreach_sm_io_done; // @[sm_x667_inr_Foreach.scala 137:22:@73021.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_864 & _T_865; // @[sm_x667_inr_Foreach.scala 137:22:@73014.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_baseEn = _T_853 & _T_862; // @[sm_x667_inr_Foreach.scala 137:22:@73013.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_break = x667_inr_Foreach_sm_io_break; // @[sm_x667_inr_Foreach.scala 137:22:@73012.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{28{x655_ctrchain_io_output_counts_0[3]}},x655_ctrchain_io_output_counts_0}; // @[sm_x667_inr_Foreach.scala 137:22:@73007.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x655_ctrchain_io_output_oobs_0; // @[sm_x667_inr_Foreach.scala 137:22:@73006.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x667_inr_Foreach.scala 136:18:@73002.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_631 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_631 <= 1'h0;
    end else begin
      _T_631 <= _T_628;
    end
  end
endmodule
module x724_outr_UnitPipe_DenseTransfer_sm( // @[:@73229.2]
  input   clock, // @[:@73230.4]
  input   reset, // @[:@73231.4]
  input   io_enable, // @[:@73232.4]
  output  io_done, // @[:@73232.4]
  input   io_parentAck, // @[:@73232.4]
  input   io_doneIn_0, // @[:@73232.4]
  output  io_enableOut_0, // @[:@73232.4]
  output  io_childAck_0, // @[:@73232.4]
  input   io_ctrCopyDone_0 // @[:@73232.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@73235.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@73235.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@73235.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@73235.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@73235.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@73235.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@73238.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@73238.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@73238.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@73238.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@73238.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@73238.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@73255.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@73255.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@73255.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@73255.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@73255.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@73255.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@73286.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@73286.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@73286.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@73286.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@73286.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@73300.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@73300.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@73300.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@73300.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@73300.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@73318.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@73318.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@73318.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@73318.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@73318.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@73355.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@73355.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@73355.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@73355.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@73355.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@73372.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@73372.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@73372.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@73372.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@73372.4]
  wire  _T_105; // @[Controllers.scala 165:35:@73270.4]
  wire  _T_107; // @[Controllers.scala 165:60:@73271.4]
  wire  _T_108; // @[Controllers.scala 165:58:@73272.4]
  wire  _T_110; // @[Controllers.scala 165:76:@73273.4]
  wire  _T_111; // @[Controllers.scala 165:74:@73274.4]
  wire  _T_115; // @[Controllers.scala 165:109:@73277.4]
  wire  _T_118; // @[Controllers.scala 165:141:@73279.4]
  wire  _T_126; // @[package.scala 96:25:@73291.4 package.scala 96:25:@73292.4]
  wire  _T_130; // @[Controllers.scala 167:54:@73294.4]
  wire  _T_131; // @[Controllers.scala 167:52:@73295.4]
  wire  _T_138; // @[package.scala 96:25:@73305.4 package.scala 96:25:@73306.4]
  wire  _T_156; // @[package.scala 96:25:@73323.4 package.scala 96:25:@73324.4]
  wire  _T_160; // @[Controllers.scala 169:67:@73326.4]
  wire  _T_161; // @[Controllers.scala 169:86:@73327.4]
  wire  _T_174; // @[Controllers.scala 213:68:@73341.4]
  wire  _T_176; // @[Controllers.scala 213:90:@73343.4]
  wire  _T_178; // @[Controllers.scala 213:132:@73345.4]
  reg  _T_186; // @[package.scala 48:56:@73351.4]
  reg [31:0] _RAND_0;
  wire  _T_187; // @[package.scala 100:41:@73353.4]
  reg  _T_200; // @[package.scala 48:56:@73369.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@73235.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@73238.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@73255.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@73286.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@73300.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@73318.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@73355.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@73372.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_105 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@73270.4]
  assign _T_107 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@73271.4]
  assign _T_108 = _T_105 & _T_107; // @[Controllers.scala 165:58:@73272.4]
  assign _T_110 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@73273.4]
  assign _T_111 = _T_108 & _T_110; // @[Controllers.scala 165:74:@73274.4]
  assign _T_115 = _T_111 & io_enable; // @[Controllers.scala 165:109:@73277.4]
  assign _T_118 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@73279.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@73291.4 package.scala 96:25:@73292.4]
  assign _T_130 = _T_126 == 1'h0; // @[Controllers.scala 167:54:@73294.4]
  assign _T_131 = io_doneIn_0 | _T_130; // @[Controllers.scala 167:52:@73295.4]
  assign _T_138 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@73305.4 package.scala 96:25:@73306.4]
  assign _T_156 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@73323.4 package.scala 96:25:@73324.4]
  assign _T_160 = _T_156 == 1'h0; // @[Controllers.scala 169:67:@73326.4]
  assign _T_161 = _T_160 & io_enable; // @[Controllers.scala 169:86:@73327.4]
  assign _T_174 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@73341.4]
  assign _T_176 = _T_174 & _T_105; // @[Controllers.scala 213:90:@73343.4]
  assign _T_178 = ~ done_0_io_output; // @[Controllers.scala 213:132:@73345.4]
  assign _T_187 = done_0_io_output & _T_186; // @[package.scala 100:41:@73353.4]
  assign io_done = RetimeWrapper_4_io_out; // @[Controllers.scala 245:13:@73379.4]
  assign io_enableOut_0 = _T_176 & _T_178; // @[Controllers.scala 213:55:@73349.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@73340.4]
  assign active_0_clock = clock; // @[:@73236.4]
  assign active_0_reset = reset; // @[:@73237.4]
  assign active_0_io_input_set = _T_115 & _T_118; // @[Controllers.scala 165:32:@73281.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@73285.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@73243.4]
  assign done_0_clock = clock; // @[:@73239.4]
  assign done_0_reset = reset; // @[:@73240.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_161; // @[Controllers.scala 169:30:@73331.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@73253.4 Controllers.scala 170:32:@73338.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@73244.4]
  assign iterDone_0_clock = clock; // @[:@73256.4]
  assign iterDone_0_reset = reset; // @[:@73257.4]
  assign iterDone_0_io_input_set = _T_131 & io_enable; // @[Controllers.scala 167:34:@73299.4]
  assign iterDone_0_io_input_reset = _T_138 | io_parentAck; // @[Controllers.scala 92:37:@73267.4 Controllers.scala 168:36:@73315.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@73258.4]
  assign RetimeWrapper_clock = clock; // @[:@73287.4]
  assign RetimeWrapper_reset = reset; // @[:@73288.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@73290.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@73289.4]
  assign RetimeWrapper_1_clock = clock; // @[:@73301.4]
  assign RetimeWrapper_1_reset = reset; // @[:@73302.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@73304.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@73303.4]
  assign RetimeWrapper_2_clock = clock; // @[:@73319.4]
  assign RetimeWrapper_2_reset = reset; // @[:@73320.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@73322.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@73321.4]
  assign RetimeWrapper_3_clock = clock; // @[:@73356.4]
  assign RetimeWrapper_3_reset = reset; // @[:@73357.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@73359.4]
  assign RetimeWrapper_3_io_in = _T_187 | io_parentAck; // @[package.scala 94:16:@73358.4]
  assign RetimeWrapper_4_clock = clock; // @[:@73373.4]
  assign RetimeWrapper_4_reset = reset; // @[:@73374.4]
  assign RetimeWrapper_4_io_flow = io_enable; // @[package.scala 95:18:@73376.4]
  assign RetimeWrapper_4_io_in = done_0_io_output & _T_200; // @[package.scala 94:16:@73375.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_200 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= _T_110;
    end
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_110;
    end
  end
endmodule
module x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1( // @[:@76452.2]
  input         clock, // @[:@76453.4]
  input         reset, // @[:@76454.4]
  output [31:0] io_in_x677_reg_wPort_0_data_0, // @[:@76455.4]
  output        io_in_x677_reg_wPort_0_reset, // @[:@76455.4]
  output        io_in_x677_reg_wPort_0_en_0, // @[:@76455.4]
  output        io_in_x677_reg_reset, // @[:@76455.4]
  output [31:0] io_in_x678_reg_wPort_0_data_0, // @[:@76455.4]
  output        io_in_x678_reg_wPort_0_reset, // @[:@76455.4]
  output        io_in_x678_reg_wPort_0_en_0, // @[:@76455.4]
  output        io_in_x678_reg_reset, // @[:@76455.4]
  input         io_in_x669_ready, // @[:@76455.4]
  output        io_in_x669_valid, // @[:@76455.4]
  output [63:0] io_in_x669_bits_addr, // @[:@76455.4]
  output [31:0] io_in_x669_bits_size, // @[:@76455.4]
  input  [31:0] io_in_b674_number, // @[:@76455.4]
  input  [63:0] io_in_x470_out_host_number, // @[:@76455.4]
  output [31:0] io_in_x676_reg_wPort_0_data_0, // @[:@76455.4]
  output        io_in_x676_reg_wPort_0_reset, // @[:@76455.4]
  output        io_in_x676_reg_wPort_0_en_0, // @[:@76455.4]
  output        io_in_x676_reg_reset, // @[:@76455.4]
  output [63:0] io_in_instrctrs_21_cycs, // @[:@76455.4]
  output [63:0] io_in_instrctrs_21_iters, // @[:@76455.4]
  output [63:0] io_in_instrctrs_21_stalls, // @[:@76455.4]
  output [63:0] io_in_instrctrs_21_idles, // @[:@76455.4]
  input         io_sigsIn_done, // @[:@76455.4]
  input         io_sigsIn_backpressure, // @[:@76455.4]
  input         io_sigsIn_datapathEn, // @[:@76455.4]
  input         io_sigsIn_baseEn, // @[:@76455.4]
  input         io_sigsIn_break, // @[:@76455.4]
  input         io_rr // @[:@76455.4]
);
  wire  cycles_x698_inr_UnitPipe_clock; // @[sm_x698_inr_UnitPipe.scala 80:44:@76600.4]
  wire  cycles_x698_inr_UnitPipe_reset; // @[sm_x698_inr_UnitPipe.scala 80:44:@76600.4]
  wire  cycles_x698_inr_UnitPipe_io_enable; // @[sm_x698_inr_UnitPipe.scala 80:44:@76600.4]
  wire [63:0] cycles_x698_inr_UnitPipe_io_count; // @[sm_x698_inr_UnitPipe.scala 80:44:@76600.4]
  wire  iters_x698_inr_UnitPipe_clock; // @[sm_x698_inr_UnitPipe.scala 81:43:@76603.4]
  wire  iters_x698_inr_UnitPipe_reset; // @[sm_x698_inr_UnitPipe.scala 81:43:@76603.4]
  wire  iters_x698_inr_UnitPipe_io_enable; // @[sm_x698_inr_UnitPipe.scala 81:43:@76603.4]
  wire [63:0] iters_x698_inr_UnitPipe_io_count; // @[sm_x698_inr_UnitPipe.scala 81:43:@76603.4]
  wire  stalls_x698_inr_UnitPipe_clock; // @[sm_x698_inr_UnitPipe.scala 84:44:@76612.4]
  wire  stalls_x698_inr_UnitPipe_reset; // @[sm_x698_inr_UnitPipe.scala 84:44:@76612.4]
  wire  stalls_x698_inr_UnitPipe_io_enable; // @[sm_x698_inr_UnitPipe.scala 84:44:@76612.4]
  wire [63:0] stalls_x698_inr_UnitPipe_io_count; // @[sm_x698_inr_UnitPipe.scala 84:44:@76612.4]
  wire  idles_x698_inr_UnitPipe_clock; // @[sm_x698_inr_UnitPipe.scala 85:43:@76615.4]
  wire  idles_x698_inr_UnitPipe_reset; // @[sm_x698_inr_UnitPipe.scala 85:43:@76615.4]
  wire  idles_x698_inr_UnitPipe_io_enable; // @[sm_x698_inr_UnitPipe.scala 85:43:@76615.4]
  wire [63:0] idles_x698_inr_UnitPipe_io_count; // @[sm_x698_inr_UnitPipe.scala 85:43:@76615.4]
  wire  x753_sum_1_clock; // @[Math.scala 150:24:@76637.4]
  wire  x753_sum_1_reset; // @[Math.scala 150:24:@76637.4]
  wire [31:0] x753_sum_1_io_a; // @[Math.scala 150:24:@76637.4]
  wire [31:0] x753_sum_1_io_b; // @[Math.scala 150:24:@76637.4]
  wire  x753_sum_1_io_flow; // @[Math.scala 150:24:@76637.4]
  wire [31:0] x753_sum_1_io_result; // @[Math.scala 150:24:@76637.4]
  wire  x683_sub_1_clock; // @[Math.scala 191:24:@76674.4]
  wire  x683_sub_1_reset; // @[Math.scala 191:24:@76674.4]
  wire [31:0] x683_sub_1_io_a; // @[Math.scala 191:24:@76674.4]
  wire [31:0] x683_sub_1_io_b; // @[Math.scala 191:24:@76674.4]
  wire  x683_sub_1_io_flow; // @[Math.scala 191:24:@76674.4]
  wire [31:0] x683_sub_1_io_result; // @[Math.scala 191:24:@76674.4]
  wire  x684_sum_1_clock; // @[Math.scala 150:24:@76686.4]
  wire  x684_sum_1_reset; // @[Math.scala 150:24:@76686.4]
  wire [31:0] x684_sum_1_io_a; // @[Math.scala 150:24:@76686.4]
  wire [31:0] x684_sum_1_io_b; // @[Math.scala 150:24:@76686.4]
  wire  x684_sum_1_io_flow; // @[Math.scala 150:24:@76686.4]
  wire [31:0] x684_sum_1_io_result; // @[Math.scala 150:24:@76686.4]
  wire  x685_sum_1_clock; // @[Math.scala 150:24:@76698.4]
  wire  x685_sum_1_reset; // @[Math.scala 150:24:@76698.4]
  wire [31:0] x685_sum_1_io_a; // @[Math.scala 150:24:@76698.4]
  wire [31:0] x685_sum_1_io_b; // @[Math.scala 150:24:@76698.4]
  wire  x685_sum_1_io_flow; // @[Math.scala 150:24:@76698.4]
  wire [31:0] x685_sum_1_io_result; // @[Math.scala 150:24:@76698.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@76727.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@76727.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@76727.4]
  wire [35:0] RetimeWrapper_io_in; // @[package.scala 93:22:@76727.4]
  wire [35:0] RetimeWrapper_io_out; // @[package.scala 93:22:@76727.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@76739.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@76739.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@76739.4]
  wire [37:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@76739.4]
  wire [37:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@76739.4]
  wire [31:0] x689_1_io_b; // @[Math.scala 720:24:@76749.4]
  wire [63:0] x689_1_io_result; // @[Math.scala 720:24:@76749.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@76759.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@76759.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@76759.4]
  wire [63:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@76759.4]
  wire [63:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@76759.4]
  wire  x691_sum_1_clock; // @[Math.scala 150:24:@76768.4]
  wire  x691_sum_1_reset; // @[Math.scala 150:24:@76768.4]
  wire [63:0] x691_sum_1_io_a; // @[Math.scala 150:24:@76768.4]
  wire [63:0] x691_sum_1_io_b; // @[Math.scala 150:24:@76768.4]
  wire  x691_sum_1_io_flow; // @[Math.scala 150:24:@76768.4]
  wire [63:0] x691_sum_1_io_result; // @[Math.scala 150:24:@76768.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@76779.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@76779.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@76779.4]
  wire [63:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@76779.4]
  wire [63:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@76779.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@76793.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@76793.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@76793.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@76793.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@76793.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@76803.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@76803.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@76803.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@76803.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@76803.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@76822.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@76822.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@76822.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@76822.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@76822.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@76842.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@76842.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@76842.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@76842.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@76842.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@76862.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@76862.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@76862.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@76862.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@76862.4]
  wire  _T_512; // @[package.scala 100:49:@76607.4]
  reg  _T_515; // @[package.scala 48:56:@76608.4]
  reg [31:0] _RAND_0;
  wire  _T_517; // @[sm_x698_inr_UnitPipe.scala 86:64:@76618.4]
  wire [32:0] _GEN_0; // @[Math.scala 461:32:@76633.4]
  wire [32:0] _T_527; // @[Math.scala 461:32:@76633.4]
  wire [31:0] x753_sum_number; // @[Math.scala 154:22:@76643.4 Math.scala 155:14:@76644.4]
  wire  _T_533; // @[FixedPoint.scala 50:25:@76648.4]
  wire [3:0] _T_537; // @[Bitwise.scala 72:12:@76650.4]
  wire [27:0] _T_538; // @[FixedPoint.scala 18:52:@76651.4]
  wire  _T_544; // @[Math.scala 451:55:@76653.4]
  wire [3:0] _T_545; // @[FixedPoint.scala 18:52:@76654.4]
  wire  _T_551; // @[Math.scala 451:110:@76656.4]
  wire  _T_552; // @[Math.scala 451:94:@76657.4]
  wire [31:0] _T_554; // @[Cat.scala 30:58:@76659.4]
  wire [31:0] x680_1_number; // @[Math.scala 454:20:@76660.4]
  wire [35:0] _GEN_1; // @[Math.scala 461:32:@76665.4]
  wire [35:0] _T_559; // @[Math.scala 461:32:@76665.4]
  wire [37:0] _GEN_2; // @[Math.scala 461:32:@76670.4]
  wire [37:0] _T_562; // @[Math.scala 461:32:@76670.4]
  wire [31:0] x685_sum_number; // @[Math.scala 154:22:@76704.4 Math.scala 155:14:@76705.4]
  wire  _T_582; // @[FixedPoint.scala 50:25:@76709.4]
  wire [3:0] _T_586; // @[Bitwise.scala 72:12:@76711.4]
  wire [27:0] _T_587; // @[FixedPoint.scala 18:52:@76712.4]
  wire  _T_593; // @[Math.scala 451:55:@76714.4]
  wire [3:0] _T_594; // @[FixedPoint.scala 18:52:@76715.4]
  wire  _T_600; // @[Math.scala 451:110:@76717.4]
  wire  _T_601; // @[Math.scala 451:94:@76718.4]
  wire [31:0] _T_603; // @[Cat.scala 30:58:@76720.4]
  wire [31:0] x686_1_number; // @[Math.scala 454:20:@76721.4]
  wire [35:0] _GEN_3; // @[Math.scala 461:32:@76726.4]
  wire [37:0] _GEN_4; // @[Math.scala 461:32:@76738.4]
  wire [37:0] _T_615; // @[package.scala 96:25:@76744.4 package.scala 96:25:@76745.4]
  wire [31:0] x755_1_number; // @[Math.scala 459:22:@76737.4 Math.scala 461:14:@76746.4]
  wire [63:0] x802_x691_sum_D1_number; // @[package.scala 96:25:@76784.4 package.scala 96:25:@76785.4]
  wire [96:0] x692_tuple; // @[Cat.scala 30:58:@76789.4]
  wire  _T_645; // @[package.scala 96:25:@76808.4 package.scala 96:25:@76809.4]
  wire  _T_647; // @[implicits.scala 56:10:@76810.4]
  wire  x803_x693_D4; // @[package.scala 96:25:@76798.4 package.scala 96:25:@76799.4]
  wire  _T_648; // @[sm_x698_inr_UnitPipe.scala 127:121:@76811.4]
  wire  _T_652; // @[sm_x698_inr_UnitPipe.scala 134:116:@76818.4]
  wire  _T_658; // @[package.scala 96:25:@76827.4 package.scala 96:25:@76828.4]
  wire  _T_660; // @[implicits.scala 56:10:@76829.4]
  wire  _T_661; // @[sm_x698_inr_UnitPipe.scala 134:133:@76830.4]
  wire  _T_663; // @[sm_x698_inr_UnitPipe.scala 134:230:@76832.4]
  wire  _T_673; // @[package.scala 96:25:@76847.4 package.scala 96:25:@76848.4]
  wire  _T_675; // @[implicits.scala 56:10:@76849.4]
  wire  _T_676; // @[sm_x698_inr_UnitPipe.scala 139:133:@76850.4]
  wire  _T_678; // @[sm_x698_inr_UnitPipe.scala 139:230:@76852.4]
  wire  _T_688; // @[package.scala 96:25:@76867.4 package.scala 96:25:@76868.4]
  wire  _T_690; // @[implicits.scala 56:10:@76869.4]
  wire  _T_691; // @[sm_x698_inr_UnitPipe.scala 144:133:@76870.4]
  wire  _T_693; // @[sm_x698_inr_UnitPipe.scala 144:230:@76872.4]
  wire [35:0] _T_610; // @[package.scala 96:25:@76732.4 package.scala 96:25:@76733.4]
  InstrumentationCounter cycles_x698_inr_UnitPipe ( // @[sm_x698_inr_UnitPipe.scala 80:44:@76600.4]
    .clock(cycles_x698_inr_UnitPipe_clock),
    .reset(cycles_x698_inr_UnitPipe_reset),
    .io_enable(cycles_x698_inr_UnitPipe_io_enable),
    .io_count(cycles_x698_inr_UnitPipe_io_count)
  );
  InstrumentationCounter iters_x698_inr_UnitPipe ( // @[sm_x698_inr_UnitPipe.scala 81:43:@76603.4]
    .clock(iters_x698_inr_UnitPipe_clock),
    .reset(iters_x698_inr_UnitPipe_reset),
    .io_enable(iters_x698_inr_UnitPipe_io_enable),
    .io_count(iters_x698_inr_UnitPipe_io_count)
  );
  InstrumentationCounter stalls_x698_inr_UnitPipe ( // @[sm_x698_inr_UnitPipe.scala 84:44:@76612.4]
    .clock(stalls_x698_inr_UnitPipe_clock),
    .reset(stalls_x698_inr_UnitPipe_reset),
    .io_enable(stalls_x698_inr_UnitPipe_io_enable),
    .io_count(stalls_x698_inr_UnitPipe_io_count)
  );
  InstrumentationCounter idles_x698_inr_UnitPipe ( // @[sm_x698_inr_UnitPipe.scala 85:43:@76615.4]
    .clock(idles_x698_inr_UnitPipe_clock),
    .reset(idles_x698_inr_UnitPipe_reset),
    .io_enable(idles_x698_inr_UnitPipe_io_enable),
    .io_count(idles_x698_inr_UnitPipe_io_count)
  );
  x739_sum x753_sum_1 ( // @[Math.scala 150:24:@76637.4]
    .clock(x753_sum_1_clock),
    .reset(x753_sum_1_reset),
    .io_a(x753_sum_1_io_a),
    .io_b(x753_sum_1_io_b),
    .io_flow(x753_sum_1_io_flow),
    .io_result(x753_sum_1_io_result)
  );
  x485_sub x683_sub_1 ( // @[Math.scala 191:24:@76674.4]
    .clock(x683_sub_1_clock),
    .reset(x683_sub_1_reset),
    .io_a(x683_sub_1_io_a),
    .io_b(x683_sub_1_io_b),
    .io_flow(x683_sub_1_io_flow),
    .io_result(x683_sub_1_io_result)
  );
  x739_sum x684_sum_1 ( // @[Math.scala 150:24:@76686.4]
    .clock(x684_sum_1_clock),
    .reset(x684_sum_1_reset),
    .io_a(x684_sum_1_io_a),
    .io_b(x684_sum_1_io_b),
    .io_flow(x684_sum_1_io_flow),
    .io_result(x684_sum_1_io_result)
  );
  x739_sum x685_sum_1 ( // @[Math.scala 150:24:@76698.4]
    .clock(x685_sum_1_clock),
    .reset(x685_sum_1_reset),
    .io_a(x685_sum_1_io_a),
    .io_b(x685_sum_1_io_b),
    .io_flow(x685_sum_1_io_flow),
    .io_result(x685_sum_1_io_result)
  );
  RetimeWrapper_36 RetimeWrapper ( // @[package.scala 93:22:@76727.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_37 RetimeWrapper_1 ( // @[package.scala 93:22:@76739.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x491 x689_1 ( // @[Math.scala 720:24:@76749.4]
    .io_b(x689_1_io_b),
    .io_result(x689_1_io_result)
  );
  RetimeWrapper_38 RetimeWrapper_2 ( // @[package.scala 93:22:@76759.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x493_sum x691_sum_1 ( // @[Math.scala 150:24:@76768.4]
    .clock(x691_sum_1_clock),
    .reset(x691_sum_1_reset),
    .io_a(x691_sum_1_io_a),
    .io_b(x691_sum_1_io_b),
    .io_flow(x691_sum_1_io_flow),
    .io_result(x691_sum_1_io_result)
  );
  RetimeWrapper_38 RetimeWrapper_3 ( // @[package.scala 93:22:@76779.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@76793.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_5 ( // @[package.scala 93:22:@76803.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@76822.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_59 RetimeWrapper_7 ( // @[package.scala 93:22:@76842.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_8 ( // @[package.scala 93:22:@76862.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  assign _T_512 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@76607.4]
  assign _T_517 = ~ io_in_x669_ready; // @[sm_x698_inr_UnitPipe.scala 86:64:@76618.4]
  assign _GEN_0 = {{1'd0}, io_in_b674_number}; // @[Math.scala 461:32:@76633.4]
  assign _T_527 = _GEN_0 << 1; // @[Math.scala 461:32:@76633.4]
  assign x753_sum_number = x753_sum_1_io_result; // @[Math.scala 154:22:@76643.4 Math.scala 155:14:@76644.4]
  assign _T_533 = x753_sum_number[31]; // @[FixedPoint.scala 50:25:@76648.4]
  assign _T_537 = _T_533 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@76650.4]
  assign _T_538 = x753_sum_number[31:4]; // @[FixedPoint.scala 18:52:@76651.4]
  assign _T_544 = _T_538 == 28'hfffffff; // @[Math.scala 451:55:@76653.4]
  assign _T_545 = x753_sum_number[3:0]; // @[FixedPoint.scala 18:52:@76654.4]
  assign _T_551 = _T_545 != 4'h0; // @[Math.scala 451:110:@76656.4]
  assign _T_552 = _T_544 & _T_551; // @[Math.scala 451:94:@76657.4]
  assign _T_554 = {_T_537,_T_538}; // @[Cat.scala 30:58:@76659.4]
  assign x680_1_number = _T_552 ? 32'h0 : _T_554; // @[Math.scala 454:20:@76660.4]
  assign _GEN_1 = {{4'd0}, x680_1_number}; // @[Math.scala 461:32:@76665.4]
  assign _T_559 = _GEN_1 << 4; // @[Math.scala 461:32:@76665.4]
  assign _GEN_2 = {{6'd0}, x680_1_number}; // @[Math.scala 461:32:@76670.4]
  assign _T_562 = _GEN_2 << 6; // @[Math.scala 461:32:@76670.4]
  assign x685_sum_number = x685_sum_1_io_result; // @[Math.scala 154:22:@76704.4 Math.scala 155:14:@76705.4]
  assign _T_582 = x685_sum_number[31]; // @[FixedPoint.scala 50:25:@76709.4]
  assign _T_586 = _T_582 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@76711.4]
  assign _T_587 = x685_sum_number[31:4]; // @[FixedPoint.scala 18:52:@76712.4]
  assign _T_593 = _T_587 == 28'hfffffff; // @[Math.scala 451:55:@76714.4]
  assign _T_594 = x685_sum_number[3:0]; // @[FixedPoint.scala 18:52:@76715.4]
  assign _T_600 = _T_594 != 4'h0; // @[Math.scala 451:110:@76717.4]
  assign _T_601 = _T_593 & _T_600; // @[Math.scala 451:94:@76718.4]
  assign _T_603 = {_T_586,_T_587}; // @[Cat.scala 30:58:@76720.4]
  assign x686_1_number = _T_601 ? 32'h0 : _T_603; // @[Math.scala 454:20:@76721.4]
  assign _GEN_3 = {{4'd0}, x686_1_number}; // @[Math.scala 461:32:@76726.4]
  assign _GEN_4 = {{6'd0}, x686_1_number}; // @[Math.scala 461:32:@76738.4]
  assign _T_615 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@76744.4 package.scala 96:25:@76745.4]
  assign x755_1_number = _T_615[31:0]; // @[Math.scala 459:22:@76737.4 Math.scala 461:14:@76746.4]
  assign x802_x691_sum_D1_number = RetimeWrapper_3_io_out; // @[package.scala 96:25:@76784.4 package.scala 96:25:@76785.4]
  assign x692_tuple = {1'h0,x755_1_number,x802_x691_sum_D1_number}; // @[Cat.scala 30:58:@76789.4]
  assign _T_645 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@76808.4 package.scala 96:25:@76809.4]
  assign _T_647 = io_rr ? _T_645 : 1'h0; // @[implicits.scala 56:10:@76810.4]
  assign x803_x693_D4 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@76798.4 package.scala 96:25:@76799.4]
  assign _T_648 = _T_647 & x803_x693_D4; // @[sm_x698_inr_UnitPipe.scala 127:121:@76811.4]
  assign _T_652 = ~ io_sigsIn_break; // @[sm_x698_inr_UnitPipe.scala 134:116:@76818.4]
  assign _T_658 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@76827.4 package.scala 96:25:@76828.4]
  assign _T_660 = io_rr ? _T_658 : 1'h0; // @[implicits.scala 56:10:@76829.4]
  assign _T_661 = _T_652 & _T_660; // @[sm_x698_inr_UnitPipe.scala 134:133:@76830.4]
  assign _T_663 = _T_661 & _T_652; // @[sm_x698_inr_UnitPipe.scala 134:230:@76832.4]
  assign _T_673 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@76847.4 package.scala 96:25:@76848.4]
  assign _T_675 = io_rr ? _T_673 : 1'h0; // @[implicits.scala 56:10:@76849.4]
  assign _T_676 = _T_652 & _T_675; // @[sm_x698_inr_UnitPipe.scala 139:133:@76850.4]
  assign _T_678 = _T_676 & _T_652; // @[sm_x698_inr_UnitPipe.scala 139:230:@76852.4]
  assign _T_688 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@76867.4 package.scala 96:25:@76868.4]
  assign _T_690 = io_rr ? _T_688 : 1'h0; // @[implicits.scala 56:10:@76869.4]
  assign _T_691 = _T_652 & _T_690; // @[sm_x698_inr_UnitPipe.scala 144:133:@76870.4]
  assign _T_693 = _T_691 & _T_652; // @[sm_x698_inr_UnitPipe.scala 144:230:@76872.4]
  assign _T_610 = RetimeWrapper_io_out; // @[package.scala 96:25:@76732.4 package.scala 96:25:@76733.4]
  assign io_in_x677_reg_wPort_0_data_0 = x684_sum_1_io_result; // @[MemInterfaceType.scala 90:56:@76855.4]
  assign io_in_x677_reg_wPort_0_reset = io_in_x677_reg_reset; // @[MemInterfaceType.scala 91:23:@76856.4]
  assign io_in_x677_reg_wPort_0_en_0 = _T_678 & io_sigsIn_backpressure; // @[MemInterfaceType.scala 93:57:@76857.4]
  assign io_in_x677_reg_reset = 1'h0;
  assign io_in_x678_reg_wPort_0_data_0 = _T_610[31:0]; // @[MemInterfaceType.scala 90:56:@76875.4]
  assign io_in_x678_reg_wPort_0_reset = io_in_x678_reg_reset; // @[MemInterfaceType.scala 91:23:@76876.4]
  assign io_in_x678_reg_wPort_0_en_0 = _T_693 & io_sigsIn_backpressure; // @[MemInterfaceType.scala 93:57:@76877.4]
  assign io_in_x678_reg_reset = 1'h0;
  assign io_in_x669_valid = _T_648 & io_sigsIn_backpressure; // @[sm_x698_inr_UnitPipe.scala 127:18:@76813.4]
  assign io_in_x669_bits_addr = x692_tuple[63:0]; // @[sm_x698_inr_UnitPipe.scala 128:22:@76815.4]
  assign io_in_x669_bits_size = x692_tuple[95:64]; // @[sm_x698_inr_UnitPipe.scala 129:22:@76817.4]
  assign io_in_x676_reg_wPort_0_data_0 = x683_sub_1_io_result; // @[MemInterfaceType.scala 90:56:@76835.4]
  assign io_in_x676_reg_wPort_0_reset = io_in_x676_reg_reset; // @[MemInterfaceType.scala 91:23:@76836.4]
  assign io_in_x676_reg_wPort_0_en_0 = _T_663 & io_sigsIn_backpressure; // @[MemInterfaceType.scala 93:57:@76837.4]
  assign io_in_x676_reg_reset = 1'h0;
  assign io_in_instrctrs_21_cycs = cycles_x698_inr_UnitPipe_io_count; // @[Ledger.scala 293:21:@76625.4]
  assign io_in_instrctrs_21_iters = iters_x698_inr_UnitPipe_io_count; // @[Ledger.scala 294:22:@76626.4]
  assign io_in_instrctrs_21_stalls = stalls_x698_inr_UnitPipe_io_count; // @[Ledger.scala 295:23:@76627.4]
  assign io_in_instrctrs_21_idles = idles_x698_inr_UnitPipe_io_count; // @[Ledger.scala 296:22:@76628.4]
  assign cycles_x698_inr_UnitPipe_clock = clock; // @[:@76601.4]
  assign cycles_x698_inr_UnitPipe_reset = reset; // @[:@76602.4]
  assign cycles_x698_inr_UnitPipe_io_enable = io_sigsIn_baseEn; // @[sm_x698_inr_UnitPipe.scala 82:42:@76606.4]
  assign iters_x698_inr_UnitPipe_clock = clock; // @[:@76604.4]
  assign iters_x698_inr_UnitPipe_reset = reset; // @[:@76605.4]
  assign iters_x698_inr_UnitPipe_io_enable = io_sigsIn_done & _T_515; // @[sm_x698_inr_UnitPipe.scala 83:41:@76611.4]
  assign stalls_x698_inr_UnitPipe_clock = clock; // @[:@76613.4]
  assign stalls_x698_inr_UnitPipe_reset = reset; // @[:@76614.4]
  assign stalls_x698_inr_UnitPipe_io_enable = io_sigsIn_baseEn & _T_517; // @[sm_x698_inr_UnitPipe.scala 86:42:@76620.4]
  assign idles_x698_inr_UnitPipe_clock = clock; // @[:@76616.4]
  assign idles_x698_inr_UnitPipe_reset = reset; // @[:@76617.4]
  assign idles_x698_inr_UnitPipe_io_enable = 1'h0; // @[sm_x698_inr_UnitPipe.scala 87:41:@76624.4]
  assign x753_sum_1_clock = clock; // @[:@76638.4]
  assign x753_sum_1_reset = reset; // @[:@76639.4]
  assign x753_sum_1_io_a = _T_527[31:0]; // @[Math.scala 151:17:@76640.4]
  assign x753_sum_1_io_b = io_in_b674_number; // @[Math.scala 152:17:@76641.4]
  assign x753_sum_1_io_flow = io_in_x669_ready; // @[Math.scala 153:20:@76642.4]
  assign x683_sub_1_clock = clock; // @[:@76675.4]
  assign x683_sub_1_reset = reset; // @[:@76676.4]
  assign x683_sub_1_io_a = x753_sum_1_io_result; // @[Math.scala 192:17:@76677.4]
  assign x683_sub_1_io_b = _T_559[31:0]; // @[Math.scala 193:17:@76678.4]
  assign x683_sub_1_io_flow = io_in_x669_ready; // @[Math.scala 194:20:@76679.4]
  assign x684_sum_1_clock = clock; // @[:@76687.4]
  assign x684_sum_1_reset = reset; // @[:@76688.4]
  assign x684_sum_1_io_a = x683_sub_1_io_result; // @[Math.scala 151:17:@76689.4]
  assign x684_sum_1_io_b = 32'h3; // @[Math.scala 152:17:@76690.4]
  assign x684_sum_1_io_flow = io_in_x669_ready; // @[Math.scala 153:20:@76691.4]
  assign x685_sum_1_clock = clock; // @[:@76699.4]
  assign x685_sum_1_reset = reset; // @[:@76700.4]
  assign x685_sum_1_io_a = x683_sub_1_io_result; // @[Math.scala 151:17:@76701.4]
  assign x685_sum_1_io_b = 32'h12; // @[Math.scala 152:17:@76702.4]
  assign x685_sum_1_io_flow = io_in_x669_ready; // @[Math.scala 153:20:@76703.4]
  assign RetimeWrapper_clock = clock; // @[:@76728.4]
  assign RetimeWrapper_reset = reset; // @[:@76729.4]
  assign RetimeWrapper_io_flow = io_in_x669_ready; // @[package.scala 95:18:@76731.4]
  assign RetimeWrapper_io_in = _GEN_3 << 4; // @[package.scala 94:16:@76730.4]
  assign RetimeWrapper_1_clock = clock; // @[:@76740.4]
  assign RetimeWrapper_1_reset = reset; // @[:@76741.4]
  assign RetimeWrapper_1_io_flow = io_in_x669_ready; // @[package.scala 95:18:@76743.4]
  assign RetimeWrapper_1_io_in = _GEN_4 << 6; // @[package.scala 94:16:@76742.4]
  assign x689_1_io_b = _T_562[31:0]; // @[Math.scala 721:17:@76752.4]
  assign RetimeWrapper_2_clock = clock; // @[:@76760.4]
  assign RetimeWrapper_2_reset = reset; // @[:@76761.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@76763.4]
  assign RetimeWrapper_2_io_in = io_in_x470_out_host_number; // @[package.scala 94:16:@76762.4]
  assign x691_sum_1_clock = clock; // @[:@76769.4]
  assign x691_sum_1_reset = reset; // @[:@76770.4]
  assign x691_sum_1_io_a = x689_1_io_result; // @[Math.scala 151:17:@76771.4]
  assign x691_sum_1_io_b = RetimeWrapper_2_io_out; // @[Math.scala 152:17:@76772.4]
  assign x691_sum_1_io_flow = io_in_x669_ready; // @[Math.scala 153:20:@76773.4]
  assign RetimeWrapper_3_clock = clock; // @[:@76780.4]
  assign RetimeWrapper_3_reset = reset; // @[:@76781.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@76783.4]
  assign RetimeWrapper_3_io_in = x691_sum_1_io_result; // @[package.scala 94:16:@76782.4]
  assign RetimeWrapper_4_clock = clock; // @[:@76794.4]
  assign RetimeWrapper_4_reset = reset; // @[:@76795.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@76797.4]
  assign RetimeWrapper_4_io_in = 1'h1; // @[package.scala 94:16:@76796.4]
  assign RetimeWrapper_5_clock = clock; // @[:@76804.4]
  assign RetimeWrapper_5_reset = reset; // @[:@76805.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@76807.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@76806.4]
  assign RetimeWrapper_6_clock = clock; // @[:@76823.4]
  assign RetimeWrapper_6_reset = reset; // @[:@76824.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@76826.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@76825.4]
  assign RetimeWrapper_7_clock = clock; // @[:@76843.4]
  assign RetimeWrapper_7_reset = reset; // @[:@76844.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@76846.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@76845.4]
  assign RetimeWrapper_8_clock = clock; // @[:@76863.4]
  assign RetimeWrapper_8_reset = reset; // @[:@76864.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@76866.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@76865.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_515 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_515 <= 1'h0;
    end else begin
      _T_515 <= _T_512;
    end
  end
endmodule
module x717_inr_Foreach_kernelx717_inr_Foreach_concrete1( // @[:@78327.2]
  input         clock, // @[:@78328.4]
  input         reset, // @[:@78329.4]
  input  [31:0] io_in_x677_reg_rPort_0_output_0, // @[:@78330.4]
  input         io_in_x670_ready, // @[:@78330.4]
  output        io_in_x670_valid, // @[:@78330.4]
  output [31:0] io_in_x670_bits_wdata_0, // @[:@78330.4]
  output        io_in_x670_bits_wstrb, // @[:@78330.4]
  input  [31:0] io_in_b674_number, // @[:@78330.4]
  output [8:0]  io_in_x539_out_sram_0_rPort_0_ofs_0, // @[:@78330.4]
  output        io_in_x539_out_sram_0_rPort_0_en_0, // @[:@78330.4]
  output        io_in_x539_out_sram_0_rPort_0_backpressure, // @[:@78330.4]
  input  [31:0] io_in_x539_out_sram_0_rPort_0_output_0, // @[:@78330.4]
  input  [31:0] io_in_x676_reg_rPort_0_output_0, // @[:@78330.4]
  output [63:0] io_in_instrctrs_22_cycs, // @[:@78330.4]
  output [63:0] io_in_instrctrs_22_iters, // @[:@78330.4]
  output [63:0] io_in_instrctrs_22_stalls, // @[:@78330.4]
  output [63:0] io_in_instrctrs_22_idles, // @[:@78330.4]
  input         io_sigsIn_done, // @[:@78330.4]
  input         io_sigsIn_backpressure, // @[:@78330.4]
  input         io_sigsIn_datapathEn, // @[:@78330.4]
  input         io_sigsIn_baseEn, // @[:@78330.4]
  input         io_sigsIn_break, // @[:@78330.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@78330.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@78330.4]
  input         io_rr // @[:@78330.4]
);
  wire  cycles_x717_inr_Foreach_clock; // @[sm_x717_inr_Foreach.scala 76:43:@78475.4]
  wire  cycles_x717_inr_Foreach_reset; // @[sm_x717_inr_Foreach.scala 76:43:@78475.4]
  wire  cycles_x717_inr_Foreach_io_enable; // @[sm_x717_inr_Foreach.scala 76:43:@78475.4]
  wire [63:0] cycles_x717_inr_Foreach_io_count; // @[sm_x717_inr_Foreach.scala 76:43:@78475.4]
  wire  iters_x717_inr_Foreach_clock; // @[sm_x717_inr_Foreach.scala 77:42:@78478.4]
  wire  iters_x717_inr_Foreach_reset; // @[sm_x717_inr_Foreach.scala 77:42:@78478.4]
  wire  iters_x717_inr_Foreach_io_enable; // @[sm_x717_inr_Foreach.scala 77:42:@78478.4]
  wire [63:0] iters_x717_inr_Foreach_io_count; // @[sm_x717_inr_Foreach.scala 77:42:@78478.4]
  wire  stalls_x717_inr_Foreach_clock; // @[sm_x717_inr_Foreach.scala 80:43:@78487.4]
  wire  stalls_x717_inr_Foreach_reset; // @[sm_x717_inr_Foreach.scala 80:43:@78487.4]
  wire  stalls_x717_inr_Foreach_io_enable; // @[sm_x717_inr_Foreach.scala 80:43:@78487.4]
  wire [63:0] stalls_x717_inr_Foreach_io_count; // @[sm_x717_inr_Foreach.scala 80:43:@78487.4]
  wire  idles_x717_inr_Foreach_clock; // @[sm_x717_inr_Foreach.scala 81:42:@78490.4]
  wire  idles_x717_inr_Foreach_reset; // @[sm_x717_inr_Foreach.scala 81:42:@78490.4]
  wire  idles_x717_inr_Foreach_io_enable; // @[sm_x717_inr_Foreach.scala 81:42:@78490.4]
  wire [63:0] idles_x717_inr_Foreach_io_count; // @[sm_x717_inr_Foreach.scala 81:42:@78490.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@78508.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@78508.4]
  wire  x709_sub_1_clock; // @[Math.scala 191:24:@78561.4]
  wire  x709_sub_1_reset; // @[Math.scala 191:24:@78561.4]
  wire [31:0] x709_sub_1_io_a; // @[Math.scala 191:24:@78561.4]
  wire [31:0] x709_sub_1_io_b; // @[Math.scala 191:24:@78561.4]
  wire  x709_sub_1_io_flow; // @[Math.scala 191:24:@78561.4]
  wire [31:0] x709_sub_1_io_result; // @[Math.scala 191:24:@78561.4]
  wire  x757_sum_1_clock; // @[Math.scala 150:24:@78576.4]
  wire  x757_sum_1_reset; // @[Math.scala 150:24:@78576.4]
  wire [31:0] x757_sum_1_io_a; // @[Math.scala 150:24:@78576.4]
  wire [31:0] x757_sum_1_io_b; // @[Math.scala 150:24:@78576.4]
  wire  x757_sum_1_io_flow; // @[Math.scala 150:24:@78576.4]
  wire [31:0] x757_sum_1_io_result; // @[Math.scala 150:24:@78576.4]
  wire  x712_sum_1_clock; // @[Math.scala 150:24:@78586.4]
  wire  x712_sum_1_reset; // @[Math.scala 150:24:@78586.4]
  wire [31:0] x712_sum_1_io_a; // @[Math.scala 150:24:@78586.4]
  wire [31:0] x712_sum_1_io_b; // @[Math.scala 150:24:@78586.4]
  wire  x712_sum_1_io_flow; // @[Math.scala 150:24:@78586.4]
  wire [31:0] x712_sum_1_io_result; // @[Math.scala 150:24:@78586.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@78597.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@78597.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@78597.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@78597.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@78597.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@78607.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@78607.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@78607.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@78607.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@78607.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@78619.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@78619.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@78619.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@78619.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@78619.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@78631.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@78631.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@78631.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@78631.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@78631.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@78652.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@78652.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@78652.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@78652.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@78652.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@78665.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@78665.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@78665.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@78665.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@78665.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@78675.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@78675.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@78675.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@78675.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@78675.4]
  wire  _T_518; // @[package.scala 100:49:@78482.4]
  reg  _T_521; // @[package.scala 48:56:@78483.4]
  reg [31:0] _RAND_0;
  wire  _T_523; // @[sm_x717_inr_Foreach.scala 82:63:@78493.4]
  wire  _T_542; // @[sm_x717_inr_Foreach.scala 91:119:@78520.4]
  wire [31:0] _T_554; // @[Math.scala 493:37:@78534.4]
  wire [31:0] b702_number; // @[Math.scala 723:22:@78513.4 Math.scala 724:14:@78514.4]
  wire [31:0] _T_555; // @[Math.scala 493:51:@78535.4]
  wire  x705; // @[Math.scala 493:44:@78536.4]
  wire [31:0] _T_574; // @[Math.scala 476:50:@78554.4]
  wire  x707; // @[Math.scala 476:44:@78555.4]
  wire [32:0] _GEN_0; // @[Math.scala 461:32:@78572.4]
  wire [32:0] _T_583; // @[Math.scala 461:32:@78572.4]
  wire  _T_613; // @[package.scala 96:25:@78624.4 package.scala 96:25:@78625.4]
  wire  _T_615; // @[implicits.scala 56:10:@78626.4]
  wire  _T_617; // @[sm_x717_inr_Foreach.scala 123:111:@78628.4]
  wire  _T_622; // @[package.scala 96:25:@78636.4 package.scala 96:25:@78637.4]
  wire  _T_624; // @[implicits.scala 56:10:@78638.4]
  wire  _T_625; // @[sm_x717_inr_Foreach.scala 123:131:@78639.4]
  wire  x805_x708_D2; // @[package.scala 96:25:@78612.4 package.scala 96:25:@78613.4]
  wire  _T_626; // @[sm_x717_inr_Foreach.scala 123:228:@78640.4]
  wire  x804_b703_D2; // @[package.scala 96:25:@78602.4 package.scala 96:25:@78603.4]
  wire  x806_x708_D4; // @[package.scala 96:25:@78657.4 package.scala 96:25:@78658.4]
  wire [32:0] x715_tuple; // @[Cat.scala 30:58:@78661.4]
  wire  _T_645; // @[package.scala 96:25:@78680.4 package.scala 96:25:@78681.4]
  wire  _T_647; // @[implicits.scala 56:10:@78682.4]
  wire  x807_b703_D4; // @[package.scala 96:25:@78670.4 package.scala 96:25:@78671.4]
  wire  _T_648; // @[sm_x717_inr_Foreach.scala 134:121:@78683.4]
  wire [31:0] x712_sum_number; // @[Math.scala 154:22:@78592.4 Math.scala 155:14:@78593.4]
  InstrumentationCounter cycles_x717_inr_Foreach ( // @[sm_x717_inr_Foreach.scala 76:43:@78475.4]
    .clock(cycles_x717_inr_Foreach_clock),
    .reset(cycles_x717_inr_Foreach_reset),
    .io_enable(cycles_x717_inr_Foreach_io_enable),
    .io_count(cycles_x717_inr_Foreach_io_count)
  );
  InstrumentationCounter iters_x717_inr_Foreach ( // @[sm_x717_inr_Foreach.scala 77:42:@78478.4]
    .clock(iters_x717_inr_Foreach_clock),
    .reset(iters_x717_inr_Foreach_reset),
    .io_enable(iters_x717_inr_Foreach_io_enable),
    .io_count(iters_x717_inr_Foreach_io_count)
  );
  InstrumentationCounter stalls_x717_inr_Foreach ( // @[sm_x717_inr_Foreach.scala 80:43:@78487.4]
    .clock(stalls_x717_inr_Foreach_clock),
    .reset(stalls_x717_inr_Foreach_reset),
    .io_enable(stalls_x717_inr_Foreach_io_enable),
    .io_count(stalls_x717_inr_Foreach_io_count)
  );
  InstrumentationCounter idles_x717_inr_Foreach ( // @[sm_x717_inr_Foreach.scala 81:42:@78490.4]
    .clock(idles_x717_inr_Foreach_clock),
    .reset(idles_x717_inr_Foreach_reset),
    .io_enable(idles_x717_inr_Foreach_io_enable),
    .io_count(idles_x717_inr_Foreach_io_count)
  );
  _ _ ( // @[Math.scala 720:24:@78508.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x485_sub x709_sub_1 ( // @[Math.scala 191:24:@78561.4]
    .clock(x709_sub_1_clock),
    .reset(x709_sub_1_reset),
    .io_a(x709_sub_1_io_a),
    .io_b(x709_sub_1_io_b),
    .io_flow(x709_sub_1_io_flow),
    .io_result(x709_sub_1_io_result)
  );
  x739_sum x757_sum_1 ( // @[Math.scala 150:24:@78576.4]
    .clock(x757_sum_1_clock),
    .reset(x757_sum_1_reset),
    .io_a(x757_sum_1_io_a),
    .io_b(x757_sum_1_io_b),
    .io_flow(x757_sum_1_io_flow),
    .io_result(x757_sum_1_io_result)
  );
  x739_sum x712_sum_1 ( // @[Math.scala 150:24:@78586.4]
    .clock(x712_sum_1_clock),
    .reset(x712_sum_1_reset),
    .io_a(x712_sum_1_io_a),
    .io_b(x712_sum_1_io_b),
    .io_flow(x712_sum_1_io_flow),
    .io_result(x712_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@78597.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@78607.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@78619.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@78631.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@78652.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_5 ( // @[package.scala 93:22:@78665.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_6 ( // @[package.scala 93:22:@78675.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  assign _T_518 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@78482.4]
  assign _T_523 = ~ io_in_x670_ready; // @[sm_x717_inr_Foreach.scala 82:63:@78493.4]
  assign _T_542 = ~ io_sigsIn_break; // @[sm_x717_inr_Foreach.scala 91:119:@78520.4]
  assign _T_554 = $signed(io_in_x676_reg_rPort_0_output_0); // @[Math.scala 493:37:@78534.4]
  assign b702_number = __io_result; // @[Math.scala 723:22:@78513.4 Math.scala 724:14:@78514.4]
  assign _T_555 = $signed(b702_number); // @[Math.scala 493:51:@78535.4]
  assign x705 = $signed(_T_554) <= $signed(_T_555); // @[Math.scala 493:44:@78536.4]
  assign _T_574 = $signed(io_in_x677_reg_rPort_0_output_0); // @[Math.scala 476:50:@78554.4]
  assign x707 = $signed(_T_555) < $signed(_T_574); // @[Math.scala 476:44:@78555.4]
  assign _GEN_0 = {{1'd0}, io_in_b674_number}; // @[Math.scala 461:32:@78572.4]
  assign _T_583 = _GEN_0 << 1; // @[Math.scala 461:32:@78572.4]
  assign _T_613 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@78624.4 package.scala 96:25:@78625.4]
  assign _T_615 = io_rr ? _T_613 : 1'h0; // @[implicits.scala 56:10:@78626.4]
  assign _T_617 = _T_615 & _T_542; // @[sm_x717_inr_Foreach.scala 123:111:@78628.4]
  assign _T_622 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@78636.4 package.scala 96:25:@78637.4]
  assign _T_624 = io_rr ? _T_622 : 1'h0; // @[implicits.scala 56:10:@78638.4]
  assign _T_625 = _T_617 & _T_624; // @[sm_x717_inr_Foreach.scala 123:131:@78639.4]
  assign x805_x708_D2 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@78612.4 package.scala 96:25:@78613.4]
  assign _T_626 = _T_625 & x805_x708_D2; // @[sm_x717_inr_Foreach.scala 123:228:@78640.4]
  assign x804_b703_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@78602.4 package.scala 96:25:@78603.4]
  assign x806_x708_D4 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@78657.4 package.scala 96:25:@78658.4]
  assign x715_tuple = {x806_x708_D4,io_in_x539_out_sram_0_rPort_0_output_0}; // @[Cat.scala 30:58:@78661.4]
  assign _T_645 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@78680.4 package.scala 96:25:@78681.4]
  assign _T_647 = io_rr ? _T_645 : 1'h0; // @[implicits.scala 56:10:@78682.4]
  assign x807_b703_D4 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@78670.4 package.scala 96:25:@78671.4]
  assign _T_648 = _T_647 & x807_b703_D4; // @[sm_x717_inr_Foreach.scala 134:121:@78683.4]
  assign x712_sum_number = x712_sum_1_io_result; // @[Math.scala 154:22:@78592.4 Math.scala 155:14:@78593.4]
  assign io_in_x670_valid = _T_648 & io_sigsIn_backpressure; // @[sm_x717_inr_Foreach.scala 134:18:@78685.4]
  assign io_in_x670_bits_wdata_0 = x715_tuple[31:0]; // @[sm_x717_inr_Foreach.scala 135:26:@78687.4]
  assign io_in_x670_bits_wstrb = x715_tuple[32]; // @[sm_x717_inr_Foreach.scala 136:23:@78689.4]
  assign io_in_x539_out_sram_0_rPort_0_ofs_0 = x712_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@78644.4]
  assign io_in_x539_out_sram_0_rPort_0_en_0 = _T_626 & x804_b703_D2; // @[MemInterfaceType.scala 110:79:@78646.4]
  assign io_in_x539_out_sram_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@78645.4]
  assign io_in_instrctrs_22_cycs = cycles_x717_inr_Foreach_io_count; // @[Ledger.scala 293:21:@78500.4]
  assign io_in_instrctrs_22_iters = iters_x717_inr_Foreach_io_count; // @[Ledger.scala 294:22:@78501.4]
  assign io_in_instrctrs_22_stalls = stalls_x717_inr_Foreach_io_count; // @[Ledger.scala 295:23:@78502.4]
  assign io_in_instrctrs_22_idles = idles_x717_inr_Foreach_io_count; // @[Ledger.scala 296:22:@78503.4]
  assign cycles_x717_inr_Foreach_clock = clock; // @[:@78476.4]
  assign cycles_x717_inr_Foreach_reset = reset; // @[:@78477.4]
  assign cycles_x717_inr_Foreach_io_enable = io_sigsIn_baseEn; // @[sm_x717_inr_Foreach.scala 78:41:@78481.4]
  assign iters_x717_inr_Foreach_clock = clock; // @[:@78479.4]
  assign iters_x717_inr_Foreach_reset = reset; // @[:@78480.4]
  assign iters_x717_inr_Foreach_io_enable = io_sigsIn_done & _T_521; // @[sm_x717_inr_Foreach.scala 79:40:@78486.4]
  assign stalls_x717_inr_Foreach_clock = clock; // @[:@78488.4]
  assign stalls_x717_inr_Foreach_reset = reset; // @[:@78489.4]
  assign stalls_x717_inr_Foreach_io_enable = io_sigsIn_baseEn & _T_523; // @[sm_x717_inr_Foreach.scala 82:41:@78495.4]
  assign idles_x717_inr_Foreach_clock = clock; // @[:@78491.4]
  assign idles_x717_inr_Foreach_reset = reset; // @[:@78492.4]
  assign idles_x717_inr_Foreach_io_enable = 1'h0; // @[sm_x717_inr_Foreach.scala 83:40:@78499.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@78511.4]
  assign x709_sub_1_clock = clock; // @[:@78562.4]
  assign x709_sub_1_reset = reset; // @[:@78563.4]
  assign x709_sub_1_io_a = __io_result; // @[Math.scala 192:17:@78564.4]
  assign x709_sub_1_io_b = io_in_x676_reg_rPort_0_output_0; // @[Math.scala 193:17:@78565.4]
  assign x709_sub_1_io_flow = io_in_x670_ready; // @[Math.scala 194:20:@78566.4]
  assign x757_sum_1_clock = clock; // @[:@78577.4]
  assign x757_sum_1_reset = reset; // @[:@78578.4]
  assign x757_sum_1_io_a = _T_583[31:0]; // @[Math.scala 151:17:@78579.4]
  assign x757_sum_1_io_b = io_in_b674_number; // @[Math.scala 152:17:@78580.4]
  assign x757_sum_1_io_flow = io_in_x670_ready; // @[Math.scala 153:20:@78581.4]
  assign x712_sum_1_clock = clock; // @[:@78587.4]
  assign x712_sum_1_reset = reset; // @[:@78588.4]
  assign x712_sum_1_io_a = x757_sum_1_io_result; // @[Math.scala 151:17:@78589.4]
  assign x712_sum_1_io_b = x709_sub_1_io_result; // @[Math.scala 152:17:@78590.4]
  assign x712_sum_1_io_flow = io_in_x670_ready; // @[Math.scala 153:20:@78591.4]
  assign RetimeWrapper_clock = clock; // @[:@78598.4]
  assign RetimeWrapper_reset = reset; // @[:@78599.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@78601.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@78600.4]
  assign RetimeWrapper_1_clock = clock; // @[:@78608.4]
  assign RetimeWrapper_1_reset = reset; // @[:@78609.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@78611.4]
  assign RetimeWrapper_1_io_in = x705 & x707; // @[package.scala 94:16:@78610.4]
  assign RetimeWrapper_2_clock = clock; // @[:@78620.4]
  assign RetimeWrapper_2_reset = reset; // @[:@78621.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@78623.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@78622.4]
  assign RetimeWrapper_3_clock = clock; // @[:@78632.4]
  assign RetimeWrapper_3_reset = reset; // @[:@78633.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@78635.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@78634.4]
  assign RetimeWrapper_4_clock = clock; // @[:@78653.4]
  assign RetimeWrapper_4_reset = reset; // @[:@78654.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@78656.4]
  assign RetimeWrapper_4_io_in = x705 & x707; // @[package.scala 94:16:@78655.4]
  assign RetimeWrapper_5_clock = clock; // @[:@78666.4]
  assign RetimeWrapper_5_reset = reset; // @[:@78667.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@78669.4]
  assign RetimeWrapper_5_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@78668.4]
  assign RetimeWrapper_6_clock = clock; // @[:@78676.4]
  assign RetimeWrapper_6_reset = reset; // @[:@78677.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@78679.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@78678.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_521 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_521 <= 1'h0;
    end else begin
      _T_521 <= _T_518;
    end
  end
endmodule
module x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1( // @[:@78691.2]
  input         clock, // @[:@78692.4]
  input         reset, // @[:@78693.4]
  input         io_in_x670_ready, // @[:@78694.4]
  output        io_in_x670_valid, // @[:@78694.4]
  output [31:0] io_in_x670_bits_wdata_0, // @[:@78694.4]
  output        io_in_x670_bits_wstrb, // @[:@78694.4]
  input         io_in_x669_ready, // @[:@78694.4]
  output        io_in_x669_valid, // @[:@78694.4]
  output [63:0] io_in_x669_bits_addr, // @[:@78694.4]
  output [31:0] io_in_x669_bits_size, // @[:@78694.4]
  input  [31:0] io_in_b674_number, // @[:@78694.4]
  input  [63:0] io_in_x470_out_host_number, // @[:@78694.4]
  output [8:0]  io_in_x539_out_sram_0_rPort_0_ofs_0, // @[:@78694.4]
  output        io_in_x539_out_sram_0_rPort_0_en_0, // @[:@78694.4]
  output        io_in_x539_out_sram_0_rPort_0_backpressure, // @[:@78694.4]
  input  [31:0] io_in_x539_out_sram_0_rPort_0_output_0, // @[:@78694.4]
  output [63:0] io_in_instrctrs_20_cycs, // @[:@78694.4]
  output [63:0] io_in_instrctrs_20_iters, // @[:@78694.4]
  output [63:0] io_in_instrctrs_21_cycs, // @[:@78694.4]
  output [63:0] io_in_instrctrs_21_iters, // @[:@78694.4]
  output [63:0] io_in_instrctrs_21_stalls, // @[:@78694.4]
  output [63:0] io_in_instrctrs_21_idles, // @[:@78694.4]
  output [63:0] io_in_instrctrs_22_cycs, // @[:@78694.4]
  output [63:0] io_in_instrctrs_22_iters, // @[:@78694.4]
  output [63:0] io_in_instrctrs_22_stalls, // @[:@78694.4]
  output [63:0] io_in_instrctrs_22_idles, // @[:@78694.4]
  input         io_sigsIn_done, // @[:@78694.4]
  input         io_sigsIn_baseEn, // @[:@78694.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@78694.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@78694.4]
  input         io_sigsIn_smChildAcks_0, // @[:@78694.4]
  input         io_sigsIn_smChildAcks_1, // @[:@78694.4]
  output        io_sigsOut_smDoneIn_0, // @[:@78694.4]
  output        io_sigsOut_smDoneIn_1, // @[:@78694.4]
  output        io_sigsOut_smMaskIn_1, // @[:@78694.4]
  input         io_rr // @[:@78694.4]
);
  wire  cycles_x718_outr_UnitPipe_clock; // @[sm_x718_outr_UnitPipe.scala 82:45:@78815.4]
  wire  cycles_x718_outr_UnitPipe_reset; // @[sm_x718_outr_UnitPipe.scala 82:45:@78815.4]
  wire  cycles_x718_outr_UnitPipe_io_enable; // @[sm_x718_outr_UnitPipe.scala 82:45:@78815.4]
  wire [63:0] cycles_x718_outr_UnitPipe_io_count; // @[sm_x718_outr_UnitPipe.scala 82:45:@78815.4]
  wire  iters_x718_outr_UnitPipe_clock; // @[sm_x718_outr_UnitPipe.scala 83:44:@78818.4]
  wire  iters_x718_outr_UnitPipe_reset; // @[sm_x718_outr_UnitPipe.scala 83:44:@78818.4]
  wire  iters_x718_outr_UnitPipe_io_enable; // @[sm_x718_outr_UnitPipe.scala 83:44:@78818.4]
  wire [63:0] iters_x718_outr_UnitPipe_io_count; // @[sm_x718_outr_UnitPipe.scala 83:44:@78818.4]
  wire  x676_reg_clock; // @[m_x676_reg.scala 27:22:@78831.4]
  wire  x676_reg_reset; // @[m_x676_reg.scala 27:22:@78831.4]
  wire [31:0] x676_reg_io_rPort_0_output_0; // @[m_x676_reg.scala 27:22:@78831.4]
  wire [31:0] x676_reg_io_wPort_0_data_0; // @[m_x676_reg.scala 27:22:@78831.4]
  wire  x676_reg_io_wPort_0_reset; // @[m_x676_reg.scala 27:22:@78831.4]
  wire  x676_reg_io_wPort_0_en_0; // @[m_x676_reg.scala 27:22:@78831.4]
  wire  x677_reg_clock; // @[m_x677_reg.scala 27:22:@78848.4]
  wire  x677_reg_reset; // @[m_x677_reg.scala 27:22:@78848.4]
  wire [31:0] x677_reg_io_rPort_0_output_0; // @[m_x677_reg.scala 27:22:@78848.4]
  wire [31:0] x677_reg_io_wPort_0_data_0; // @[m_x677_reg.scala 27:22:@78848.4]
  wire  x677_reg_io_wPort_0_reset; // @[m_x677_reg.scala 27:22:@78848.4]
  wire  x677_reg_io_wPort_0_en_0; // @[m_x677_reg.scala 27:22:@78848.4]
  wire  x678_reg_clock; // @[m_x678_reg.scala 27:22:@78865.4]
  wire  x678_reg_reset; // @[m_x678_reg.scala 27:22:@78865.4]
  wire [31:0] x678_reg_io_rPort_0_output_0; // @[m_x678_reg.scala 27:22:@78865.4]
  wire [31:0] x678_reg_io_wPort_0_data_0; // @[m_x678_reg.scala 27:22:@78865.4]
  wire  x678_reg_io_wPort_0_reset; // @[m_x678_reg.scala 27:22:@78865.4]
  wire  x678_reg_io_wPort_0_en_0; // @[m_x678_reg.scala 27:22:@78865.4]
  wire  x698_inr_UnitPipe_sm_clock; // @[sm_x698_inr_UnitPipe.scala 34:18:@78918.4]
  wire  x698_inr_UnitPipe_sm_reset; // @[sm_x698_inr_UnitPipe.scala 34:18:@78918.4]
  wire  x698_inr_UnitPipe_sm_io_enable; // @[sm_x698_inr_UnitPipe.scala 34:18:@78918.4]
  wire  x698_inr_UnitPipe_sm_io_done; // @[sm_x698_inr_UnitPipe.scala 34:18:@78918.4]
  wire  x698_inr_UnitPipe_sm_io_doneLatch; // @[sm_x698_inr_UnitPipe.scala 34:18:@78918.4]
  wire  x698_inr_UnitPipe_sm_io_rst; // @[sm_x698_inr_UnitPipe.scala 34:18:@78918.4]
  wire  x698_inr_UnitPipe_sm_io_ctrDone; // @[sm_x698_inr_UnitPipe.scala 34:18:@78918.4]
  wire  x698_inr_UnitPipe_sm_io_datapathEn; // @[sm_x698_inr_UnitPipe.scala 34:18:@78918.4]
  wire  x698_inr_UnitPipe_sm_io_ctrInc; // @[sm_x698_inr_UnitPipe.scala 34:18:@78918.4]
  wire  x698_inr_UnitPipe_sm_io_ctrRst; // @[sm_x698_inr_UnitPipe.scala 34:18:@78918.4]
  wire  x698_inr_UnitPipe_sm_io_parentAck; // @[sm_x698_inr_UnitPipe.scala 34:18:@78918.4]
  wire  x698_inr_UnitPipe_sm_io_backpressure; // @[sm_x698_inr_UnitPipe.scala 34:18:@78918.4]
  wire  x698_inr_UnitPipe_sm_io_break; // @[sm_x698_inr_UnitPipe.scala 34:18:@78918.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@78976.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@78976.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@78976.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@78976.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@78976.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@78984.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@78984.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@78984.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@78984.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@78984.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_clock; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_reset; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire [31:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_data_0; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_reset; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_en_0; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_reset; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire [31:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_data_0; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_reset; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_en_0; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_reset; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_ready; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_valid; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire [63:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_bits_addr; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire [31:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_bits_size; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire [31:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_b674_number; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire [63:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x470_out_host_number; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire [31:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_data_0; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_reset; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_en_0; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_reset; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire [63:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_instrctrs_21_cycs; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire [63:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_instrctrs_21_iters; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire [63:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_instrctrs_21_stalls; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire [63:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_instrctrs_21_idles; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_done; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_baseEn; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_break; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_rr; // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
  wire  x701_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@79257.4]
  wire  x701_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@79257.4]
  wire [31:0] x701_ctrchain_io_setup_stops_0; // @[SpatialBlocks.scala 37:22:@79257.4]
  wire  x701_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@79257.4]
  wire  x701_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@79257.4]
  wire [31:0] x701_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@79257.4]
  wire  x701_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@79257.4]
  wire  x701_ctrchain_io_output_noop; // @[SpatialBlocks.scala 37:22:@79257.4]
  wire  x701_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@79257.4]
  wire  x717_inr_Foreach_sm_clock; // @[sm_x717_inr_Foreach.scala 34:18:@79312.4]
  wire  x717_inr_Foreach_sm_reset; // @[sm_x717_inr_Foreach.scala 34:18:@79312.4]
  wire  x717_inr_Foreach_sm_io_enable; // @[sm_x717_inr_Foreach.scala 34:18:@79312.4]
  wire  x717_inr_Foreach_sm_io_done; // @[sm_x717_inr_Foreach.scala 34:18:@79312.4]
  wire  x717_inr_Foreach_sm_io_doneLatch; // @[sm_x717_inr_Foreach.scala 34:18:@79312.4]
  wire  x717_inr_Foreach_sm_io_ctrDone; // @[sm_x717_inr_Foreach.scala 34:18:@79312.4]
  wire  x717_inr_Foreach_sm_io_datapathEn; // @[sm_x717_inr_Foreach.scala 34:18:@79312.4]
  wire  x717_inr_Foreach_sm_io_ctrInc; // @[sm_x717_inr_Foreach.scala 34:18:@79312.4]
  wire  x717_inr_Foreach_sm_io_ctrRst; // @[sm_x717_inr_Foreach.scala 34:18:@79312.4]
  wire  x717_inr_Foreach_sm_io_parentAck; // @[sm_x717_inr_Foreach.scala 34:18:@79312.4]
  wire  x717_inr_Foreach_sm_io_backpressure; // @[sm_x717_inr_Foreach.scala 34:18:@79312.4]
  wire  x717_inr_Foreach_sm_io_break; // @[sm_x717_inr_Foreach.scala 34:18:@79312.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@79341.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@79341.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@79341.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@79341.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@79341.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@79381.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@79381.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@79381.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@79381.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@79381.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@79389.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@79389.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@79389.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@79389.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@79389.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_clock; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_reset; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire [31:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x677_reg_rPort_0_output_0; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_ready; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_valid; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire [31:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_bits_wdata_0; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_bits_wstrb; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire [31:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_b674_number; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire [8:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_en_0; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire [31:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_output_0; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire [31:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x676_reg_rPort_0_output_0; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire [63:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_instrctrs_22_cycs; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire [63:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_instrctrs_22_iters; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire [63:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_instrctrs_22_stalls; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire [63:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_instrctrs_22_idles; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_done; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire [31:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_rr; // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
  wire  _T_276; // @[package.scala 100:49:@78822.4]
  reg  _T_279; // @[package.scala 48:56:@78823.4]
  reg [31:0] _RAND_0;
  wire  _T_344; // @[package.scala 100:49:@78946.4]
  reg  _T_347; // @[package.scala 48:56:@78947.4]
  reg [31:0] _RAND_1;
  wire  _T_362; // @[package.scala 96:25:@78981.4 package.scala 96:25:@78982.4]
  wire  _T_368; // @[package.scala 96:25:@78989.4 package.scala 96:25:@78990.4]
  wire  _T_371; // @[SpatialBlocks.scala 137:99:@78992.4]
  wire [31:0] x737_rd_x678_number; // @[sm_x718_outr_UnitPipe.scala 99:30:@79243.4 sm_x718_outr_UnitPipe.scala 104:202:@79256.4]
  wire  _T_459; // @[package.scala 96:25:@79346.4 package.scala 96:25:@79347.4]
  wire  x717_inr_Foreach_mySignalsIn_mask; // @[sm_x718_outr_UnitPipe.scala 115:32:@79357.4]
  wire  _T_475; // @[package.scala 96:25:@79386.4 package.scala 96:25:@79387.4]
  wire  _T_481; // @[package.scala 96:25:@79394.4 package.scala 96:25:@79395.4]
  wire  _T_484; // @[SpatialBlocks.scala 137:99:@79397.4]
  wire  _T_486; // @[SpatialBlocks.scala 156:36:@79406.4]
  wire  _T_487; // @[SpatialBlocks.scala 156:78:@79407.4]
  InstrumentationCounter cycles_x718_outr_UnitPipe ( // @[sm_x718_outr_UnitPipe.scala 82:45:@78815.4]
    .clock(cycles_x718_outr_UnitPipe_clock),
    .reset(cycles_x718_outr_UnitPipe_reset),
    .io_enable(cycles_x718_outr_UnitPipe_io_enable),
    .io_count(cycles_x718_outr_UnitPipe_io_count)
  );
  InstrumentationCounter iters_x718_outr_UnitPipe ( // @[sm_x718_outr_UnitPipe.scala 83:44:@78818.4]
    .clock(iters_x718_outr_UnitPipe_clock),
    .reset(iters_x718_outr_UnitPipe_reset),
    .io_enable(iters_x718_outr_UnitPipe_io_enable),
    .io_count(iters_x718_outr_UnitPipe_io_count)
  );
  x505_reg x676_reg ( // @[m_x676_reg.scala 27:22:@78831.4]
    .clock(x676_reg_clock),
    .reset(x676_reg_reset),
    .io_rPort_0_output_0(x676_reg_io_rPort_0_output_0),
    .io_wPort_0_data_0(x676_reg_io_wPort_0_data_0),
    .io_wPort_0_reset(x676_reg_io_wPort_0_reset),
    .io_wPort_0_en_0(x676_reg_io_wPort_0_en_0)
  );
  x505_reg x677_reg ( // @[m_x677_reg.scala 27:22:@78848.4]
    .clock(x677_reg_clock),
    .reset(x677_reg_reset),
    .io_rPort_0_output_0(x677_reg_io_rPort_0_output_0),
    .io_wPort_0_data_0(x677_reg_io_wPort_0_data_0),
    .io_wPort_0_reset(x677_reg_io_wPort_0_reset),
    .io_wPort_0_en_0(x677_reg_io_wPort_0_en_0)
  );
  x505_reg x678_reg ( // @[m_x678_reg.scala 27:22:@78865.4]
    .clock(x678_reg_clock),
    .reset(x678_reg_reset),
    .io_rPort_0_output_0(x678_reg_io_rPort_0_output_0),
    .io_wPort_0_data_0(x678_reg_io_wPort_0_data_0),
    .io_wPort_0_reset(x678_reg_io_wPort_0_reset),
    .io_wPort_0_en_0(x678_reg_io_wPort_0_en_0)
  );
  x499_inr_Foreach_sm x698_inr_UnitPipe_sm ( // @[sm_x698_inr_UnitPipe.scala 34:18:@78918.4]
    .clock(x698_inr_UnitPipe_sm_clock),
    .reset(x698_inr_UnitPipe_sm_reset),
    .io_enable(x698_inr_UnitPipe_sm_io_enable),
    .io_done(x698_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x698_inr_UnitPipe_sm_io_doneLatch),
    .io_rst(x698_inr_UnitPipe_sm_io_rst),
    .io_ctrDone(x698_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x698_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x698_inr_UnitPipe_sm_io_ctrInc),
    .io_ctrRst(x698_inr_UnitPipe_sm_io_ctrRst),
    .io_parentAck(x698_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x698_inr_UnitPipe_sm_io_backpressure),
    .io_break(x698_inr_UnitPipe_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@78976.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@78984.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1 x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1 ( // @[sm_x698_inr_UnitPipe.scala 146:24:@79013.4]
    .clock(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_clock),
    .reset(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_reset),
    .io_in_x677_reg_wPort_0_data_0(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_data_0),
    .io_in_x677_reg_wPort_0_reset(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_reset),
    .io_in_x677_reg_wPort_0_en_0(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_en_0),
    .io_in_x677_reg_reset(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_reset),
    .io_in_x678_reg_wPort_0_data_0(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_data_0),
    .io_in_x678_reg_wPort_0_reset(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_reset),
    .io_in_x678_reg_wPort_0_en_0(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_en_0),
    .io_in_x678_reg_reset(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_reset),
    .io_in_x669_ready(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_ready),
    .io_in_x669_valid(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_valid),
    .io_in_x669_bits_addr(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_bits_addr),
    .io_in_x669_bits_size(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_bits_size),
    .io_in_b674_number(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_b674_number),
    .io_in_x470_out_host_number(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x470_out_host_number),
    .io_in_x676_reg_wPort_0_data_0(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_data_0),
    .io_in_x676_reg_wPort_0_reset(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_reset),
    .io_in_x676_reg_wPort_0_en_0(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_en_0),
    .io_in_x676_reg_reset(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_reset),
    .io_in_instrctrs_21_cycs(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_instrctrs_21_cycs),
    .io_in_instrctrs_21_iters(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_instrctrs_21_iters),
    .io_in_instrctrs_21_stalls(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_instrctrs_21_stalls),
    .io_in_instrctrs_21_idles(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_instrctrs_21_idles),
    .io_sigsIn_done(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_done),
    .io_sigsIn_backpressure(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_break),
    .io_rr(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_rr)
  );
  x519_ctrchain x701_ctrchain ( // @[SpatialBlocks.scala 37:22:@79257.4]
    .clock(x701_ctrchain_clock),
    .reset(x701_ctrchain_reset),
    .io_setup_stops_0(x701_ctrchain_io_setup_stops_0),
    .io_input_reset(x701_ctrchain_io_input_reset),
    .io_input_enable(x701_ctrchain_io_input_enable),
    .io_output_counts_0(x701_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x701_ctrchain_io_output_oobs_0),
    .io_output_noop(x701_ctrchain_io_output_noop),
    .io_output_done(x701_ctrchain_io_output_done)
  );
  x652_inr_Foreach_sm x717_inr_Foreach_sm ( // @[sm_x717_inr_Foreach.scala 34:18:@79312.4]
    .clock(x717_inr_Foreach_sm_clock),
    .reset(x717_inr_Foreach_sm_reset),
    .io_enable(x717_inr_Foreach_sm_io_enable),
    .io_done(x717_inr_Foreach_sm_io_done),
    .io_doneLatch(x717_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x717_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x717_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x717_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x717_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x717_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x717_inr_Foreach_sm_io_backpressure),
    .io_break(x717_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@79341.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@79381.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@79389.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1 x717_inr_Foreach_kernelx717_inr_Foreach_concrete1 ( // @[sm_x717_inr_Foreach.scala 138:24:@79423.4]
    .clock(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_clock),
    .reset(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_reset),
    .io_in_x677_reg_rPort_0_output_0(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x677_reg_rPort_0_output_0),
    .io_in_x670_ready(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_ready),
    .io_in_x670_valid(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_valid),
    .io_in_x670_bits_wdata_0(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_bits_wdata_0),
    .io_in_x670_bits_wstrb(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_bits_wstrb),
    .io_in_b674_number(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_b674_number),
    .io_in_x539_out_sram_0_rPort_0_ofs_0(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0),
    .io_in_x539_out_sram_0_rPort_0_en_0(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_en_0),
    .io_in_x539_out_sram_0_rPort_0_backpressure(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure),
    .io_in_x539_out_sram_0_rPort_0_output_0(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_output_0),
    .io_in_x676_reg_rPort_0_output_0(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x676_reg_rPort_0_output_0),
    .io_in_instrctrs_22_cycs(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_instrctrs_22_cycs),
    .io_in_instrctrs_22_iters(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_instrctrs_22_iters),
    .io_in_instrctrs_22_stalls(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_instrctrs_22_stalls),
    .io_in_instrctrs_22_idles(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_instrctrs_22_idles),
    .io_sigsIn_done(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_backpressure(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_rr)
  );
  assign _T_276 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@78822.4]
  assign _T_344 = x698_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@78946.4]
  assign _T_362 = RetimeWrapper_io_out; // @[package.scala 96:25:@78981.4 package.scala 96:25:@78982.4]
  assign _T_368 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@78989.4 package.scala 96:25:@78990.4]
  assign _T_371 = ~ _T_368; // @[SpatialBlocks.scala 137:99:@78992.4]
  assign x737_rd_x678_number = x678_reg_io_rPort_0_output_0; // @[sm_x718_outr_UnitPipe.scala 99:30:@79243.4 sm_x718_outr_UnitPipe.scala 104:202:@79256.4]
  assign _T_459 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@79346.4 package.scala 96:25:@79347.4]
  assign x717_inr_Foreach_mySignalsIn_mask = ~ x701_ctrchain_io_output_noop; // @[sm_x718_outr_UnitPipe.scala 115:32:@79357.4]
  assign _T_475 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@79386.4 package.scala 96:25:@79387.4]
  assign _T_481 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@79394.4 package.scala 96:25:@79395.4]
  assign _T_484 = ~ _T_481; // @[SpatialBlocks.scala 137:99:@79397.4]
  assign _T_486 = x717_inr_Foreach_sm_io_datapathEn & x717_inr_Foreach_mySignalsIn_mask; // @[SpatialBlocks.scala 156:36:@79406.4]
  assign _T_487 = ~ x717_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 156:78:@79407.4]
  assign io_in_x670_valid = x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_valid; // @[sm_x717_inr_Foreach.scala 58:23:@79601.4]
  assign io_in_x670_bits_wdata_0 = x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_bits_wdata_0; // @[sm_x717_inr_Foreach.scala 58:23:@79600.4]
  assign io_in_x670_bits_wstrb = x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_bits_wstrb; // @[sm_x717_inr_Foreach.scala 58:23:@79599.4]
  assign io_in_x669_valid = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_valid; // @[sm_x698_inr_UnitPipe.scala 61:23:@79201.4]
  assign io_in_x669_bits_addr = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_bits_addr; // @[sm_x698_inr_UnitPipe.scala 61:23:@79200.4]
  assign io_in_x669_bits_size = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_bits_size; // @[sm_x698_inr_UnitPipe.scala 61:23:@79199.4]
  assign io_in_x539_out_sram_0_rPort_0_ofs_0 = x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@79607.4]
  assign io_in_x539_out_sram_0_rPort_0_en_0 = x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@79606.4]
  assign io_in_x539_out_sram_0_rPort_0_backpressure = x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@79605.4]
  assign io_in_instrctrs_20_cycs = cycles_x718_outr_UnitPipe_io_count; // @[Ledger.scala 293:21:@78827.4]
  assign io_in_instrctrs_20_iters = iters_x718_outr_UnitPipe_io_count; // @[Ledger.scala 294:22:@78828.4]
  assign io_in_instrctrs_21_cycs = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_instrctrs_21_cycs; // @[Ledger.scala 302:78:@79215.4]
  assign io_in_instrctrs_21_iters = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_instrctrs_21_iters; // @[Ledger.scala 302:78:@79214.4]
  assign io_in_instrctrs_21_stalls = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_instrctrs_21_stalls; // @[Ledger.scala 302:78:@79213.4]
  assign io_in_instrctrs_21_idles = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_instrctrs_21_idles; // @[Ledger.scala 302:78:@79212.4]
  assign io_in_instrctrs_22_cycs = x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_instrctrs_22_cycs; // @[Ledger.scala 302:78:@79617.4]
  assign io_in_instrctrs_22_iters = x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_instrctrs_22_iters; // @[Ledger.scala 302:78:@79616.4]
  assign io_in_instrctrs_22_stalls = x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_instrctrs_22_stalls; // @[Ledger.scala 302:78:@79615.4]
  assign io_in_instrctrs_22_idles = x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_instrctrs_22_idles; // @[Ledger.scala 302:78:@79614.4]
  assign io_sigsOut_smDoneIn_0 = x698_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 155:56:@78999.4]
  assign io_sigsOut_smDoneIn_1 = x717_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@79404.4]
  assign io_sigsOut_smMaskIn_1 = ~ x701_ctrchain_io_output_noop; // @[SpatialBlocks.scala 155:86:@79405.4]
  assign cycles_x718_outr_UnitPipe_clock = clock; // @[:@78816.4]
  assign cycles_x718_outr_UnitPipe_reset = reset; // @[:@78817.4]
  assign cycles_x718_outr_UnitPipe_io_enable = io_sigsIn_baseEn; // @[sm_x718_outr_UnitPipe.scala 84:43:@78821.4]
  assign iters_x718_outr_UnitPipe_clock = clock; // @[:@78819.4]
  assign iters_x718_outr_UnitPipe_reset = reset; // @[:@78820.4]
  assign iters_x718_outr_UnitPipe_io_enable = io_sigsIn_done & _T_279; // @[sm_x718_outr_UnitPipe.scala 85:42:@78826.4]
  assign x676_reg_clock = clock; // @[:@78832.4]
  assign x676_reg_reset = reset; // @[:@78833.4]
  assign x676_reg_io_wPort_0_data_0 = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@79209.4]
  assign x676_reg_io_wPort_0_reset = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_reset; // @[MemInterfaceType.scala 67:44:@79208.4]
  assign x676_reg_io_wPort_0_en_0 = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@79205.4]
  assign x677_reg_clock = clock; // @[:@78849.4]
  assign x677_reg_reset = reset; // @[:@78850.4]
  assign x677_reg_io_wPort_0_data_0 = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@79189.4]
  assign x677_reg_io_wPort_0_reset = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_reset; // @[MemInterfaceType.scala 67:44:@79188.4]
  assign x677_reg_io_wPort_0_en_0 = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@79185.4]
  assign x678_reg_clock = clock; // @[:@78866.4]
  assign x678_reg_reset = reset; // @[:@78867.4]
  assign x678_reg_io_wPort_0_data_0 = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@79196.4]
  assign x678_reg_io_wPort_0_reset = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_reset; // @[MemInterfaceType.scala 67:44:@79195.4]
  assign x678_reg_io_wPort_0_en_0 = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@79192.4]
  assign x698_inr_UnitPipe_sm_clock = clock; // @[:@78919.4]
  assign x698_inr_UnitPipe_sm_reset = reset; // @[:@78920.4]
  assign x698_inr_UnitPipe_sm_io_enable = _T_362 & _T_371; // @[SpatialBlocks.scala 139:18:@78996.4]
  assign x698_inr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 133:15:@78971.4]
  assign x698_inr_UnitPipe_sm_io_ctrDone = x698_inr_UnitPipe_sm_io_ctrInc & _T_347; // @[sm_x718_outr_UnitPipe.scala 91:39:@78950.4]
  assign x698_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@78998.4]
  assign x698_inr_UnitPipe_sm_io_backpressure = io_in_x669_ready | x698_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 132:24:@78970.4]
  assign x698_inr_UnitPipe_sm_io_break = 1'h0; // @[sm_x718_outr_UnitPipe.scala 95:37:@78957.4]
  assign RetimeWrapper_clock = clock; // @[:@78977.4]
  assign RetimeWrapper_reset = reset; // @[:@78978.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@78980.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@78979.4]
  assign RetimeWrapper_1_clock = clock; // @[:@78985.4]
  assign RetimeWrapper_1_reset = reset; // @[:@78986.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@78988.4]
  assign RetimeWrapper_1_io_in = x698_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@78987.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_clock = clock; // @[:@79014.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_reset = reset; // @[:@79015.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_ready = io_in_x669_ready; // @[sm_x698_inr_UnitPipe.scala 61:23:@79202.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_b674_number = io_in_b674_number; // @[sm_x698_inr_UnitPipe.scala 62:23:@79203.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x470_out_host_number = io_in_x470_out_host_number; // @[sm_x698_inr_UnitPipe.scala 63:32:@79204.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_done = x698_inr_UnitPipe_sm_io_done; // @[sm_x698_inr_UnitPipe.scala 152:22:@79235.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x669_ready | x698_inr_UnitPipe_sm_io_doneLatch; // @[sm_x698_inr_UnitPipe.scala 152:22:@79230.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x698_inr_UnitPipe_sm_io_datapathEn; // @[sm_x698_inr_UnitPipe.scala 152:22:@79228.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_baseEn = _T_362 & _T_371; // @[sm_x698_inr_UnitPipe.scala 152:22:@79227.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_break = x698_inr_UnitPipe_sm_io_break; // @[sm_x698_inr_UnitPipe.scala 152:22:@79226.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x698_inr_UnitPipe.scala 151:18:@79216.4]
  assign x701_ctrchain_clock = clock; // @[:@79258.4]
  assign x701_ctrchain_reset = reset; // @[:@79259.4]
  assign x701_ctrchain_io_setup_stops_0 = $signed(x737_rd_x678_number); // @[SpatialBlocks.scala 40:87:@79273.4]
  assign x701_ctrchain_io_input_reset = x717_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@79422.4]
  assign x701_ctrchain_io_input_enable = x717_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 158:42:@79421.4]
  assign x717_inr_Foreach_sm_clock = clock; // @[:@79313.4]
  assign x717_inr_Foreach_sm_reset = reset; // @[:@79314.4]
  assign x717_inr_Foreach_sm_io_enable = _T_475 & _T_484; // @[SpatialBlocks.scala 139:18:@79401.4]
  assign x717_inr_Foreach_sm_io_ctrDone = io_rr ? _T_459 : 1'h0; // @[sm_x718_outr_UnitPipe.scala 110:38:@79349.4]
  assign x717_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 141:21:@79403.4]
  assign x717_inr_Foreach_sm_io_backpressure = io_in_x670_ready | x717_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 132:24:@79375.4]
  assign x717_inr_Foreach_sm_io_break = 1'h0; // @[sm_x718_outr_UnitPipe.scala 114:36:@79356.4]
  assign RetimeWrapper_2_clock = clock; // @[:@79342.4]
  assign RetimeWrapper_2_reset = reset; // @[:@79343.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@79345.4]
  assign RetimeWrapper_2_io_in = x701_ctrchain_io_output_done; // @[package.scala 94:16:@79344.4]
  assign RetimeWrapper_3_clock = clock; // @[:@79382.4]
  assign RetimeWrapper_3_reset = reset; // @[:@79383.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@79385.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@79384.4]
  assign RetimeWrapper_4_clock = clock; // @[:@79390.4]
  assign RetimeWrapper_4_reset = reset; // @[:@79391.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@79393.4]
  assign RetimeWrapper_4_io_in = x717_inr_Foreach_sm_io_done; // @[package.scala 94:16:@79392.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_clock = clock; // @[:@79424.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_reset = reset; // @[:@79425.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x677_reg_rPort_0_output_0 = x677_reg_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@79594.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_ready = io_in_x670_ready; // @[sm_x717_inr_Foreach.scala 58:23:@79602.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_b674_number = io_in_b674_number; // @[sm_x717_inr_Foreach.scala 59:23:@79603.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_output_0 = io_in_x539_out_sram_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@79604.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x676_reg_rPort_0_output_0 = x676_reg_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@79609.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_done = x717_inr_Foreach_sm_io_done; // @[sm_x717_inr_Foreach.scala 144:22:@79637.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x670_ready | x717_inr_Foreach_sm_io_doneLatch; // @[sm_x717_inr_Foreach.scala 144:22:@79632.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_486 & _T_487; // @[sm_x717_inr_Foreach.scala 144:22:@79630.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_baseEn = _T_475 & _T_484; // @[sm_x717_inr_Foreach.scala 144:22:@79629.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_break = x717_inr_Foreach_sm_io_break; // @[sm_x717_inr_Foreach.scala 144:22:@79628.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x701_ctrchain_io_output_counts_0; // @[sm_x717_inr_Foreach.scala 144:22:@79623.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x701_ctrchain_io_output_oobs_0; // @[sm_x717_inr_Foreach.scala 144:22:@79622.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x717_inr_Foreach.scala 143:18:@79618.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_279 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_347 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_279 <= 1'h0;
    end else begin
      _T_279 <= _T_276;
    end
    if (reset) begin
      _T_347 <= 1'h0;
    end else begin
      _T_347 <= _T_344;
    end
  end
endmodule
module x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1( // @[:@80026.2]
  input         clock, // @[:@80027.4]
  input         reset, // @[:@80028.4]
  output        io_in_x671_ready, // @[:@80029.4]
  input         io_in_x671_valid, // @[:@80029.4]
  output [63:0] io_in_instrctrs_23_cycs, // @[:@80029.4]
  output [63:0] io_in_instrctrs_23_iters, // @[:@80029.4]
  output [63:0] io_in_instrctrs_23_stalls, // @[:@80029.4]
  output [63:0] io_in_instrctrs_23_idles, // @[:@80029.4]
  input         io_sigsIn_done, // @[:@80029.4]
  input         io_sigsIn_datapathEn, // @[:@80029.4]
  input         io_sigsIn_baseEn // @[:@80029.4]
);
  wire  cycles_x722_inr_UnitPipe_clock; // @[sm_x722_inr_UnitPipe.scala 63:44:@80135.4]
  wire  cycles_x722_inr_UnitPipe_reset; // @[sm_x722_inr_UnitPipe.scala 63:44:@80135.4]
  wire  cycles_x722_inr_UnitPipe_io_enable; // @[sm_x722_inr_UnitPipe.scala 63:44:@80135.4]
  wire [63:0] cycles_x722_inr_UnitPipe_io_count; // @[sm_x722_inr_UnitPipe.scala 63:44:@80135.4]
  wire  iters_x722_inr_UnitPipe_clock; // @[sm_x722_inr_UnitPipe.scala 64:43:@80138.4]
  wire  iters_x722_inr_UnitPipe_reset; // @[sm_x722_inr_UnitPipe.scala 64:43:@80138.4]
  wire  iters_x722_inr_UnitPipe_io_enable; // @[sm_x722_inr_UnitPipe.scala 64:43:@80138.4]
  wire [63:0] iters_x722_inr_UnitPipe_io_count; // @[sm_x722_inr_UnitPipe.scala 64:43:@80138.4]
  wire  stalls_x722_inr_UnitPipe_clock; // @[sm_x722_inr_UnitPipe.scala 67:44:@80147.4]
  wire  stalls_x722_inr_UnitPipe_reset; // @[sm_x722_inr_UnitPipe.scala 67:44:@80147.4]
  wire  stalls_x722_inr_UnitPipe_io_enable; // @[sm_x722_inr_UnitPipe.scala 67:44:@80147.4]
  wire [63:0] stalls_x722_inr_UnitPipe_io_count; // @[sm_x722_inr_UnitPipe.scala 67:44:@80147.4]
  wire  idles_x722_inr_UnitPipe_clock; // @[sm_x722_inr_UnitPipe.scala 68:43:@80150.4]
  wire  idles_x722_inr_UnitPipe_reset; // @[sm_x722_inr_UnitPipe.scala 68:43:@80150.4]
  wire  idles_x722_inr_UnitPipe_io_enable; // @[sm_x722_inr_UnitPipe.scala 68:43:@80150.4]
  wire [63:0] idles_x722_inr_UnitPipe_io_count; // @[sm_x722_inr_UnitPipe.scala 68:43:@80150.4]
  wire  _T_138; // @[package.scala 100:49:@80142.4]
  reg  _T_141; // @[package.scala 48:56:@80143.4]
  reg [31:0] _RAND_0;
  wire  _T_148; // @[sm_x722_inr_UnitPipe.scala 70:63:@80157.4]
  InstrumentationCounter cycles_x722_inr_UnitPipe ( // @[sm_x722_inr_UnitPipe.scala 63:44:@80135.4]
    .clock(cycles_x722_inr_UnitPipe_clock),
    .reset(cycles_x722_inr_UnitPipe_reset),
    .io_enable(cycles_x722_inr_UnitPipe_io_enable),
    .io_count(cycles_x722_inr_UnitPipe_io_count)
  );
  InstrumentationCounter iters_x722_inr_UnitPipe ( // @[sm_x722_inr_UnitPipe.scala 64:43:@80138.4]
    .clock(iters_x722_inr_UnitPipe_clock),
    .reset(iters_x722_inr_UnitPipe_reset),
    .io_enable(iters_x722_inr_UnitPipe_io_enable),
    .io_count(iters_x722_inr_UnitPipe_io_count)
  );
  InstrumentationCounter stalls_x722_inr_UnitPipe ( // @[sm_x722_inr_UnitPipe.scala 67:44:@80147.4]
    .clock(stalls_x722_inr_UnitPipe_clock),
    .reset(stalls_x722_inr_UnitPipe_reset),
    .io_enable(stalls_x722_inr_UnitPipe_io_enable),
    .io_count(stalls_x722_inr_UnitPipe_io_count)
  );
  InstrumentationCounter idles_x722_inr_UnitPipe ( // @[sm_x722_inr_UnitPipe.scala 68:43:@80150.4]
    .clock(idles_x722_inr_UnitPipe_clock),
    .reset(idles_x722_inr_UnitPipe_reset),
    .io_enable(idles_x722_inr_UnitPipe_io_enable),
    .io_count(idles_x722_inr_UnitPipe_io_count)
  );
  assign _T_138 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@80142.4]
  assign _T_148 = ~ io_in_x671_valid; // @[sm_x722_inr_UnitPipe.scala 70:63:@80157.4]
  assign io_in_x671_ready = io_sigsIn_datapathEn; // @[sm_x722_inr_UnitPipe.scala 73:18:@80166.4]
  assign io_in_instrctrs_23_cycs = cycles_x722_inr_UnitPipe_io_count; // @[Ledger.scala 293:21:@80160.4]
  assign io_in_instrctrs_23_iters = iters_x722_inr_UnitPipe_io_count; // @[Ledger.scala 294:22:@80161.4]
  assign io_in_instrctrs_23_stalls = stalls_x722_inr_UnitPipe_io_count; // @[Ledger.scala 295:23:@80162.4]
  assign io_in_instrctrs_23_idles = idles_x722_inr_UnitPipe_io_count; // @[Ledger.scala 296:22:@80163.4]
  assign cycles_x722_inr_UnitPipe_clock = clock; // @[:@80136.4]
  assign cycles_x722_inr_UnitPipe_reset = reset; // @[:@80137.4]
  assign cycles_x722_inr_UnitPipe_io_enable = io_sigsIn_baseEn; // @[sm_x722_inr_UnitPipe.scala 65:42:@80141.4]
  assign iters_x722_inr_UnitPipe_clock = clock; // @[:@80139.4]
  assign iters_x722_inr_UnitPipe_reset = reset; // @[:@80140.4]
  assign iters_x722_inr_UnitPipe_io_enable = io_sigsIn_done & _T_141; // @[sm_x722_inr_UnitPipe.scala 66:41:@80146.4]
  assign stalls_x722_inr_UnitPipe_clock = clock; // @[:@80148.4]
  assign stalls_x722_inr_UnitPipe_reset = reset; // @[:@80149.4]
  assign stalls_x722_inr_UnitPipe_io_enable = 1'h0; // @[sm_x722_inr_UnitPipe.scala 69:42:@80155.4]
  assign idles_x722_inr_UnitPipe_clock = clock; // @[:@80151.4]
  assign idles_x722_inr_UnitPipe_reset = reset; // @[:@80152.4]
  assign idles_x722_inr_UnitPipe_io_enable = io_sigsIn_baseEn & _T_148; // @[sm_x722_inr_UnitPipe.scala 70:41:@80159.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_141 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_141 <= 1'h0;
    end else begin
      _T_141 <= _T_138;
    end
  end
endmodule
module x723_outr_Foreach_kernelx723_outr_Foreach_concrete1( // @[:@80169.2]
  input         clock, // @[:@80170.4]
  input         reset, // @[:@80171.4]
  input         io_in_x670_ready, // @[:@80172.4]
  output        io_in_x670_valid, // @[:@80172.4]
  output [31:0] io_in_x670_bits_wdata_0, // @[:@80172.4]
  output        io_in_x670_bits_wstrb, // @[:@80172.4]
  input         io_in_x669_ready, // @[:@80172.4]
  output        io_in_x669_valid, // @[:@80172.4]
  output [63:0] io_in_x669_bits_addr, // @[:@80172.4]
  output [31:0] io_in_x669_bits_size, // @[:@80172.4]
  input  [63:0] io_in_x470_out_host_number, // @[:@80172.4]
  output [8:0]  io_in_x539_out_sram_0_rPort_0_ofs_0, // @[:@80172.4]
  output        io_in_x539_out_sram_0_rPort_0_en_0, // @[:@80172.4]
  output        io_in_x539_out_sram_0_rPort_0_backpressure, // @[:@80172.4]
  input  [31:0] io_in_x539_out_sram_0_rPort_0_output_0, // @[:@80172.4]
  output        io_in_x671_ready, // @[:@80172.4]
  input         io_in_x671_valid, // @[:@80172.4]
  output [63:0] io_in_instrctrs_19_cycs, // @[:@80172.4]
  output [63:0] io_in_instrctrs_19_iters, // @[:@80172.4]
  output [63:0] io_in_instrctrs_20_cycs, // @[:@80172.4]
  output [63:0] io_in_instrctrs_20_iters, // @[:@80172.4]
  output [63:0] io_in_instrctrs_21_cycs, // @[:@80172.4]
  output [63:0] io_in_instrctrs_21_iters, // @[:@80172.4]
  output [63:0] io_in_instrctrs_21_stalls, // @[:@80172.4]
  output [63:0] io_in_instrctrs_21_idles, // @[:@80172.4]
  output [63:0] io_in_instrctrs_22_cycs, // @[:@80172.4]
  output [63:0] io_in_instrctrs_22_iters, // @[:@80172.4]
  output [63:0] io_in_instrctrs_22_stalls, // @[:@80172.4]
  output [63:0] io_in_instrctrs_22_idles, // @[:@80172.4]
  output [63:0] io_in_instrctrs_23_cycs, // @[:@80172.4]
  output [63:0] io_in_instrctrs_23_iters, // @[:@80172.4]
  output [63:0] io_in_instrctrs_23_stalls, // @[:@80172.4]
  output [63:0] io_in_instrctrs_23_idles, // @[:@80172.4]
  input         io_sigsIn_done, // @[:@80172.4]
  input         io_sigsIn_baseEn, // @[:@80172.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@80172.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@80172.4]
  input         io_sigsIn_smChildAcks_0, // @[:@80172.4]
  input         io_sigsIn_smChildAcks_1, // @[:@80172.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@80172.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@80172.4]
  output        io_sigsOut_smDoneIn_0, // @[:@80172.4]
  output        io_sigsOut_smDoneIn_1, // @[:@80172.4]
  output        io_sigsOut_smMaskIn_0, // @[:@80172.4]
  output        io_sigsOut_smMaskIn_1, // @[:@80172.4]
  input         io_rr // @[:@80172.4]
);
  wire  cycles_x723_outr_Foreach_clock; // @[sm_x723_outr_Foreach.scala 78:44:@80293.4]
  wire  cycles_x723_outr_Foreach_reset; // @[sm_x723_outr_Foreach.scala 78:44:@80293.4]
  wire  cycles_x723_outr_Foreach_io_enable; // @[sm_x723_outr_Foreach.scala 78:44:@80293.4]
  wire [63:0] cycles_x723_outr_Foreach_io_count; // @[sm_x723_outr_Foreach.scala 78:44:@80293.4]
  wire  iters_x723_outr_Foreach_clock; // @[sm_x723_outr_Foreach.scala 79:43:@80296.4]
  wire  iters_x723_outr_Foreach_reset; // @[sm_x723_outr_Foreach.scala 79:43:@80296.4]
  wire  iters_x723_outr_Foreach_io_enable; // @[sm_x723_outr_Foreach.scala 79:43:@80296.4]
  wire [63:0] iters_x723_outr_Foreach_io_count; // @[sm_x723_outr_Foreach.scala 79:43:@80296.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@80313.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@80313.4]
  wire  x718_outr_UnitPipe_sm_clock; // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
  wire  x718_outr_UnitPipe_sm_reset; // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
  wire  x718_outr_UnitPipe_sm_io_enable; // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
  wire  x718_outr_UnitPipe_sm_io_done; // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
  wire  x718_outr_UnitPipe_sm_io_ctrDone; // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
  wire  x718_outr_UnitPipe_sm_io_ctrInc; // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
  wire  x718_outr_UnitPipe_sm_io_ctrRst; // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
  wire  x718_outr_UnitPipe_sm_io_parentAck; // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
  wire  x718_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
  wire  x718_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
  wire  x718_outr_UnitPipe_sm_io_maskIn_0; // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
  wire  x718_outr_UnitPipe_sm_io_maskIn_1; // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
  wire  x718_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
  wire  x718_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
  wire  x718_outr_UnitPipe_sm_io_childAck_0; // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
  wire  x718_outr_UnitPipe_sm_io_childAck_1; // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@80431.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@80431.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@80431.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@80431.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@80431.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@80439.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@80439.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@80439.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@80439.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@80439.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_clock; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_reset; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_ready; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_valid; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [31:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_bits_wdata_0; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_bits_wstrb; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_ready; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_valid; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [63:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_bits_addr; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [31:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_bits_size; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [31:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_b674_number; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [63:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x470_out_host_number; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [8:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_en_0; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [31:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_output_0; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [63:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_20_cycs; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [63:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_20_iters; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [63:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_21_cycs; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [63:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_21_iters; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [63:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_21_stalls; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [63:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_21_idles; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [63:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_22_cycs; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [63:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_22_iters; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [63:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_22_stalls; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire [63:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_22_idles; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_done; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_baseEn; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smMaskIn_1; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_rr; // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
  wire  x722_inr_UnitPipe_sm_clock; // @[sm_x722_inr_UnitPipe.scala 33:18:@80720.4]
  wire  x722_inr_UnitPipe_sm_reset; // @[sm_x722_inr_UnitPipe.scala 33:18:@80720.4]
  wire  x722_inr_UnitPipe_sm_io_enable; // @[sm_x722_inr_UnitPipe.scala 33:18:@80720.4]
  wire  x722_inr_UnitPipe_sm_io_done; // @[sm_x722_inr_UnitPipe.scala 33:18:@80720.4]
  wire  x722_inr_UnitPipe_sm_io_doneLatch; // @[sm_x722_inr_UnitPipe.scala 33:18:@80720.4]
  wire  x722_inr_UnitPipe_sm_io_ctrDone; // @[sm_x722_inr_UnitPipe.scala 33:18:@80720.4]
  wire  x722_inr_UnitPipe_sm_io_datapathEn; // @[sm_x722_inr_UnitPipe.scala 33:18:@80720.4]
  wire  x722_inr_UnitPipe_sm_io_ctrInc; // @[sm_x722_inr_UnitPipe.scala 33:18:@80720.4]
  wire  x722_inr_UnitPipe_sm_io_parentAck; // @[sm_x722_inr_UnitPipe.scala 33:18:@80720.4]
  wire  x722_inr_UnitPipe_sm_io_backpressure; // @[sm_x722_inr_UnitPipe.scala 33:18:@80720.4]
  wire  x722_inr_UnitPipe_sm_io_break; // @[sm_x722_inr_UnitPipe.scala 33:18:@80720.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@80778.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@80778.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@80778.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@80778.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@80778.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@80786.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@80786.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@80786.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@80786.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@80786.4]
  wire  x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_clock; // @[sm_x722_inr_UnitPipe.scala 76:24:@80815.4]
  wire  x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_reset; // @[sm_x722_inr_UnitPipe.scala 76:24:@80815.4]
  wire  x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_x671_ready; // @[sm_x722_inr_UnitPipe.scala 76:24:@80815.4]
  wire  x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_x671_valid; // @[sm_x722_inr_UnitPipe.scala 76:24:@80815.4]
  wire [63:0] x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_instrctrs_23_cycs; // @[sm_x722_inr_UnitPipe.scala 76:24:@80815.4]
  wire [63:0] x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_instrctrs_23_iters; // @[sm_x722_inr_UnitPipe.scala 76:24:@80815.4]
  wire [63:0] x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_instrctrs_23_stalls; // @[sm_x722_inr_UnitPipe.scala 76:24:@80815.4]
  wire [63:0] x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_instrctrs_23_idles; // @[sm_x722_inr_UnitPipe.scala 76:24:@80815.4]
  wire  x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_sigsIn_done; // @[sm_x722_inr_UnitPipe.scala 76:24:@80815.4]
  wire  x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x722_inr_UnitPipe.scala 76:24:@80815.4]
  wire  x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_sigsIn_baseEn; // @[sm_x722_inr_UnitPipe.scala 76:24:@80815.4]
  wire  _T_284; // @[package.scala 100:49:@80300.4]
  reg  _T_287; // @[package.scala 48:56:@80301.4]
  reg [31:0] _RAND_0;
  wire  b675; // @[sm_x723_outr_Foreach.scala 84:18:@80321.4]
  wire  _T_356; // @[package.scala 100:49:@80396.4]
  reg  _T_359; // @[package.scala 48:56:@80397.4]
  reg [31:0] _RAND_1;
  wire  _T_374; // @[package.scala 96:25:@80436.4 package.scala 96:25:@80437.4]
  wire  _T_380; // @[package.scala 96:25:@80444.4 package.scala 96:25:@80445.4]
  wire  _T_383; // @[SpatialBlocks.scala 137:99:@80447.4]
  wire  _T_451; // @[package.scala 100:49:@80748.4]
  reg  _T_454; // @[package.scala 48:56:@80749.4]
  reg [31:0] _RAND_2;
  wire  x722_inr_UnitPipe_mySignalsIn_forwardpressure; // @[sm_x723_outr_Foreach.scala 97:69:@80756.4]
  wire  _T_468; // @[package.scala 96:25:@80783.4 package.scala 96:25:@80784.4]
  wire  _T_474; // @[package.scala 96:25:@80791.4 package.scala 96:25:@80792.4]
  wire  _T_477; // @[SpatialBlocks.scala 137:99:@80794.4]
  wire  x722_inr_UnitPipe_mySignalsIn_baseEn; // @[SpatialBlocks.scala 137:96:@80795.4]
  InstrumentationCounter cycles_x723_outr_Foreach ( // @[sm_x723_outr_Foreach.scala 78:44:@80293.4]
    .clock(cycles_x723_outr_Foreach_clock),
    .reset(cycles_x723_outr_Foreach_reset),
    .io_enable(cycles_x723_outr_Foreach_io_enable),
    .io_count(cycles_x723_outr_Foreach_io_count)
  );
  InstrumentationCounter iters_x723_outr_Foreach ( // @[sm_x723_outr_Foreach.scala 79:43:@80296.4]
    .clock(iters_x723_outr_Foreach_clock),
    .reset(iters_x723_outr_Foreach_reset),
    .io_enable(iters_x723_outr_Foreach_io_enable),
    .io_count(iters_x723_outr_Foreach_io_count)
  );
  _ _ ( // @[Math.scala 720:24:@80313.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x537_outr_Foreach_sm x718_outr_UnitPipe_sm ( // @[sm_x718_outr_UnitPipe.scala 36:18:@80363.4]
    .clock(x718_outr_UnitPipe_sm_clock),
    .reset(x718_outr_UnitPipe_sm_reset),
    .io_enable(x718_outr_UnitPipe_sm_io_enable),
    .io_done(x718_outr_UnitPipe_sm_io_done),
    .io_ctrDone(x718_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x718_outr_UnitPipe_sm_io_ctrInc),
    .io_ctrRst(x718_outr_UnitPipe_sm_io_ctrRst),
    .io_parentAck(x718_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x718_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x718_outr_UnitPipe_sm_io_doneIn_1),
    .io_maskIn_0(x718_outr_UnitPipe_sm_io_maskIn_0),
    .io_maskIn_1(x718_outr_UnitPipe_sm_io_maskIn_1),
    .io_enableOut_0(x718_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x718_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x718_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x718_outr_UnitPipe_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@80431.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@80439.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1 x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1 ( // @[sm_x718_outr_UnitPipe.scala 119:24:@80468.4]
    .clock(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_clock),
    .reset(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_reset),
    .io_in_x670_ready(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_ready),
    .io_in_x670_valid(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_valid),
    .io_in_x670_bits_wdata_0(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_bits_wdata_0),
    .io_in_x670_bits_wstrb(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_bits_wstrb),
    .io_in_x669_ready(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_ready),
    .io_in_x669_valid(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_valid),
    .io_in_x669_bits_addr(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_bits_addr),
    .io_in_x669_bits_size(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_bits_size),
    .io_in_b674_number(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_b674_number),
    .io_in_x470_out_host_number(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x470_out_host_number),
    .io_in_x539_out_sram_0_rPort_0_ofs_0(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0),
    .io_in_x539_out_sram_0_rPort_0_en_0(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_en_0),
    .io_in_x539_out_sram_0_rPort_0_backpressure(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure),
    .io_in_x539_out_sram_0_rPort_0_output_0(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_output_0),
    .io_in_instrctrs_20_cycs(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_20_cycs),
    .io_in_instrctrs_20_iters(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_20_iters),
    .io_in_instrctrs_21_cycs(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_21_cycs),
    .io_in_instrctrs_21_iters(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_21_iters),
    .io_in_instrctrs_21_stalls(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_21_stalls),
    .io_in_instrctrs_21_idles(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_21_idles),
    .io_in_instrctrs_22_cycs(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_22_cycs),
    .io_in_instrctrs_22_iters(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_22_iters),
    .io_in_instrctrs_22_stalls(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_22_stalls),
    .io_in_instrctrs_22_idles(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_22_idles),
    .io_sigsIn_done(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smEnableOuts_0(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smMaskIn_1(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smMaskIn_1),
    .io_rr(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_rr)
  );
  x516_inr_UnitPipe_sm x722_inr_UnitPipe_sm ( // @[sm_x722_inr_UnitPipe.scala 33:18:@80720.4]
    .clock(x722_inr_UnitPipe_sm_clock),
    .reset(x722_inr_UnitPipe_sm_reset),
    .io_enable(x722_inr_UnitPipe_sm_io_enable),
    .io_done(x722_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x722_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x722_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x722_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x722_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x722_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x722_inr_UnitPipe_sm_io_backpressure),
    .io_break(x722_inr_UnitPipe_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@80778.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@80786.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1 x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1 ( // @[sm_x722_inr_UnitPipe.scala 76:24:@80815.4]
    .clock(x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_clock),
    .reset(x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_reset),
    .io_in_x671_ready(x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_x671_ready),
    .io_in_x671_valid(x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_x671_valid),
    .io_in_instrctrs_23_cycs(x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_instrctrs_23_cycs),
    .io_in_instrctrs_23_iters(x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_instrctrs_23_iters),
    .io_in_instrctrs_23_stalls(x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_instrctrs_23_stalls),
    .io_in_instrctrs_23_idles(x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_instrctrs_23_idles),
    .io_sigsIn_done(x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_sigsIn_done),
    .io_sigsIn_datapathEn(x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_sigsIn_baseEn)
  );
  assign _T_284 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@80300.4]
  assign b675 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x723_outr_Foreach.scala 84:18:@80321.4]
  assign _T_356 = x718_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@80396.4]
  assign _T_374 = RetimeWrapper_io_out; // @[package.scala 96:25:@80436.4 package.scala 96:25:@80437.4]
  assign _T_380 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@80444.4 package.scala 96:25:@80445.4]
  assign _T_383 = ~ _T_380; // @[SpatialBlocks.scala 137:99:@80447.4]
  assign _T_451 = x722_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@80748.4]
  assign x722_inr_UnitPipe_mySignalsIn_forwardpressure = io_in_x671_valid | x722_inr_UnitPipe_sm_io_doneLatch; // @[sm_x723_outr_Foreach.scala 97:69:@80756.4]
  assign _T_468 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@80783.4 package.scala 96:25:@80784.4]
  assign _T_474 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@80791.4 package.scala 96:25:@80792.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 137:99:@80794.4]
  assign x722_inr_UnitPipe_mySignalsIn_baseEn = _T_468 & _T_477; // @[SpatialBlocks.scala 137:96:@80795.4]
  assign io_in_x670_valid = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_valid; // @[sm_x718_outr_UnitPipe.scala 61:23:@80626.4]
  assign io_in_x670_bits_wdata_0 = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_bits_wdata_0; // @[sm_x718_outr_UnitPipe.scala 61:23:@80625.4]
  assign io_in_x670_bits_wstrb = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_bits_wstrb; // @[sm_x718_outr_UnitPipe.scala 61:23:@80624.4]
  assign io_in_x669_valid = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_valid; // @[sm_x718_outr_UnitPipe.scala 62:23:@80630.4]
  assign io_in_x669_bits_addr = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_bits_addr; // @[sm_x718_outr_UnitPipe.scala 62:23:@80629.4]
  assign io_in_x669_bits_size = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_bits_size; // @[sm_x718_outr_UnitPipe.scala 62:23:@80628.4]
  assign io_in_x539_out_sram_0_rPort_0_ofs_0 = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@80638.4]
  assign io_in_x539_out_sram_0_rPort_0_en_0 = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@80637.4]
  assign io_in_x539_out_sram_0_rPort_0_backpressure = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@80636.4]
  assign io_in_x671_ready = x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_x671_ready; // @[sm_x722_inr_UnitPipe.scala 51:23:@80949.4]
  assign io_in_instrctrs_19_cycs = cycles_x723_outr_Foreach_io_count; // @[Ledger.scala 293:21:@80305.4]
  assign io_in_instrctrs_19_iters = iters_x723_outr_Foreach_io_count; // @[Ledger.scala 294:22:@80306.4]
  assign io_in_instrctrs_20_cycs = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_20_cycs; // @[Ledger.scala 302:78:@80643.4]
  assign io_in_instrctrs_20_iters = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_20_iters; // @[Ledger.scala 302:78:@80642.4]
  assign io_in_instrctrs_21_cycs = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_21_cycs; // @[Ledger.scala 302:78:@80647.4]
  assign io_in_instrctrs_21_iters = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_21_iters; // @[Ledger.scala 302:78:@80646.4]
  assign io_in_instrctrs_21_stalls = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_21_stalls; // @[Ledger.scala 302:78:@80645.4]
  assign io_in_instrctrs_21_idles = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_21_idles; // @[Ledger.scala 302:78:@80644.4]
  assign io_in_instrctrs_22_cycs = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_22_cycs; // @[Ledger.scala 302:78:@80651.4]
  assign io_in_instrctrs_22_iters = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_22_iters; // @[Ledger.scala 302:78:@80650.4]
  assign io_in_instrctrs_22_stalls = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_22_stalls; // @[Ledger.scala 302:78:@80649.4]
  assign io_in_instrctrs_22_idles = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_instrctrs_22_idles; // @[Ledger.scala 302:78:@80648.4]
  assign io_in_instrctrs_23_cycs = x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_instrctrs_23_cycs; // @[Ledger.scala 302:78:@80953.4]
  assign io_in_instrctrs_23_iters = x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_instrctrs_23_iters; // @[Ledger.scala 302:78:@80952.4]
  assign io_in_instrctrs_23_stalls = x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_instrctrs_23_stalls; // @[Ledger.scala 302:78:@80951.4]
  assign io_in_instrctrs_23_idles = x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_instrctrs_23_idles; // @[Ledger.scala 302:78:@80950.4]
  assign io_sigsOut_smDoneIn_0 = x718_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 155:56:@80454.4]
  assign io_sigsOut_smDoneIn_1 = x722_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 155:56:@80801.4]
  assign io_sigsOut_smMaskIn_0 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[SpatialBlocks.scala 155:86:@80455.4]
  assign io_sigsOut_smMaskIn_1 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[SpatialBlocks.scala 155:86:@80802.4]
  assign cycles_x723_outr_Foreach_clock = clock; // @[:@80294.4]
  assign cycles_x723_outr_Foreach_reset = reset; // @[:@80295.4]
  assign cycles_x723_outr_Foreach_io_enable = io_sigsIn_baseEn; // @[sm_x723_outr_Foreach.scala 80:42:@80299.4]
  assign iters_x723_outr_Foreach_clock = clock; // @[:@80297.4]
  assign iters_x723_outr_Foreach_reset = reset; // @[:@80298.4]
  assign iters_x723_outr_Foreach_io_enable = io_sigsIn_done & _T_287; // @[sm_x723_outr_Foreach.scala 81:41:@80304.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@80316.4]
  assign x718_outr_UnitPipe_sm_clock = clock; // @[:@80364.4]
  assign x718_outr_UnitPipe_sm_reset = reset; // @[:@80365.4]
  assign x718_outr_UnitPipe_sm_io_enable = _T_374 & _T_383; // @[SpatialBlocks.scala 139:18:@80451.4]
  assign x718_outr_UnitPipe_sm_io_ctrDone = x718_outr_UnitPipe_sm_io_ctrInc & _T_359; // @[sm_x723_outr_Foreach.scala 86:40:@80400.4]
  assign x718_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@80453.4]
  assign x718_outr_UnitPipe_sm_io_doneIn_0 = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@80421.4]
  assign x718_outr_UnitPipe_sm_io_doneIn_1 = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:72:@80422.4]
  assign x718_outr_UnitPipe_sm_io_maskIn_0 = 1'h1; // @[SpatialBlocks.scala 131:72:@80423.4]
  assign x718_outr_UnitPipe_sm_io_maskIn_1 = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smMaskIn_1; // @[SpatialBlocks.scala 131:72:@80424.4]
  assign RetimeWrapper_clock = clock; // @[:@80432.4]
  assign RetimeWrapper_reset = reset; // @[:@80433.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@80435.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@80434.4]
  assign RetimeWrapper_1_clock = clock; // @[:@80440.4]
  assign RetimeWrapper_1_reset = reset; // @[:@80441.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@80443.4]
  assign RetimeWrapper_1_io_in = x718_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@80442.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_clock = clock; // @[:@80469.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_reset = reset; // @[:@80470.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_ready = io_in_x670_ready; // @[sm_x718_outr_UnitPipe.scala 61:23:@80627.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_ready = io_in_x669_ready; // @[sm_x718_outr_UnitPipe.scala 62:23:@80631.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_b674_number = __io_result; // @[sm_x718_outr_UnitPipe.scala 63:23:@80632.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x470_out_host_number = io_in_x470_out_host_number; // @[sm_x718_outr_UnitPipe.scala 65:32:@80634.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_output_0 = io_in_x539_out_sram_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@80635.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_done = x718_outr_UnitPipe_sm_io_done; // @[sm_x718_outr_UnitPipe.scala 125:22:@80674.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_baseEn = _T_374 & _T_383; // @[sm_x718_outr_UnitPipe.scala 125:22:@80666.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x718_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x718_outr_UnitPipe.scala 125:22:@80662.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x718_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x718_outr_UnitPipe.scala 125:22:@80663.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x718_outr_UnitPipe_sm_io_childAck_0; // @[sm_x718_outr_UnitPipe.scala 125:22:@80658.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x718_outr_UnitPipe_sm_io_childAck_1; // @[sm_x718_outr_UnitPipe.scala 125:22:@80659.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x718_outr_UnitPipe.scala 124:18:@80652.4]
  assign x722_inr_UnitPipe_sm_clock = clock; // @[:@80721.4]
  assign x722_inr_UnitPipe_sm_reset = reset; // @[:@80722.4]
  assign x722_inr_UnitPipe_sm_io_enable = x722_inr_UnitPipe_mySignalsIn_baseEn & x722_inr_UnitPipe_mySignalsIn_forwardpressure; // @[SpatialBlocks.scala 139:18:@80798.4]
  assign x722_inr_UnitPipe_sm_io_ctrDone = x722_inr_UnitPipe_sm_io_ctrInc & _T_454; // @[sm_x723_outr_Foreach.scala 95:39:@80752.4]
  assign x722_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 141:21:@80800.4]
  assign x722_inr_UnitPipe_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@80772.4]
  assign x722_inr_UnitPipe_sm_io_break = 1'h0; // @[sm_x723_outr_Foreach.scala 99:37:@80759.4]
  assign RetimeWrapper_2_clock = clock; // @[:@80779.4]
  assign RetimeWrapper_2_reset = reset; // @[:@80780.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@80782.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@80781.4]
  assign RetimeWrapper_3_clock = clock; // @[:@80787.4]
  assign RetimeWrapper_3_reset = reset; // @[:@80788.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@80790.4]
  assign RetimeWrapper_3_io_in = x722_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@80789.4]
  assign x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_clock = clock; // @[:@80816.4]
  assign x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_reset = reset; // @[:@80817.4]
  assign x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_x671_valid = io_in_x671_valid; // @[sm_x722_inr_UnitPipe.scala 51:23:@80948.4]
  assign x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_sigsIn_done = x722_inr_UnitPipe_sm_io_done; // @[sm_x722_inr_UnitPipe.scala 82:22:@80973.4]
  assign x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x722_inr_UnitPipe_sm_io_datapathEn & b675; // @[sm_x722_inr_UnitPipe.scala 82:22:@80966.4]
  assign x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_sigsIn_baseEn = _T_468 & _T_477; // @[sm_x722_inr_UnitPipe.scala 82:22:@80965.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_287 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_359 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_454 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_287 <= 1'h0;
    end else begin
      _T_287 <= _T_284;
    end
    if (reset) begin
      _T_359 <= 1'h0;
    end else begin
      _T_359 <= _T_356;
    end
    if (reset) begin
      _T_454 <= 1'h0;
    end else begin
      _T_454 <= _T_451;
    end
  end
endmodule
module x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1( // @[:@80982.2]
  input         clock, // @[:@80983.4]
  input         reset, // @[:@80984.4]
  input         io_in_x670_ready, // @[:@80985.4]
  output        io_in_x670_valid, // @[:@80985.4]
  output [31:0] io_in_x670_bits_wdata_0, // @[:@80985.4]
  output        io_in_x670_bits_wstrb, // @[:@80985.4]
  input         io_in_x669_ready, // @[:@80985.4]
  output        io_in_x669_valid, // @[:@80985.4]
  output [63:0] io_in_x669_bits_addr, // @[:@80985.4]
  output [31:0] io_in_x669_bits_size, // @[:@80985.4]
  input  [63:0] io_in_x470_out_host_number, // @[:@80985.4]
  output [8:0]  io_in_x539_out_sram_0_rPort_0_ofs_0, // @[:@80985.4]
  output        io_in_x539_out_sram_0_rPort_0_en_0, // @[:@80985.4]
  output        io_in_x539_out_sram_0_rPort_0_backpressure, // @[:@80985.4]
  input  [31:0] io_in_x539_out_sram_0_rPort_0_output_0, // @[:@80985.4]
  output        io_in_x671_ready, // @[:@80985.4]
  input         io_in_x671_valid, // @[:@80985.4]
  output [63:0] io_in_instrctrs_18_cycs, // @[:@80985.4]
  output [63:0] io_in_instrctrs_18_iters, // @[:@80985.4]
  output [63:0] io_in_instrctrs_19_cycs, // @[:@80985.4]
  output [63:0] io_in_instrctrs_19_iters, // @[:@80985.4]
  output [63:0] io_in_instrctrs_20_cycs, // @[:@80985.4]
  output [63:0] io_in_instrctrs_20_iters, // @[:@80985.4]
  output [63:0] io_in_instrctrs_21_cycs, // @[:@80985.4]
  output [63:0] io_in_instrctrs_21_iters, // @[:@80985.4]
  output [63:0] io_in_instrctrs_21_stalls, // @[:@80985.4]
  output [63:0] io_in_instrctrs_21_idles, // @[:@80985.4]
  output [63:0] io_in_instrctrs_22_cycs, // @[:@80985.4]
  output [63:0] io_in_instrctrs_22_iters, // @[:@80985.4]
  output [63:0] io_in_instrctrs_22_stalls, // @[:@80985.4]
  output [63:0] io_in_instrctrs_22_idles, // @[:@80985.4]
  output [63:0] io_in_instrctrs_23_cycs, // @[:@80985.4]
  output [63:0] io_in_instrctrs_23_iters, // @[:@80985.4]
  output [63:0] io_in_instrctrs_23_stalls, // @[:@80985.4]
  output [63:0] io_in_instrctrs_23_idles, // @[:@80985.4]
  input         io_sigsIn_done, // @[:@80985.4]
  input         io_sigsIn_baseEn, // @[:@80985.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@80985.4]
  input         io_sigsIn_smChildAcks_0, // @[:@80985.4]
  output        io_sigsOut_smDoneIn_0, // @[:@80985.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@80985.4]
  input         io_rr // @[:@80985.4]
);
  wire  cycles_x724_outr_UnitPipe_DenseTransfer_clock; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 78:59:@81104.4]
  wire  cycles_x724_outr_UnitPipe_DenseTransfer_reset; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 78:59:@81104.4]
  wire  cycles_x724_outr_UnitPipe_DenseTransfer_io_enable; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 78:59:@81104.4]
  wire [63:0] cycles_x724_outr_UnitPipe_DenseTransfer_io_count; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 78:59:@81104.4]
  wire  iters_x724_outr_UnitPipe_DenseTransfer_clock; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 79:58:@81107.4]
  wire  iters_x724_outr_UnitPipe_DenseTransfer_reset; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 79:58:@81107.4]
  wire  iters_x724_outr_UnitPipe_DenseTransfer_io_enable; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 79:58:@81107.4]
  wire [63:0] iters_x724_outr_UnitPipe_DenseTransfer_io_count; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 79:58:@81107.4]
  wire  x673_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@81120.4]
  wire  x673_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@81120.4]
  wire  x673_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@81120.4]
  wire  x673_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@81120.4]
  wire [8:0] x673_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@81120.4]
  wire  x673_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@81120.4]
  wire  x673_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@81120.4]
  wire  x723_outr_Foreach_sm_clock; // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
  wire  x723_outr_Foreach_sm_reset; // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
  wire  x723_outr_Foreach_sm_io_enable; // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
  wire  x723_outr_Foreach_sm_io_done; // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
  wire  x723_outr_Foreach_sm_io_ctrDone; // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
  wire  x723_outr_Foreach_sm_io_ctrInc; // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
  wire  x723_outr_Foreach_sm_io_ctrRst; // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
  wire  x723_outr_Foreach_sm_io_parentAck; // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
  wire  x723_outr_Foreach_sm_io_doneIn_0; // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
  wire  x723_outr_Foreach_sm_io_doneIn_1; // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
  wire  x723_outr_Foreach_sm_io_maskIn_0; // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
  wire  x723_outr_Foreach_sm_io_maskIn_1; // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
  wire  x723_outr_Foreach_sm_io_enableOut_0; // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
  wire  x723_outr_Foreach_sm_io_enableOut_1; // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
  wire  x723_outr_Foreach_sm_io_childAck_0; // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
  wire  x723_outr_Foreach_sm_io_childAck_1; // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@81212.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@81212.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@81212.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@81212.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@81212.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@81257.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@81257.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@81257.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@81257.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@81257.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@81265.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@81265.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@81265.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@81265.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@81265.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_clock; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_reset; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_ready; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_valid; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [31:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_bits_wdata_0; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_bits_wstrb; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_ready; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_valid; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_bits_addr; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [31:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_bits_size; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x470_out_host_number; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [8:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_en_0; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [31:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_output_0; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x671_ready; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x671_valid; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_19_cycs; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_19_iters; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_20_cycs; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_20_iters; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_21_cycs; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_21_iters; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_21_stalls; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_21_idles; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_22_cycs; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_22_iters; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_22_stalls; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_22_idles; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_23_cycs; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_23_iters; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_23_stalls; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_23_idles; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_done; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire [31:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_rr; // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
  wire  _T_284; // @[package.scala 100:49:@81111.4]
  reg  _T_287; // @[package.scala 48:56:@81112.4]
  reg [31:0] _RAND_0;
  wire  _T_353; // @[package.scala 96:25:@81217.4 package.scala 96:25:@81218.4]
  wire  _T_370; // @[package.scala 96:25:@81262.4 package.scala 96:25:@81263.4]
  wire  _T_376; // @[package.scala 96:25:@81270.4 package.scala 96:25:@81271.4]
  wire  _T_379; // @[SpatialBlocks.scala 137:99:@81273.4]
  InstrumentationCounter cycles_x724_outr_UnitPipe_DenseTransfer ( // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 78:59:@81104.4]
    .clock(cycles_x724_outr_UnitPipe_DenseTransfer_clock),
    .reset(cycles_x724_outr_UnitPipe_DenseTransfer_reset),
    .io_enable(cycles_x724_outr_UnitPipe_DenseTransfer_io_enable),
    .io_count(cycles_x724_outr_UnitPipe_DenseTransfer_io_count)
  );
  InstrumentationCounter iters_x724_outr_UnitPipe_DenseTransfer ( // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 79:58:@81107.4]
    .clock(iters_x724_outr_UnitPipe_DenseTransfer_clock),
    .reset(iters_x724_outr_UnitPipe_DenseTransfer_reset),
    .io_enable(iters_x724_outr_UnitPipe_DenseTransfer_io_enable),
    .io_count(iters_x724_outr_UnitPipe_DenseTransfer_io_count)
  );
  x478_ctrchain x673_ctrchain ( // @[SpatialBlocks.scala 37:22:@81120.4]
    .clock(x673_ctrchain_clock),
    .reset(x673_ctrchain_reset),
    .io_input_reset(x673_ctrchain_io_input_reset),
    .io_input_enable(x673_ctrchain_io_input_enable),
    .io_output_counts_0(x673_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x673_ctrchain_io_output_oobs_0),
    .io_output_done(x673_ctrchain_io_output_done)
  );
  x537_outr_Foreach_sm x723_outr_Foreach_sm ( // @[sm_x723_outr_Foreach.scala 36:18:@81178.4]
    .clock(x723_outr_Foreach_sm_clock),
    .reset(x723_outr_Foreach_sm_reset),
    .io_enable(x723_outr_Foreach_sm_io_enable),
    .io_done(x723_outr_Foreach_sm_io_done),
    .io_ctrDone(x723_outr_Foreach_sm_io_ctrDone),
    .io_ctrInc(x723_outr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x723_outr_Foreach_sm_io_ctrRst),
    .io_parentAck(x723_outr_Foreach_sm_io_parentAck),
    .io_doneIn_0(x723_outr_Foreach_sm_io_doneIn_0),
    .io_doneIn_1(x723_outr_Foreach_sm_io_doneIn_1),
    .io_maskIn_0(x723_outr_Foreach_sm_io_maskIn_0),
    .io_maskIn_1(x723_outr_Foreach_sm_io_maskIn_1),
    .io_enableOut_0(x723_outr_Foreach_sm_io_enableOut_0),
    .io_enableOut_1(x723_outr_Foreach_sm_io_enableOut_1),
    .io_childAck_0(x723_outr_Foreach_sm_io_childAck_0),
    .io_childAck_1(x723_outr_Foreach_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@81212.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@81257.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@81265.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1 x723_outr_Foreach_kernelx723_outr_Foreach_concrete1 ( // @[sm_x723_outr_Foreach.scala 104:24:@81300.4]
    .clock(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_clock),
    .reset(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_reset),
    .io_in_x670_ready(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_ready),
    .io_in_x670_valid(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_valid),
    .io_in_x670_bits_wdata_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_bits_wdata_0),
    .io_in_x670_bits_wstrb(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_bits_wstrb),
    .io_in_x669_ready(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_ready),
    .io_in_x669_valid(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_valid),
    .io_in_x669_bits_addr(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_bits_addr),
    .io_in_x669_bits_size(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_bits_size),
    .io_in_x470_out_host_number(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x470_out_host_number),
    .io_in_x539_out_sram_0_rPort_0_ofs_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0),
    .io_in_x539_out_sram_0_rPort_0_en_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_en_0),
    .io_in_x539_out_sram_0_rPort_0_backpressure(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure),
    .io_in_x539_out_sram_0_rPort_0_output_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_output_0),
    .io_in_x671_ready(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x671_ready),
    .io_in_x671_valid(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x671_valid),
    .io_in_instrctrs_19_cycs(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_19_cycs),
    .io_in_instrctrs_19_iters(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_19_iters),
    .io_in_instrctrs_20_cycs(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_20_cycs),
    .io_in_instrctrs_20_iters(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_20_iters),
    .io_in_instrctrs_21_cycs(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_21_cycs),
    .io_in_instrctrs_21_iters(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_21_iters),
    .io_in_instrctrs_21_stalls(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_21_stalls),
    .io_in_instrctrs_21_idles(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_21_idles),
    .io_in_instrctrs_22_cycs(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_22_cycs),
    .io_in_instrctrs_22_iters(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_22_iters),
    .io_in_instrctrs_22_stalls(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_22_stalls),
    .io_in_instrctrs_22_idles(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_22_idles),
    .io_in_instrctrs_23_cycs(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_23_cycs),
    .io_in_instrctrs_23_iters(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_23_iters),
    .io_in_instrctrs_23_stalls(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_23_stalls),
    .io_in_instrctrs_23_idles(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_23_idles),
    .io_sigsIn_done(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smEnableOuts_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsOut_smDoneIn_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smMaskIn_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0),
    .io_sigsOut_smMaskIn_1(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1),
    .io_rr(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_rr)
  );
  assign _T_284 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@81111.4]
  assign _T_353 = RetimeWrapper_io_out; // @[package.scala 96:25:@81217.4 package.scala 96:25:@81218.4]
  assign _T_370 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@81262.4 package.scala 96:25:@81263.4]
  assign _T_376 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@81270.4 package.scala 96:25:@81271.4]
  assign _T_379 = ~ _T_376; // @[SpatialBlocks.scala 137:99:@81273.4]
  assign io_in_x670_valid = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_valid; // @[sm_x723_outr_Foreach.scala 59:23:@81459.4]
  assign io_in_x670_bits_wdata_0 = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_bits_wdata_0; // @[sm_x723_outr_Foreach.scala 59:23:@81458.4]
  assign io_in_x670_bits_wstrb = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_bits_wstrb; // @[sm_x723_outr_Foreach.scala 59:23:@81457.4]
  assign io_in_x669_valid = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_valid; // @[sm_x723_outr_Foreach.scala 60:23:@81463.4]
  assign io_in_x669_bits_addr = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_bits_addr; // @[sm_x723_outr_Foreach.scala 60:23:@81462.4]
  assign io_in_x669_bits_size = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_bits_size; // @[sm_x723_outr_Foreach.scala 60:23:@81461.4]
  assign io_in_x539_out_sram_0_rPort_0_ofs_0 = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@81469.4]
  assign io_in_x539_out_sram_0_rPort_0_en_0 = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@81468.4]
  assign io_in_x539_out_sram_0_rPort_0_backpressure = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@81467.4]
  assign io_in_x671_ready = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x671_ready; // @[sm_x723_outr_Foreach.scala 63:23:@81473.4]
  assign io_in_instrctrs_18_cycs = cycles_x724_outr_UnitPipe_DenseTransfer_io_count; // @[Ledger.scala 293:21:@81116.4]
  assign io_in_instrctrs_18_iters = iters_x724_outr_UnitPipe_DenseTransfer_io_count; // @[Ledger.scala 294:22:@81117.4]
  assign io_in_instrctrs_19_cycs = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_19_cycs; // @[Ledger.scala 302:78:@81477.4]
  assign io_in_instrctrs_19_iters = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_19_iters; // @[Ledger.scala 302:78:@81476.4]
  assign io_in_instrctrs_20_cycs = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_20_cycs; // @[Ledger.scala 302:78:@81481.4]
  assign io_in_instrctrs_20_iters = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_20_iters; // @[Ledger.scala 302:78:@81480.4]
  assign io_in_instrctrs_21_cycs = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_21_cycs; // @[Ledger.scala 302:78:@81485.4]
  assign io_in_instrctrs_21_iters = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_21_iters; // @[Ledger.scala 302:78:@81484.4]
  assign io_in_instrctrs_21_stalls = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_21_stalls; // @[Ledger.scala 302:78:@81483.4]
  assign io_in_instrctrs_21_idles = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_21_idles; // @[Ledger.scala 302:78:@81482.4]
  assign io_in_instrctrs_22_cycs = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_22_cycs; // @[Ledger.scala 302:78:@81489.4]
  assign io_in_instrctrs_22_iters = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_22_iters; // @[Ledger.scala 302:78:@81488.4]
  assign io_in_instrctrs_22_stalls = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_22_stalls; // @[Ledger.scala 302:78:@81487.4]
  assign io_in_instrctrs_22_idles = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_22_idles; // @[Ledger.scala 302:78:@81486.4]
  assign io_in_instrctrs_23_cycs = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_23_cycs; // @[Ledger.scala 302:78:@81493.4]
  assign io_in_instrctrs_23_iters = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_23_iters; // @[Ledger.scala 302:78:@81492.4]
  assign io_in_instrctrs_23_stalls = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_23_stalls; // @[Ledger.scala 302:78:@81491.4]
  assign io_in_instrctrs_23_idles = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_instrctrs_23_idles; // @[Ledger.scala 302:78:@81490.4]
  assign io_sigsOut_smDoneIn_0 = x723_outr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@81280.4]
  assign io_sigsOut_smCtrCopyDone_0 = x723_outr_Foreach_sm_io_done; // @[SpatialBlocks.scala 170:140:@81299.4]
  assign cycles_x724_outr_UnitPipe_DenseTransfer_clock = clock; // @[:@81105.4]
  assign cycles_x724_outr_UnitPipe_DenseTransfer_reset = reset; // @[:@81106.4]
  assign cycles_x724_outr_UnitPipe_DenseTransfer_io_enable = io_sigsIn_baseEn; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 80:57:@81110.4]
  assign iters_x724_outr_UnitPipe_DenseTransfer_clock = clock; // @[:@81108.4]
  assign iters_x724_outr_UnitPipe_DenseTransfer_reset = reset; // @[:@81109.4]
  assign iters_x724_outr_UnitPipe_DenseTransfer_io_enable = io_sigsIn_done & _T_287; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 81:56:@81115.4]
  assign x673_ctrchain_clock = clock; // @[:@81121.4]
  assign x673_ctrchain_reset = reset; // @[:@81122.4]
  assign x673_ctrchain_io_input_reset = x723_outr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@81298.4]
  assign x673_ctrchain_io_input_enable = x723_outr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 158:42:@81297.4]
  assign x723_outr_Foreach_sm_clock = clock; // @[:@81179.4]
  assign x723_outr_Foreach_sm_reset = reset; // @[:@81180.4]
  assign x723_outr_Foreach_sm_io_enable = _T_370 & _T_379; // @[SpatialBlocks.scala 139:18:@81277.4]
  assign x723_outr_Foreach_sm_io_ctrDone = io_rr ? _T_353 : 1'h0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 88:39:@81220.4]
  assign x723_outr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@81279.4]
  assign x723_outr_Foreach_sm_io_doneIn_0 = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@81247.4]
  assign x723_outr_Foreach_sm_io_doneIn_1 = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:72:@81248.4]
  assign x723_outr_Foreach_sm_io_maskIn_0 = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0; // @[SpatialBlocks.scala 131:72:@81249.4]
  assign x723_outr_Foreach_sm_io_maskIn_1 = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1; // @[SpatialBlocks.scala 131:72:@81250.4]
  assign RetimeWrapper_clock = clock; // @[:@81213.4]
  assign RetimeWrapper_reset = reset; // @[:@81214.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@81216.4]
  assign RetimeWrapper_io_in = x673_ctrchain_io_output_done; // @[package.scala 94:16:@81215.4]
  assign RetimeWrapper_1_clock = clock; // @[:@81258.4]
  assign RetimeWrapper_1_reset = reset; // @[:@81259.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@81261.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@81260.4]
  assign RetimeWrapper_2_clock = clock; // @[:@81266.4]
  assign RetimeWrapper_2_reset = reset; // @[:@81267.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@81269.4]
  assign RetimeWrapper_2_io_in = x723_outr_Foreach_sm_io_done; // @[package.scala 94:16:@81268.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_clock = clock; // @[:@81301.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_reset = reset; // @[:@81302.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_ready = io_in_x670_ready; // @[sm_x723_outr_Foreach.scala 59:23:@81460.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_ready = io_in_x669_ready; // @[sm_x723_outr_Foreach.scala 60:23:@81464.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x470_out_host_number = io_in_x470_out_host_number; // @[sm_x723_outr_Foreach.scala 61:32:@81465.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_output_0 = io_in_x539_out_sram_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@81466.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x671_valid = io_in_x671_valid; // @[sm_x723_outr_Foreach.scala 63:23:@81472.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_done = x723_outr_Foreach_sm_io_done; // @[sm_x723_outr_Foreach.scala 110:22:@81516.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_baseEn = _T_370 & _T_379; // @[sm_x723_outr_Foreach.scala 110:22:@81508.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0 = x723_outr_Foreach_sm_io_enableOut_0; // @[sm_x723_outr_Foreach.scala 110:22:@81504.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1 = x723_outr_Foreach_sm_io_enableOut_1; // @[sm_x723_outr_Foreach.scala 110:22:@81505.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0 = x723_outr_Foreach_sm_io_childAck_0; // @[sm_x723_outr_Foreach.scala 110:22:@81500.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1 = x723_outr_Foreach_sm_io_childAck_1; // @[sm_x723_outr_Foreach.scala 110:22:@81501.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{23{x673_ctrchain_io_output_counts_0[8]}},x673_ctrchain_io_output_counts_0}; // @[sm_x723_outr_Foreach.scala 110:22:@81499.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x673_ctrchain_io_output_oobs_0; // @[sm_x723_outr_Foreach.scala 110:22:@81498.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_rr = io_rr; // @[sm_x723_outr_Foreach.scala 109:18:@81494.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_287 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_287 <= 1'h0;
    end else begin
      _T_287 <= _T_284;
    end
  end
endmodule
module RootController_kernelRootController_concrete1( // @[:@81527.2]
  input         clock, // @[:@81528.4]
  input         reset, // @[:@81529.4]
  input  [63:0] io_in_x468_A_dram_number, // @[:@81530.4]
  input         io_in_x670_ready, // @[:@81530.4]
  output        io_in_x670_valid, // @[:@81530.4]
  output [31:0] io_in_x670_bits_wdata_0, // @[:@81530.4]
  output        io_in_x670_bits_wstrb, // @[:@81530.4]
  input         io_in_x669_ready, // @[:@81530.4]
  output        io_in_x669_valid, // @[:@81530.4]
  output [63:0] io_in_x669_bits_addr, // @[:@81530.4]
  output [31:0] io_in_x669_bits_size, // @[:@81530.4]
  output        io_in_x476_ready, // @[:@81530.4]
  input         io_in_x476_valid, // @[:@81530.4]
  input  [31:0] io_in_x476_bits_rdata_0, // @[:@81530.4]
  input  [63:0] io_in_x470_out_host_number, // @[:@81530.4]
  output        io_in_x671_ready, // @[:@81530.4]
  input         io_in_x671_valid, // @[:@81530.4]
  input         io_in_x474_ready, // @[:@81530.4]
  output        io_in_x474_valid, // @[:@81530.4]
  output [63:0] io_in_x474_bits_addr, // @[:@81530.4]
  output [31:0] io_in_x474_bits_size, // @[:@81530.4]
  output [63:0] io_in_instrctrs_0_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_0_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_1_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_1_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_2_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_2_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_2_stalls, // @[:@81530.4]
  output [63:0] io_in_instrctrs_2_idles, // @[:@81530.4]
  output [63:0] io_in_instrctrs_3_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_3_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_4_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_4_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_4_stalls, // @[:@81530.4]
  output [63:0] io_in_instrctrs_4_idles, // @[:@81530.4]
  output [63:0] io_in_instrctrs_5_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_5_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_5_stalls, // @[:@81530.4]
  output [63:0] io_in_instrctrs_5_idles, // @[:@81530.4]
  output [63:0] io_in_instrctrs_6_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_6_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_7_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_7_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_8_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_8_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_9_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_9_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_10_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_10_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_11_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_11_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_12_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_12_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_13_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_13_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_14_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_14_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_15_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_15_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_16_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_16_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_17_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_17_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_18_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_18_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_19_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_19_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_20_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_20_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_21_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_21_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_21_stalls, // @[:@81530.4]
  output [63:0] io_in_instrctrs_21_idles, // @[:@81530.4]
  output [63:0] io_in_instrctrs_22_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_22_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_22_stalls, // @[:@81530.4]
  output [63:0] io_in_instrctrs_22_idles, // @[:@81530.4]
  output [63:0] io_in_instrctrs_23_cycs, // @[:@81530.4]
  output [63:0] io_in_instrctrs_23_iters, // @[:@81530.4]
  output [63:0] io_in_instrctrs_23_stalls, // @[:@81530.4]
  output [63:0] io_in_instrctrs_23_idles, // @[:@81530.4]
  input         io_sigsIn_done, // @[:@81530.4]
  input         io_sigsIn_baseEn, // @[:@81530.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@81530.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@81530.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@81530.4]
  input         io_sigsIn_smChildAcks_0, // @[:@81530.4]
  input         io_sigsIn_smChildAcks_1, // @[:@81530.4]
  input         io_sigsIn_smChildAcks_2, // @[:@81530.4]
  output        io_sigsOut_smDoneIn_0, // @[:@81530.4]
  output        io_sigsOut_smDoneIn_1, // @[:@81530.4]
  output        io_sigsOut_smDoneIn_2, // @[:@81530.4]
  input         io_rr // @[:@81530.4]
);
  wire  cycles_RootController_clock; // @[sm_RootController.scala 86:41:@81640.4]
  wire  cycles_RootController_reset; // @[sm_RootController.scala 86:41:@81640.4]
  wire  cycles_RootController_io_enable; // @[sm_RootController.scala 86:41:@81640.4]
  wire [63:0] cycles_RootController_io_count; // @[sm_RootController.scala 86:41:@81640.4]
  wire  iters_RootController_clock; // @[sm_RootController.scala 87:40:@81643.4]
  wire  iters_RootController_reset; // @[sm_RootController.scala 87:40:@81643.4]
  wire  iters_RootController_io_enable; // @[sm_RootController.scala 87:40:@81643.4]
  wire [63:0] iters_RootController_io_count; // @[sm_RootController.scala 87:40:@81643.4]
  wire  x471_A_sram_0_clock; // @[m_x471_A_sram_0.scala 27:22:@81656.4]
  wire  x471_A_sram_0_reset; // @[m_x471_A_sram_0.scala 27:22:@81656.4]
  wire [8:0] x471_A_sram_0_io_rPort_0_ofs_0; // @[m_x471_A_sram_0.scala 27:22:@81656.4]
  wire  x471_A_sram_0_io_rPort_0_en_0; // @[m_x471_A_sram_0.scala 27:22:@81656.4]
  wire  x471_A_sram_0_io_rPort_0_backpressure; // @[m_x471_A_sram_0.scala 27:22:@81656.4]
  wire [31:0] x471_A_sram_0_io_rPort_0_output_0; // @[m_x471_A_sram_0.scala 27:22:@81656.4]
  wire [8:0] x471_A_sram_0_io_wPort_0_ofs_0; // @[m_x471_A_sram_0.scala 27:22:@81656.4]
  wire [31:0] x471_A_sram_0_io_wPort_0_data_0; // @[m_x471_A_sram_0.scala 27:22:@81656.4]
  wire  x471_A_sram_0_io_wPort_0_en_0; // @[m_x471_A_sram_0.scala 27:22:@81656.4]
  wire  x472_A_sram_1_clock; // @[m_x472_A_sram_1.scala 27:22:@81673.4]
  wire  x472_A_sram_1_reset; // @[m_x472_A_sram_1.scala 27:22:@81673.4]
  wire [8:0] x472_A_sram_1_io_rPort_0_ofs_0; // @[m_x472_A_sram_1.scala 27:22:@81673.4]
  wire  x472_A_sram_1_io_rPort_0_en_0; // @[m_x472_A_sram_1.scala 27:22:@81673.4]
  wire  x472_A_sram_1_io_rPort_0_backpressure; // @[m_x472_A_sram_1.scala 27:22:@81673.4]
  wire [31:0] x472_A_sram_1_io_rPort_0_output_0; // @[m_x472_A_sram_1.scala 27:22:@81673.4]
  wire [8:0] x472_A_sram_1_io_wPort_0_ofs_0; // @[m_x472_A_sram_1.scala 27:22:@81673.4]
  wire [31:0] x472_A_sram_1_io_wPort_0_data_0; // @[m_x472_A_sram_1.scala 27:22:@81673.4]
  wire  x472_A_sram_1_io_wPort_0_en_0; // @[m_x472_A_sram_1.scala 27:22:@81673.4]
  wire  x473_A_sram_2_clock; // @[m_x473_A_sram_2.scala 27:22:@81690.4]
  wire  x473_A_sram_2_reset; // @[m_x473_A_sram_2.scala 27:22:@81690.4]
  wire [8:0] x473_A_sram_2_io_rPort_0_ofs_0; // @[m_x473_A_sram_2.scala 27:22:@81690.4]
  wire  x473_A_sram_2_io_rPort_0_en_0; // @[m_x473_A_sram_2.scala 27:22:@81690.4]
  wire  x473_A_sram_2_io_rPort_0_backpressure; // @[m_x473_A_sram_2.scala 27:22:@81690.4]
  wire [31:0] x473_A_sram_2_io_rPort_0_output_0; // @[m_x473_A_sram_2.scala 27:22:@81690.4]
  wire [8:0] x473_A_sram_2_io_wPort_0_ofs_0; // @[m_x473_A_sram_2.scala 27:22:@81690.4]
  wire [31:0] x473_A_sram_2_io_wPort_0_data_0; // @[m_x473_A_sram_2.scala 27:22:@81690.4]
  wire  x473_A_sram_2_io_wPort_0_en_0; // @[m_x473_A_sram_2.scala 27:22:@81690.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_clock; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@81755.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_reset; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@81755.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_enable; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@81755.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_done; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@81755.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_parentAck; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@81755.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_doneIn_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@81755.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_doneIn_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@81755.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_enableOut_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@81755.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_enableOut_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@81755.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_childAck_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@81755.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_childAck_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@81755.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@81755.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@81755.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@81818.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@81818.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@81818.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@81818.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@81818.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@81826.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@81826.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@81826.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@81826.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@81826.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_clock; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_reset; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x468_A_dram_number; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [8:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [31:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_data_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_en_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [8:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [31:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_data_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_en_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_ready; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_valid; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [31:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_bits_rdata_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [8:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [31:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_data_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_en_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_ready; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_valid; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_bits_addr; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [31:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_bits_size; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_1_cycs; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_1_iters; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_2_cycs; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_2_iters; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_2_stalls; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_2_idles; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_3_cycs; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_3_iters; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_4_cycs; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_4_iters; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_4_stalls; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_4_idles; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_5_cycs; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_5_iters; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_5_stalls; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_5_idles; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_done; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_baseEn; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_rr; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
  wire  x539_out_sram_0_clock; // @[m_x539_out_sram_0.scala 27:22:@82131.4]
  wire  x539_out_sram_0_reset; // @[m_x539_out_sram_0.scala 27:22:@82131.4]
  wire [8:0] x539_out_sram_0_io_rPort_0_ofs_0; // @[m_x539_out_sram_0.scala 27:22:@82131.4]
  wire  x539_out_sram_0_io_rPort_0_en_0; // @[m_x539_out_sram_0.scala 27:22:@82131.4]
  wire  x539_out_sram_0_io_rPort_0_backpressure; // @[m_x539_out_sram_0.scala 27:22:@82131.4]
  wire [31:0] x539_out_sram_0_io_rPort_0_output_0; // @[m_x539_out_sram_0.scala 27:22:@82131.4]
  wire [8:0] x539_out_sram_0_io_wPort_0_ofs_0; // @[m_x539_out_sram_0.scala 27:22:@82131.4]
  wire [31:0] x539_out_sram_0_io_wPort_0_data_0; // @[m_x539_out_sram_0.scala 27:22:@82131.4]
  wire  x539_out_sram_0_io_wPort_0_en_0; // @[m_x539_out_sram_0.scala 27:22:@82131.4]
  wire  x541_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@82148.4]
  wire  x541_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@82148.4]
  wire  x541_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@82148.4]
  wire  x541_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@82148.4]
  wire [8:0] x541_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@82148.4]
  wire  x541_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@82148.4]
  wire  x541_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@82148.4]
  wire  x668_outr_Foreach_sm_clock; // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
  wire  x668_outr_Foreach_sm_reset; // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
  wire  x668_outr_Foreach_sm_io_enable; // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
  wire  x668_outr_Foreach_sm_io_done; // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
  wire  x668_outr_Foreach_sm_io_ctrDone; // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
  wire  x668_outr_Foreach_sm_io_ctrInc; // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
  wire  x668_outr_Foreach_sm_io_ctrRst; // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
  wire  x668_outr_Foreach_sm_io_parentAck; // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
  wire  x668_outr_Foreach_sm_io_doneIn_0; // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
  wire  x668_outr_Foreach_sm_io_doneIn_1; // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
  wire  x668_outr_Foreach_sm_io_maskIn_0; // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
  wire  x668_outr_Foreach_sm_io_maskIn_1; // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
  wire  x668_outr_Foreach_sm_io_enableOut_0; // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
  wire  x668_outr_Foreach_sm_io_enableOut_1; // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
  wire  x668_outr_Foreach_sm_io_childAck_0; // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
  wire  x668_outr_Foreach_sm_io_childAck_1; // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@82240.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@82240.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@82240.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@82240.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@82240.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@82285.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@82285.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@82285.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@82285.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@82285.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@82293.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@82293.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@82293.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@82293.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@82293.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_clock; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_reset; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [8:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_en_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [31:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_output_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [8:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_en_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [31:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_output_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [8:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_ofs_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_en_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [31:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_output_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [8:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_ofs_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [31:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_data_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_en_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_6_cycs; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_6_iters; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_7_cycs; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_7_iters; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_8_cycs; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_8_iters; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_9_cycs; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_9_iters; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_10_cycs; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_10_iters; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_11_cycs; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_11_iters; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_12_cycs; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_12_iters; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_13_cycs; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_13_iters; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_14_cycs; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_14_iters; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_15_cycs; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_15_iters; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_16_cycs; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_16_iters; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_17_cycs; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [63:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_17_iters; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_done; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire [31:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_rr; // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_clock; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@82649.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_reset; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@82649.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_io_enable; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@82649.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_io_done; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@82649.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_io_parentAck; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@82649.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_io_doneIn_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@82649.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_io_enableOut_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@82649.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_io_childAck_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@82649.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@82649.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@82702.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@82702.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@82702.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@82702.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@82702.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@82710.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@82710.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@82710.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@82710.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@82710.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_clock; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_reset; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_ready; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_valid; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [31:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_bits_wdata_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_bits_wstrb; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_ready; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_valid; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_bits_addr; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [31:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_bits_size; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x470_out_host_number; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [8:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_en_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [31:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_output_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x671_ready; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x671_valid; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_18_cycs; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_18_iters; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_19_cycs; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_19_iters; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_20_cycs; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_20_iters; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_21_cycs; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_21_iters; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_21_stalls; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_21_idles; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_22_cycs; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_22_iters; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_22_stalls; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_22_idles; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_23_cycs; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_23_iters; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_23_stalls; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_23_idles; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_done; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_baseEn; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_rr; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
  wire  _T_190; // @[package.scala 100:49:@81647.4]
  reg  _T_193; // @[package.scala 48:56:@81648.4]
  reg [31:0] _RAND_0;
  wire  _T_277; // @[package.scala 96:25:@81823.4 package.scala 96:25:@81824.4]
  wire  _T_283; // @[package.scala 96:25:@81831.4 package.scala 96:25:@81832.4]
  wire  _T_286; // @[SpatialBlocks.scala 137:99:@81834.4]
  wire  _T_359; // @[package.scala 96:25:@82245.4 package.scala 96:25:@82246.4]
  wire  _T_376; // @[package.scala 96:25:@82290.4 package.scala 96:25:@82291.4]
  wire  _T_382; // @[package.scala 96:25:@82298.4 package.scala 96:25:@82299.4]
  wire  _T_385; // @[SpatialBlocks.scala 137:99:@82301.4]
  wire  _T_468; // @[package.scala 96:25:@82707.4 package.scala 96:25:@82708.4]
  wire  _T_474; // @[package.scala 96:25:@82715.4 package.scala 96:25:@82716.4]
  wire  _T_477; // @[SpatialBlocks.scala 137:99:@82718.4]
  InstrumentationCounter cycles_RootController ( // @[sm_RootController.scala 86:41:@81640.4]
    .clock(cycles_RootController_clock),
    .reset(cycles_RootController_reset),
    .io_enable(cycles_RootController_io_enable),
    .io_count(cycles_RootController_io_count)
  );
  InstrumentationCounter iters_RootController ( // @[sm_RootController.scala 87:40:@81643.4]
    .clock(iters_RootController_clock),
    .reset(iters_RootController_reset),
    .io_enable(iters_RootController_io_enable),
    .io_count(iters_RootController_io_count)
  );
  x471_A_sram_0 x471_A_sram_0 ( // @[m_x471_A_sram_0.scala 27:22:@81656.4]
    .clock(x471_A_sram_0_clock),
    .reset(x471_A_sram_0_reset),
    .io_rPort_0_ofs_0(x471_A_sram_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x471_A_sram_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x471_A_sram_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x471_A_sram_0_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(x471_A_sram_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x471_A_sram_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x471_A_sram_0_io_wPort_0_en_0)
  );
  x471_A_sram_0 x472_A_sram_1 ( // @[m_x472_A_sram_1.scala 27:22:@81673.4]
    .clock(x472_A_sram_1_clock),
    .reset(x472_A_sram_1_reset),
    .io_rPort_0_ofs_0(x472_A_sram_1_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x472_A_sram_1_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x472_A_sram_1_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x472_A_sram_1_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(x472_A_sram_1_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x472_A_sram_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(x472_A_sram_1_io_wPort_0_en_0)
  );
  x471_A_sram_0 x473_A_sram_2 ( // @[m_x473_A_sram_2.scala 27:22:@81690.4]
    .clock(x473_A_sram_2_clock),
    .reset(x473_A_sram_2_reset),
    .io_rPort_0_ofs_0(x473_A_sram_2_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x473_A_sram_2_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x473_A_sram_2_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x473_A_sram_2_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(x473_A_sram_2_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x473_A_sram_2_io_wPort_0_data_0),
    .io_wPort_0_en_0(x473_A_sram_2_io_wPort_0_en_0)
  );
  x538_outr_UnitPipe_DenseTransfer_sm x538_outr_UnitPipe_DenseTransfer_sm ( // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@81755.4]
    .clock(x538_outr_UnitPipe_DenseTransfer_sm_clock),
    .reset(x538_outr_UnitPipe_DenseTransfer_sm_reset),
    .io_enable(x538_outr_UnitPipe_DenseTransfer_sm_io_enable),
    .io_done(x538_outr_UnitPipe_DenseTransfer_sm_io_done),
    .io_parentAck(x538_outr_UnitPipe_DenseTransfer_sm_io_parentAck),
    .io_doneIn_0(x538_outr_UnitPipe_DenseTransfer_sm_io_doneIn_0),
    .io_doneIn_1(x538_outr_UnitPipe_DenseTransfer_sm_io_doneIn_1),
    .io_enableOut_0(x538_outr_UnitPipe_DenseTransfer_sm_io_enableOut_0),
    .io_enableOut_1(x538_outr_UnitPipe_DenseTransfer_sm_io_enableOut_1),
    .io_childAck_0(x538_outr_UnitPipe_DenseTransfer_sm_io_childAck_0),
    .io_childAck_1(x538_outr_UnitPipe_DenseTransfer_sm_io_childAck_1),
    .io_ctrCopyDone_0(x538_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x538_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@81818.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@81826.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1 x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1 ( // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 114:24:@81857.4]
    .clock(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_clock),
    .reset(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_reset),
    .io_in_x468_A_dram_number(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x468_A_dram_number),
    .io_in_x472_A_sram_1_wPort_0_ofs_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0),
    .io_in_x472_A_sram_1_wPort_0_data_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_data_0),
    .io_in_x472_A_sram_1_wPort_0_en_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_en_0),
    .io_in_x471_A_sram_0_wPort_0_ofs_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0),
    .io_in_x471_A_sram_0_wPort_0_data_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_data_0),
    .io_in_x471_A_sram_0_wPort_0_en_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_en_0),
    .io_in_x476_ready(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_ready),
    .io_in_x476_valid(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_valid),
    .io_in_x476_bits_rdata_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_bits_rdata_0),
    .io_in_x473_A_sram_2_wPort_0_ofs_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0),
    .io_in_x473_A_sram_2_wPort_0_data_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_data_0),
    .io_in_x473_A_sram_2_wPort_0_en_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_en_0),
    .io_in_x474_ready(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_ready),
    .io_in_x474_valid(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_valid),
    .io_in_x474_bits_addr(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_bits_addr),
    .io_in_x474_bits_size(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_bits_size),
    .io_in_instrctrs_1_cycs(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_1_cycs),
    .io_in_instrctrs_1_iters(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_1_iters),
    .io_in_instrctrs_2_cycs(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_2_cycs),
    .io_in_instrctrs_2_iters(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_2_iters),
    .io_in_instrctrs_2_stalls(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_2_stalls),
    .io_in_instrctrs_2_idles(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_2_idles),
    .io_in_instrctrs_3_cycs(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_3_cycs),
    .io_in_instrctrs_3_iters(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_3_iters),
    .io_in_instrctrs_4_cycs(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_4_cycs),
    .io_in_instrctrs_4_iters(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_4_iters),
    .io_in_instrctrs_4_stalls(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_4_stalls),
    .io_in_instrctrs_4_idles(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_4_idles),
    .io_in_instrctrs_5_cycs(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_5_cycs),
    .io_in_instrctrs_5_iters(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_5_iters),
    .io_in_instrctrs_5_stalls(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_5_stalls),
    .io_in_instrctrs_5_idles(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_5_idles),
    .io_sigsIn_done(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smEnableOuts_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_rr)
  );
  x471_A_sram_0 x539_out_sram_0 ( // @[m_x539_out_sram_0.scala 27:22:@82131.4]
    .clock(x539_out_sram_0_clock),
    .reset(x539_out_sram_0_reset),
    .io_rPort_0_ofs_0(x539_out_sram_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x539_out_sram_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x539_out_sram_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x539_out_sram_0_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(x539_out_sram_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x539_out_sram_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x539_out_sram_0_io_wPort_0_en_0)
  );
  x478_ctrchain x541_ctrchain ( // @[SpatialBlocks.scala 37:22:@82148.4]
    .clock(x541_ctrchain_clock),
    .reset(x541_ctrchain_reset),
    .io_input_reset(x541_ctrchain_io_input_reset),
    .io_input_enable(x541_ctrchain_io_input_enable),
    .io_output_counts_0(x541_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x541_ctrchain_io_output_oobs_0),
    .io_output_done(x541_ctrchain_io_output_done)
  );
  x668_outr_Foreach_sm x668_outr_Foreach_sm ( // @[sm_x668_outr_Foreach.scala 32:18:@82206.4]
    .clock(x668_outr_Foreach_sm_clock),
    .reset(x668_outr_Foreach_sm_reset),
    .io_enable(x668_outr_Foreach_sm_io_enable),
    .io_done(x668_outr_Foreach_sm_io_done),
    .io_ctrDone(x668_outr_Foreach_sm_io_ctrDone),
    .io_ctrInc(x668_outr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x668_outr_Foreach_sm_io_ctrRst),
    .io_parentAck(x668_outr_Foreach_sm_io_parentAck),
    .io_doneIn_0(x668_outr_Foreach_sm_io_doneIn_0),
    .io_doneIn_1(x668_outr_Foreach_sm_io_doneIn_1),
    .io_maskIn_0(x668_outr_Foreach_sm_io_maskIn_0),
    .io_maskIn_1(x668_outr_Foreach_sm_io_maskIn_1),
    .io_enableOut_0(x668_outr_Foreach_sm_io_enableOut_0),
    .io_enableOut_1(x668_outr_Foreach_sm_io_enableOut_1),
    .io_childAck_0(x668_outr_Foreach_sm_io_childAck_0),
    .io_childAck_1(x668_outr_Foreach_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@82240.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@82285.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@82293.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1 x668_outr_Foreach_kernelx668_outr_Foreach_concrete1 ( // @[sm_x668_outr_Foreach.scala 120:24:@82327.4]
    .clock(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_clock),
    .reset(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_reset),
    .io_in_x472_A_sram_1_rPort_0_ofs_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0),
    .io_in_x472_A_sram_1_rPort_0_en_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_en_0),
    .io_in_x472_A_sram_1_rPort_0_output_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_output_0),
    .io_in_x471_A_sram_0_rPort_0_ofs_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0),
    .io_in_x471_A_sram_0_rPort_0_en_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_en_0),
    .io_in_x471_A_sram_0_rPort_0_output_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_output_0),
    .io_in_x473_A_sram_2_rPort_0_ofs_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_ofs_0),
    .io_in_x473_A_sram_2_rPort_0_en_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_en_0),
    .io_in_x473_A_sram_2_rPort_0_output_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_output_0),
    .io_in_x539_out_sram_0_wPort_0_ofs_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_ofs_0),
    .io_in_x539_out_sram_0_wPort_0_data_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_data_0),
    .io_in_x539_out_sram_0_wPort_0_en_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_en_0),
    .io_in_instrctrs_6_cycs(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_6_cycs),
    .io_in_instrctrs_6_iters(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_6_iters),
    .io_in_instrctrs_7_cycs(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_7_cycs),
    .io_in_instrctrs_7_iters(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_7_iters),
    .io_in_instrctrs_8_cycs(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_8_cycs),
    .io_in_instrctrs_8_iters(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_8_iters),
    .io_in_instrctrs_9_cycs(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_9_cycs),
    .io_in_instrctrs_9_iters(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_9_iters),
    .io_in_instrctrs_10_cycs(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_10_cycs),
    .io_in_instrctrs_10_iters(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_10_iters),
    .io_in_instrctrs_11_cycs(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_11_cycs),
    .io_in_instrctrs_11_iters(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_11_iters),
    .io_in_instrctrs_12_cycs(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_12_cycs),
    .io_in_instrctrs_12_iters(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_12_iters),
    .io_in_instrctrs_13_cycs(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_13_cycs),
    .io_in_instrctrs_13_iters(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_13_iters),
    .io_in_instrctrs_14_cycs(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_14_cycs),
    .io_in_instrctrs_14_iters(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_14_iters),
    .io_in_instrctrs_15_cycs(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_15_cycs),
    .io_in_instrctrs_15_iters(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_15_iters),
    .io_in_instrctrs_16_cycs(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_16_cycs),
    .io_in_instrctrs_16_iters(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_16_iters),
    .io_in_instrctrs_17_cycs(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_17_cycs),
    .io_in_instrctrs_17_iters(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_17_iters),
    .io_sigsIn_done(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smEnableOuts_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsOut_smDoneIn_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smMaskIn_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0),
    .io_sigsOut_smMaskIn_1(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1),
    .io_rr(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_rr)
  );
  x724_outr_UnitPipe_DenseTransfer_sm x724_outr_UnitPipe_DenseTransfer_sm ( // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@82649.4]
    .clock(x724_outr_UnitPipe_DenseTransfer_sm_clock),
    .reset(x724_outr_UnitPipe_DenseTransfer_sm_reset),
    .io_enable(x724_outr_UnitPipe_DenseTransfer_sm_io_enable),
    .io_done(x724_outr_UnitPipe_DenseTransfer_sm_io_done),
    .io_parentAck(x724_outr_UnitPipe_DenseTransfer_sm_io_parentAck),
    .io_doneIn_0(x724_outr_UnitPipe_DenseTransfer_sm_io_doneIn_0),
    .io_enableOut_0(x724_outr_UnitPipe_DenseTransfer_sm_io_enableOut_0),
    .io_childAck_0(x724_outr_UnitPipe_DenseTransfer_sm_io_childAck_0),
    .io_ctrCopyDone_0(x724_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@82702.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@82710.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1 x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1 ( // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 97:24:@82740.4]
    .clock(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_clock),
    .reset(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_reset),
    .io_in_x670_ready(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_ready),
    .io_in_x670_valid(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_valid),
    .io_in_x670_bits_wdata_0(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_bits_wdata_0),
    .io_in_x670_bits_wstrb(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_bits_wstrb),
    .io_in_x669_ready(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_ready),
    .io_in_x669_valid(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_valid),
    .io_in_x669_bits_addr(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_bits_addr),
    .io_in_x669_bits_size(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_bits_size),
    .io_in_x470_out_host_number(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x470_out_host_number),
    .io_in_x539_out_sram_0_rPort_0_ofs_0(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0),
    .io_in_x539_out_sram_0_rPort_0_en_0(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_en_0),
    .io_in_x539_out_sram_0_rPort_0_backpressure(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure),
    .io_in_x539_out_sram_0_rPort_0_output_0(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_output_0),
    .io_in_x671_ready(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x671_ready),
    .io_in_x671_valid(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x671_valid),
    .io_in_instrctrs_18_cycs(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_18_cycs),
    .io_in_instrctrs_18_iters(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_18_iters),
    .io_in_instrctrs_19_cycs(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_19_cycs),
    .io_in_instrctrs_19_iters(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_19_iters),
    .io_in_instrctrs_20_cycs(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_20_cycs),
    .io_in_instrctrs_20_iters(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_20_iters),
    .io_in_instrctrs_21_cycs(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_21_cycs),
    .io_in_instrctrs_21_iters(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_21_iters),
    .io_in_instrctrs_21_stalls(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_21_stalls),
    .io_in_instrctrs_21_idles(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_21_idles),
    .io_in_instrctrs_22_cycs(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_22_cycs),
    .io_in_instrctrs_22_iters(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_22_iters),
    .io_in_instrctrs_22_stalls(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_22_stalls),
    .io_in_instrctrs_22_idles(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_22_idles),
    .io_in_instrctrs_23_cycs(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_23_cycs),
    .io_in_instrctrs_23_iters(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_23_iters),
    .io_in_instrctrs_23_stalls(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_23_stalls),
    .io_in_instrctrs_23_idles(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_23_idles),
    .io_sigsIn_done(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smEnableOuts_0(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_rr)
  );
  assign _T_190 = io_sigsIn_done == 1'h0; // @[package.scala 100:49:@81647.4]
  assign _T_277 = RetimeWrapper_io_out; // @[package.scala 96:25:@81823.4 package.scala 96:25:@81824.4]
  assign _T_283 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@81831.4 package.scala 96:25:@81832.4]
  assign _T_286 = ~ _T_283; // @[SpatialBlocks.scala 137:99:@81834.4]
  assign _T_359 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@82245.4 package.scala 96:25:@82246.4]
  assign _T_376 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@82290.4 package.scala 96:25:@82291.4]
  assign _T_382 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@82298.4 package.scala 96:25:@82299.4]
  assign _T_385 = ~ _T_382; // @[SpatialBlocks.scala 137:99:@82301.4]
  assign _T_468 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@82707.4 package.scala 96:25:@82708.4]
  assign _T_474 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@82715.4 package.scala 96:25:@82716.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 137:99:@82718.4]
  assign io_in_x670_valid = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_valid; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 59:23:@82894.4]
  assign io_in_x670_bits_wdata_0 = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_bits_wdata_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 59:23:@82893.4]
  assign io_in_x670_bits_wstrb = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_bits_wstrb; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 59:23:@82892.4]
  assign io_in_x669_valid = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_valid; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 60:23:@82898.4]
  assign io_in_x669_bits_addr = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_bits_addr; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 60:23:@82897.4]
  assign io_in_x669_bits_size = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_bits_size; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 60:23:@82896.4]
  assign io_in_x476_ready = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_ready; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 63:23:@82060.4]
  assign io_in_x671_ready = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x671_ready; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 63:23:@82908.4]
  assign io_in_x474_valid = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_valid; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 65:23:@82070.4]
  assign io_in_x474_bits_addr = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_bits_addr; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 65:23:@82069.4]
  assign io_in_x474_bits_size = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_bits_size; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 65:23:@82068.4]
  assign io_in_instrctrs_0_cycs = cycles_RootController_io_count; // @[Ledger.scala 293:21:@81652.4]
  assign io_in_instrctrs_0_iters = iters_RootController_io_count; // @[Ledger.scala 294:22:@81653.4]
  assign io_in_instrctrs_1_cycs = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_1_cycs; // @[Ledger.scala 302:78:@82075.4]
  assign io_in_instrctrs_1_iters = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_1_iters; // @[Ledger.scala 302:78:@82074.4]
  assign io_in_instrctrs_2_cycs = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_2_cycs; // @[Ledger.scala 302:78:@82079.4]
  assign io_in_instrctrs_2_iters = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_2_iters; // @[Ledger.scala 302:78:@82078.4]
  assign io_in_instrctrs_2_stalls = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_2_stalls; // @[Ledger.scala 302:78:@82077.4]
  assign io_in_instrctrs_2_idles = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_2_idles; // @[Ledger.scala 302:78:@82076.4]
  assign io_in_instrctrs_3_cycs = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_3_cycs; // @[Ledger.scala 302:78:@82083.4]
  assign io_in_instrctrs_3_iters = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_3_iters; // @[Ledger.scala 302:78:@82082.4]
  assign io_in_instrctrs_4_cycs = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_4_cycs; // @[Ledger.scala 302:78:@82087.4]
  assign io_in_instrctrs_4_iters = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_4_iters; // @[Ledger.scala 302:78:@82086.4]
  assign io_in_instrctrs_4_stalls = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_4_stalls; // @[Ledger.scala 302:78:@82085.4]
  assign io_in_instrctrs_4_idles = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_4_idles; // @[Ledger.scala 302:78:@82084.4]
  assign io_in_instrctrs_5_cycs = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_5_cycs; // @[Ledger.scala 302:78:@82091.4]
  assign io_in_instrctrs_5_iters = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_5_iters; // @[Ledger.scala 302:78:@82090.4]
  assign io_in_instrctrs_5_stalls = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_5_stalls; // @[Ledger.scala 302:78:@82089.4]
  assign io_in_instrctrs_5_idles = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_5_idles; // @[Ledger.scala 302:78:@82088.4]
  assign io_in_instrctrs_6_cycs = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_6_cycs; // @[Ledger.scala 302:78:@82536.4]
  assign io_in_instrctrs_6_iters = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_6_iters; // @[Ledger.scala 302:78:@82535.4]
  assign io_in_instrctrs_7_cycs = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_7_cycs; // @[Ledger.scala 302:78:@82540.4]
  assign io_in_instrctrs_7_iters = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_7_iters; // @[Ledger.scala 302:78:@82539.4]
  assign io_in_instrctrs_8_cycs = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_8_cycs; // @[Ledger.scala 302:78:@82544.4]
  assign io_in_instrctrs_8_iters = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_8_iters; // @[Ledger.scala 302:78:@82543.4]
  assign io_in_instrctrs_9_cycs = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_9_cycs; // @[Ledger.scala 302:78:@82548.4]
  assign io_in_instrctrs_9_iters = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_9_iters; // @[Ledger.scala 302:78:@82547.4]
  assign io_in_instrctrs_10_cycs = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_10_cycs; // @[Ledger.scala 302:78:@82552.4]
  assign io_in_instrctrs_10_iters = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_10_iters; // @[Ledger.scala 302:78:@82551.4]
  assign io_in_instrctrs_11_cycs = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_11_cycs; // @[Ledger.scala 302:78:@82556.4]
  assign io_in_instrctrs_11_iters = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_11_iters; // @[Ledger.scala 302:78:@82555.4]
  assign io_in_instrctrs_12_cycs = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_12_cycs; // @[Ledger.scala 302:78:@82560.4]
  assign io_in_instrctrs_12_iters = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_12_iters; // @[Ledger.scala 302:78:@82559.4]
  assign io_in_instrctrs_13_cycs = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_13_cycs; // @[Ledger.scala 302:78:@82564.4]
  assign io_in_instrctrs_13_iters = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_13_iters; // @[Ledger.scala 302:78:@82563.4]
  assign io_in_instrctrs_14_cycs = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_14_cycs; // @[Ledger.scala 302:78:@82568.4]
  assign io_in_instrctrs_14_iters = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_14_iters; // @[Ledger.scala 302:78:@82567.4]
  assign io_in_instrctrs_15_cycs = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_15_cycs; // @[Ledger.scala 302:78:@82572.4]
  assign io_in_instrctrs_15_iters = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_15_iters; // @[Ledger.scala 302:78:@82571.4]
  assign io_in_instrctrs_16_cycs = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_16_cycs; // @[Ledger.scala 302:78:@82576.4]
  assign io_in_instrctrs_16_iters = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_16_iters; // @[Ledger.scala 302:78:@82575.4]
  assign io_in_instrctrs_17_cycs = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_17_cycs; // @[Ledger.scala 302:78:@82580.4]
  assign io_in_instrctrs_17_iters = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_instrctrs_17_iters; // @[Ledger.scala 302:78:@82579.4]
  assign io_in_instrctrs_18_cycs = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_18_cycs; // @[Ledger.scala 302:78:@82912.4]
  assign io_in_instrctrs_18_iters = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_18_iters; // @[Ledger.scala 302:78:@82911.4]
  assign io_in_instrctrs_19_cycs = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_19_cycs; // @[Ledger.scala 302:78:@82916.4]
  assign io_in_instrctrs_19_iters = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_19_iters; // @[Ledger.scala 302:78:@82915.4]
  assign io_in_instrctrs_20_cycs = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_20_cycs; // @[Ledger.scala 302:78:@82920.4]
  assign io_in_instrctrs_20_iters = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_20_iters; // @[Ledger.scala 302:78:@82919.4]
  assign io_in_instrctrs_21_cycs = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_21_cycs; // @[Ledger.scala 302:78:@82924.4]
  assign io_in_instrctrs_21_iters = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_21_iters; // @[Ledger.scala 302:78:@82923.4]
  assign io_in_instrctrs_21_stalls = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_21_stalls; // @[Ledger.scala 302:78:@82922.4]
  assign io_in_instrctrs_21_idles = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_21_idles; // @[Ledger.scala 302:78:@82921.4]
  assign io_in_instrctrs_22_cycs = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_22_cycs; // @[Ledger.scala 302:78:@82928.4]
  assign io_in_instrctrs_22_iters = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_22_iters; // @[Ledger.scala 302:78:@82927.4]
  assign io_in_instrctrs_22_stalls = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_22_stalls; // @[Ledger.scala 302:78:@82926.4]
  assign io_in_instrctrs_22_idles = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_22_idles; // @[Ledger.scala 302:78:@82925.4]
  assign io_in_instrctrs_23_cycs = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_23_cycs; // @[Ledger.scala 302:78:@82932.4]
  assign io_in_instrctrs_23_iters = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_23_iters; // @[Ledger.scala 302:78:@82931.4]
  assign io_in_instrctrs_23_stalls = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_23_stalls; // @[Ledger.scala 302:78:@82930.4]
  assign io_in_instrctrs_23_idles = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_instrctrs_23_idles; // @[Ledger.scala 302:78:@82929.4]
  assign io_sigsOut_smDoneIn_0 = x538_outr_UnitPipe_DenseTransfer_sm_io_done; // @[SpatialBlocks.scala 155:56:@81841.4]
  assign io_sigsOut_smDoneIn_1 = x668_outr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@82308.4]
  assign io_sigsOut_smDoneIn_2 = x724_outr_UnitPipe_DenseTransfer_sm_io_done; // @[SpatialBlocks.scala 155:56:@82725.4]
  assign cycles_RootController_clock = clock; // @[:@81641.4]
  assign cycles_RootController_reset = reset; // @[:@81642.4]
  assign cycles_RootController_io_enable = io_sigsIn_baseEn; // @[sm_RootController.scala 88:39:@81646.4]
  assign iters_RootController_clock = clock; // @[:@81644.4]
  assign iters_RootController_reset = reset; // @[:@81645.4]
  assign iters_RootController_io_enable = io_sigsIn_done & _T_193; // @[sm_RootController.scala 89:38:@81651.4]
  assign x471_A_sram_0_clock = clock; // @[:@81657.4]
  assign x471_A_sram_0_reset = reset; // @[:@81658.4]
  assign x471_A_sram_0_io_rPort_0_ofs_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@82519.4]
  assign x471_A_sram_0_io_rPort_0_en_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@82518.4]
  assign x471_A_sram_0_io_rPort_0_backpressure = 1'h1; // @[MemInterfaceType.scala 66:44:@82517.4]
  assign x471_A_sram_0_io_wPort_0_ofs_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@82056.4]
  assign x471_A_sram_0_io_wPort_0_data_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@82055.4]
  assign x471_A_sram_0_io_wPort_0_en_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@82051.4]
  assign x472_A_sram_1_clock = clock; // @[:@81674.4]
  assign x472_A_sram_1_reset = reset; // @[:@81675.4]
  assign x472_A_sram_1_io_rPort_0_ofs_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@82514.4]
  assign x472_A_sram_1_io_rPort_0_en_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@82513.4]
  assign x472_A_sram_1_io_rPort_0_backpressure = 1'h1; // @[MemInterfaceType.scala 66:44:@82512.4]
  assign x472_A_sram_1_io_wPort_0_ofs_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@82049.4]
  assign x472_A_sram_1_io_wPort_0_data_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@82048.4]
  assign x472_A_sram_1_io_wPort_0_en_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@82044.4]
  assign x473_A_sram_2_clock = clock; // @[:@81691.4]
  assign x473_A_sram_2_reset = reset; // @[:@81692.4]
  assign x473_A_sram_2_io_rPort_0_ofs_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@82524.4]
  assign x473_A_sram_2_io_rPort_0_en_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@82523.4]
  assign x473_A_sram_2_io_rPort_0_backpressure = 1'h1; // @[MemInterfaceType.scala 66:44:@82522.4]
  assign x473_A_sram_2_io_wPort_0_ofs_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@82066.4]
  assign x473_A_sram_2_io_wPort_0_data_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@82065.4]
  assign x473_A_sram_2_io_wPort_0_en_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@82061.4]
  assign x538_outr_UnitPipe_DenseTransfer_sm_clock = clock; // @[:@81756.4]
  assign x538_outr_UnitPipe_DenseTransfer_sm_reset = reset; // @[:@81757.4]
  assign x538_outr_UnitPipe_DenseTransfer_sm_io_enable = _T_277 & _T_286; // @[SpatialBlocks.scala 139:18:@81838.4]
  assign x538_outr_UnitPipe_DenseTransfer_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@81840.4]
  assign x538_outr_UnitPipe_DenseTransfer_sm_io_doneIn_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@81808.4]
  assign x538_outr_UnitPipe_DenseTransfer_sm_io_doneIn_1 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:72:@81809.4]
  assign x538_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:95:@81855.4]
  assign x538_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_1 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:95:@81856.4]
  assign RetimeWrapper_clock = clock; // @[:@81819.4]
  assign RetimeWrapper_reset = reset; // @[:@81820.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@81822.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@81821.4]
  assign RetimeWrapper_1_clock = clock; // @[:@81827.4]
  assign RetimeWrapper_1_reset = reset; // @[:@81828.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@81830.4]
  assign RetimeWrapper_1_io_in = x538_outr_UnitPipe_DenseTransfer_sm_io_done; // @[package.scala 94:16:@81829.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_clock = clock; // @[:@81858.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_reset = reset; // @[:@81859.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x468_A_dram_number = io_in_x468_A_dram_number; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 60:30:@82043.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_valid = io_in_x476_valid; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 63:23:@82059.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_bits_rdata_0 = io_in_x476_bits_rdata_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 63:23:@82058.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_ready = io_in_x474_ready; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 65:23:@82071.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_done = x538_outr_UnitPipe_DenseTransfer_sm_io_done; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 120:22:@82119.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_baseEn = _T_277 & _T_286; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 120:22:@82111.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_0 = x538_outr_UnitPipe_DenseTransfer_sm_io_enableOut_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 120:22:@82107.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_1 = x538_outr_UnitPipe_DenseTransfer_sm_io_enableOut_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 120:22:@82108.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_0 = x538_outr_UnitPipe_DenseTransfer_sm_io_childAck_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 120:22:@82103.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_1 = x538_outr_UnitPipe_DenseTransfer_sm_io_childAck_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 120:22:@82104.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_rr = io_rr; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 119:18:@82092.4]
  assign x539_out_sram_0_clock = clock; // @[:@82132.4]
  assign x539_out_sram_0_reset = reset; // @[:@82133.4]
  assign x539_out_sram_0_io_rPort_0_ofs_0 = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@82904.4]
  assign x539_out_sram_0_io_rPort_0_en_0 = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@82903.4]
  assign x539_out_sram_0_io_rPort_0_backpressure = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@82902.4]
  assign x539_out_sram_0_io_wPort_0_ofs_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@82531.4]
  assign x539_out_sram_0_io_wPort_0_data_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@82530.4]
  assign x539_out_sram_0_io_wPort_0_en_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@82526.4]
  assign x541_ctrchain_clock = clock; // @[:@82149.4]
  assign x541_ctrchain_reset = reset; // @[:@82150.4]
  assign x541_ctrchain_io_input_reset = x668_outr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@82326.4]
  assign x541_ctrchain_io_input_enable = x668_outr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 158:42:@82325.4]
  assign x668_outr_Foreach_sm_clock = clock; // @[:@82207.4]
  assign x668_outr_Foreach_sm_reset = reset; // @[:@82208.4]
  assign x668_outr_Foreach_sm_io_enable = _T_376 & _T_385; // @[SpatialBlocks.scala 139:18:@82305.4]
  assign x668_outr_Foreach_sm_io_ctrDone = io_rr ? _T_359 : 1'h0; // @[sm_RootController.scala 108:39:@82248.4]
  assign x668_outr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 141:21:@82307.4]
  assign x668_outr_Foreach_sm_io_doneIn_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@82275.4]
  assign x668_outr_Foreach_sm_io_doneIn_1 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:72:@82276.4]
  assign x668_outr_Foreach_sm_io_maskIn_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0; // @[SpatialBlocks.scala 131:72:@82277.4]
  assign x668_outr_Foreach_sm_io_maskIn_1 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1; // @[SpatialBlocks.scala 131:72:@82278.4]
  assign RetimeWrapper_2_clock = clock; // @[:@82241.4]
  assign RetimeWrapper_2_reset = reset; // @[:@82242.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@82244.4]
  assign RetimeWrapper_2_io_in = x541_ctrchain_io_output_done; // @[package.scala 94:16:@82243.4]
  assign RetimeWrapper_3_clock = clock; // @[:@82286.4]
  assign RetimeWrapper_3_reset = reset; // @[:@82287.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@82289.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@82288.4]
  assign RetimeWrapper_4_clock = clock; // @[:@82294.4]
  assign RetimeWrapper_4_reset = reset; // @[:@82295.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@82297.4]
  assign RetimeWrapper_4_io_in = x668_outr_Foreach_sm_io_done; // @[package.scala 94:16:@82296.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_clock = clock; // @[:@82328.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_reset = reset; // @[:@82329.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_output_0 = x472_A_sram_1_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@82511.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_output_0 = x471_A_sram_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@82516.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_output_0 = x473_A_sram_2_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@82521.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_done = x668_outr_Foreach_sm_io_done; // @[sm_x668_outr_Foreach.scala 126:22:@82603.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_baseEn = _T_376 & _T_385; // @[sm_x668_outr_Foreach.scala 126:22:@82595.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0 = x668_outr_Foreach_sm_io_enableOut_0; // @[sm_x668_outr_Foreach.scala 126:22:@82591.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1 = x668_outr_Foreach_sm_io_enableOut_1; // @[sm_x668_outr_Foreach.scala 126:22:@82592.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0 = x668_outr_Foreach_sm_io_childAck_0; // @[sm_x668_outr_Foreach.scala 126:22:@82587.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1 = x668_outr_Foreach_sm_io_childAck_1; // @[sm_x668_outr_Foreach.scala 126:22:@82588.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{23{x541_ctrchain_io_output_counts_0[8]}},x541_ctrchain_io_output_counts_0}; // @[sm_x668_outr_Foreach.scala 126:22:@82586.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x541_ctrchain_io_output_oobs_0; // @[sm_x668_outr_Foreach.scala 126:22:@82585.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_rr = io_rr; // @[sm_x668_outr_Foreach.scala 125:18:@82581.4]
  assign x724_outr_UnitPipe_DenseTransfer_sm_clock = clock; // @[:@82650.4]
  assign x724_outr_UnitPipe_DenseTransfer_sm_reset = reset; // @[:@82651.4]
  assign x724_outr_UnitPipe_DenseTransfer_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 139:18:@82722.4]
  assign x724_outr_UnitPipe_DenseTransfer_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 141:21:@82724.4]
  assign x724_outr_UnitPipe_DenseTransfer_sm_io_doneIn_0 = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@82694.4]
  assign x724_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_0 = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:95:@82739.4]
  assign RetimeWrapper_5_clock = clock; // @[:@82703.4]
  assign RetimeWrapper_5_reset = reset; // @[:@82704.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@82706.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@82705.4]
  assign RetimeWrapper_6_clock = clock; // @[:@82711.4]
  assign RetimeWrapper_6_reset = reset; // @[:@82712.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@82714.4]
  assign RetimeWrapper_6_io_in = x724_outr_UnitPipe_DenseTransfer_sm_io_done; // @[package.scala 94:16:@82713.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_clock = clock; // @[:@82741.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_reset = reset; // @[:@82742.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_ready = io_in_x670_ready; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 59:23:@82895.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_ready = io_in_x669_ready; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 60:23:@82899.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x470_out_host_number = io_in_x470_out_host_number; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 61:32:@82900.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_output_0 = x539_out_sram_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@82901.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x671_valid = io_in_x671_valid; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 63:23:@82907.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_done = x724_outr_UnitPipe_DenseTransfer_sm_io_done; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 103:22:@82952.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_baseEn = _T_468 & _T_477; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 103:22:@82944.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_0 = x724_outr_UnitPipe_DenseTransfer_sm_io_enableOut_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 103:22:@82941.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_0 = x724_outr_UnitPipe_DenseTransfer_sm_io_childAck_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 103:22:@82939.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_rr = io_rr; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 102:18:@82933.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_193 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_193 <= 1'h0;
    end else begin
      _T_193 <= _T_190;
    end
  end
endmodule
module AccelUnit( // @[:@82961.2]
  input          clock, // @[:@82962.4]
  input          reset, // @[:@82963.4]
  input          io_enable, // @[:@82964.4]
  output         io_done, // @[:@82964.4]
  input          io_reset, // @[:@82964.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@82964.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@82964.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@82964.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@82964.4]
  output         io_memStreams_loads_0_data_ready, // @[:@82964.4]
  input          io_memStreams_loads_0_data_valid, // @[:@82964.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@82964.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@82964.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@82964.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@82964.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@82964.4]
  input          io_memStreams_stores_0_data_ready, // @[:@82964.4]
  output         io_memStreams_stores_0_data_valid, // @[:@82964.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@82964.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@82964.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@82964.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@82964.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@82964.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@82964.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_16, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_17, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_18, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_19, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_20, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_21, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_22, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_23, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_24, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_25, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_26, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_27, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_28, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_29, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_30, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_31, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_32, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_33, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_34, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_35, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_36, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_37, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_38, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_39, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_40, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_41, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_42, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_43, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_44, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_45, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_46, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_47, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_48, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_49, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_50, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_51, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_52, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_53, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_54, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_55, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_56, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_57, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_58, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_59, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_60, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_61, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_62, // @[:@82964.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_63, // @[:@82964.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@82964.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_0, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_1, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_2, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_3, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_4, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_5, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_6, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_7, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_8, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_9, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_10, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_11, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_12, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_13, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_14, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_15, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_16, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_17, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_18, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_19, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_20, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_21, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_22, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_23, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_24, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_25, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_26, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_27, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_28, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_29, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_30, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_31, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_32, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_33, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_34, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_35, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_36, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_37, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_38, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_39, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_40, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_41, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_42, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_43, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_44, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_45, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_46, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_47, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_48, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_49, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_50, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_51, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_52, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_53, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_54, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_55, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_56, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_57, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_58, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_59, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_60, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_61, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_62, // @[:@82964.4]
  input  [7:0]   io_memStreams_gathers_0_data_bits_63, // @[:@82964.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@82964.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_16, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_17, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_18, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_19, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_20, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_21, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_22, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_23, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_24, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_25, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_26, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_27, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_28, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_29, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_30, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_31, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_32, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_33, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_34, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_35, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_36, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_37, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_38, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_39, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_40, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_41, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_42, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_43, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_44, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_45, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_46, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_47, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_48, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_49, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_50, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_51, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_52, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_53, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_54, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_55, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_56, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_57, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_58, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_59, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_60, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_61, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_62, // @[:@82964.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_63, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_16, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_17, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_18, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_19, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_20, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_21, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_22, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_23, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_24, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_25, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_26, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_27, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_28, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_29, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_30, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_31, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_32, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_33, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_34, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_35, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_36, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_37, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_38, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_39, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_40, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_41, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_42, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_43, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_44, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_45, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_46, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_47, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_48, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_49, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_50, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_51, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_52, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_53, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_54, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_55, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_56, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_57, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_58, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_59, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_60, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_61, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_62, // @[:@82964.4]
  output [7:0]   io_memStreams_scatters_0_cmd_bits_wdata_63, // @[:@82964.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@82964.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@82964.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@82964.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@82964.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@82964.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@82964.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@82964.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@82964.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@82964.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@82964.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@82964.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@82964.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@82964.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@82964.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@82964.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@82964.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@82964.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@82964.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@82964.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@82964.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@82964.4]
  output         io_heap_0_req_valid, // @[:@82964.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@82964.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@82964.4]
  input          io_heap_0_resp_valid, // @[:@82964.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@82964.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@82964.4]
  input  [63:0]  io_argIns_0, // @[:@82964.4]
  input  [63:0]  io_argIns_1, // @[:@82964.4]
  input          io_argOuts_0_port_ready, // @[:@82964.4]
  output         io_argOuts_0_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_0_echo, // @[:@82964.4]
  input          io_argOuts_1_port_ready, // @[:@82964.4]
  output         io_argOuts_1_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_1_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_1_echo, // @[:@82964.4]
  input          io_argOuts_2_port_ready, // @[:@82964.4]
  output         io_argOuts_2_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_2_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_2_echo, // @[:@82964.4]
  input          io_argOuts_3_port_ready, // @[:@82964.4]
  output         io_argOuts_3_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_3_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_3_echo, // @[:@82964.4]
  input          io_argOuts_4_port_ready, // @[:@82964.4]
  output         io_argOuts_4_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_4_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_4_echo, // @[:@82964.4]
  input          io_argOuts_5_port_ready, // @[:@82964.4]
  output         io_argOuts_5_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_5_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_5_echo, // @[:@82964.4]
  input          io_argOuts_6_port_ready, // @[:@82964.4]
  output         io_argOuts_6_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_6_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_6_echo, // @[:@82964.4]
  input          io_argOuts_7_port_ready, // @[:@82964.4]
  output         io_argOuts_7_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_7_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_7_echo, // @[:@82964.4]
  input          io_argOuts_8_port_ready, // @[:@82964.4]
  output         io_argOuts_8_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_8_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_8_echo, // @[:@82964.4]
  input          io_argOuts_9_port_ready, // @[:@82964.4]
  output         io_argOuts_9_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_9_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_9_echo, // @[:@82964.4]
  input          io_argOuts_10_port_ready, // @[:@82964.4]
  output         io_argOuts_10_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_10_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_10_echo, // @[:@82964.4]
  input          io_argOuts_11_port_ready, // @[:@82964.4]
  output         io_argOuts_11_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_11_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_11_echo, // @[:@82964.4]
  input          io_argOuts_12_port_ready, // @[:@82964.4]
  output         io_argOuts_12_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_12_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_12_echo, // @[:@82964.4]
  input          io_argOuts_13_port_ready, // @[:@82964.4]
  output         io_argOuts_13_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_13_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_13_echo, // @[:@82964.4]
  input          io_argOuts_14_port_ready, // @[:@82964.4]
  output         io_argOuts_14_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_14_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_14_echo, // @[:@82964.4]
  input          io_argOuts_15_port_ready, // @[:@82964.4]
  output         io_argOuts_15_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_15_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_15_echo, // @[:@82964.4]
  input          io_argOuts_16_port_ready, // @[:@82964.4]
  output         io_argOuts_16_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_16_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_16_echo, // @[:@82964.4]
  input          io_argOuts_17_port_ready, // @[:@82964.4]
  output         io_argOuts_17_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_17_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_17_echo, // @[:@82964.4]
  input          io_argOuts_18_port_ready, // @[:@82964.4]
  output         io_argOuts_18_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_18_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_18_echo, // @[:@82964.4]
  input          io_argOuts_19_port_ready, // @[:@82964.4]
  output         io_argOuts_19_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_19_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_19_echo, // @[:@82964.4]
  input          io_argOuts_20_port_ready, // @[:@82964.4]
  output         io_argOuts_20_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_20_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_20_echo, // @[:@82964.4]
  input          io_argOuts_21_port_ready, // @[:@82964.4]
  output         io_argOuts_21_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_21_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_21_echo, // @[:@82964.4]
  input          io_argOuts_22_port_ready, // @[:@82964.4]
  output         io_argOuts_22_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_22_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_22_echo, // @[:@82964.4]
  input          io_argOuts_23_port_ready, // @[:@82964.4]
  output         io_argOuts_23_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_23_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_23_echo, // @[:@82964.4]
  input          io_argOuts_24_port_ready, // @[:@82964.4]
  output         io_argOuts_24_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_24_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_24_echo, // @[:@82964.4]
  input          io_argOuts_25_port_ready, // @[:@82964.4]
  output         io_argOuts_25_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_25_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_25_echo, // @[:@82964.4]
  input          io_argOuts_26_port_ready, // @[:@82964.4]
  output         io_argOuts_26_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_26_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_26_echo, // @[:@82964.4]
  input          io_argOuts_27_port_ready, // @[:@82964.4]
  output         io_argOuts_27_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_27_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_27_echo, // @[:@82964.4]
  input          io_argOuts_28_port_ready, // @[:@82964.4]
  output         io_argOuts_28_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_28_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_28_echo, // @[:@82964.4]
  input          io_argOuts_29_port_ready, // @[:@82964.4]
  output         io_argOuts_29_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_29_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_29_echo, // @[:@82964.4]
  input          io_argOuts_30_port_ready, // @[:@82964.4]
  output         io_argOuts_30_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_30_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_30_echo, // @[:@82964.4]
  input          io_argOuts_31_port_ready, // @[:@82964.4]
  output         io_argOuts_31_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_31_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_31_echo, // @[:@82964.4]
  input          io_argOuts_32_port_ready, // @[:@82964.4]
  output         io_argOuts_32_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_32_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_32_echo, // @[:@82964.4]
  input          io_argOuts_33_port_ready, // @[:@82964.4]
  output         io_argOuts_33_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_33_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_33_echo, // @[:@82964.4]
  input          io_argOuts_34_port_ready, // @[:@82964.4]
  output         io_argOuts_34_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_34_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_34_echo, // @[:@82964.4]
  input          io_argOuts_35_port_ready, // @[:@82964.4]
  output         io_argOuts_35_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_35_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_35_echo, // @[:@82964.4]
  input          io_argOuts_36_port_ready, // @[:@82964.4]
  output         io_argOuts_36_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_36_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_36_echo, // @[:@82964.4]
  input          io_argOuts_37_port_ready, // @[:@82964.4]
  output         io_argOuts_37_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_37_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_37_echo, // @[:@82964.4]
  input          io_argOuts_38_port_ready, // @[:@82964.4]
  output         io_argOuts_38_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_38_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_38_echo, // @[:@82964.4]
  input          io_argOuts_39_port_ready, // @[:@82964.4]
  output         io_argOuts_39_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_39_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_39_echo, // @[:@82964.4]
  input          io_argOuts_40_port_ready, // @[:@82964.4]
  output         io_argOuts_40_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_40_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_40_echo, // @[:@82964.4]
  input          io_argOuts_41_port_ready, // @[:@82964.4]
  output         io_argOuts_41_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_41_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_41_echo, // @[:@82964.4]
  input          io_argOuts_42_port_ready, // @[:@82964.4]
  output         io_argOuts_42_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_42_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_42_echo, // @[:@82964.4]
  input          io_argOuts_43_port_ready, // @[:@82964.4]
  output         io_argOuts_43_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_43_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_43_echo, // @[:@82964.4]
  input          io_argOuts_44_port_ready, // @[:@82964.4]
  output         io_argOuts_44_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_44_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_44_echo, // @[:@82964.4]
  input          io_argOuts_45_port_ready, // @[:@82964.4]
  output         io_argOuts_45_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_45_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_45_echo, // @[:@82964.4]
  input          io_argOuts_46_port_ready, // @[:@82964.4]
  output         io_argOuts_46_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_46_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_46_echo, // @[:@82964.4]
  input          io_argOuts_47_port_ready, // @[:@82964.4]
  output         io_argOuts_47_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_47_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_47_echo, // @[:@82964.4]
  input          io_argOuts_48_port_ready, // @[:@82964.4]
  output         io_argOuts_48_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_48_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_48_echo, // @[:@82964.4]
  input          io_argOuts_49_port_ready, // @[:@82964.4]
  output         io_argOuts_49_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_49_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_49_echo, // @[:@82964.4]
  input          io_argOuts_50_port_ready, // @[:@82964.4]
  output         io_argOuts_50_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_50_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_50_echo, // @[:@82964.4]
  input          io_argOuts_51_port_ready, // @[:@82964.4]
  output         io_argOuts_51_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_51_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_51_echo, // @[:@82964.4]
  input          io_argOuts_52_port_ready, // @[:@82964.4]
  output         io_argOuts_52_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_52_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_52_echo, // @[:@82964.4]
  input          io_argOuts_53_port_ready, // @[:@82964.4]
  output         io_argOuts_53_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_53_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_53_echo, // @[:@82964.4]
  input          io_argOuts_54_port_ready, // @[:@82964.4]
  output         io_argOuts_54_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_54_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_54_echo, // @[:@82964.4]
  input          io_argOuts_55_port_ready, // @[:@82964.4]
  output         io_argOuts_55_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_55_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_55_echo, // @[:@82964.4]
  input          io_argOuts_56_port_ready, // @[:@82964.4]
  output         io_argOuts_56_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_56_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_56_echo, // @[:@82964.4]
  input          io_argOuts_57_port_ready, // @[:@82964.4]
  output         io_argOuts_57_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_57_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_57_echo, // @[:@82964.4]
  input          io_argOuts_58_port_ready, // @[:@82964.4]
  output         io_argOuts_58_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_58_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_58_echo, // @[:@82964.4]
  input          io_argOuts_59_port_ready, // @[:@82964.4]
  output         io_argOuts_59_port_valid, // @[:@82964.4]
  output [63:0]  io_argOuts_59_port_bits, // @[:@82964.4]
  input  [63:0]  io_argOuts_59_echo // @[:@82964.4]
);
  wire  SingleCounter_clock; // @[Main.scala 42:32:@83525.4]
  wire  SingleCounter_reset; // @[Main.scala 42:32:@83525.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 42:32:@83525.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 42:32:@83525.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@83543.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@83543.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@83543.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@83543.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@83543.4]
  wire  SRFF_clock; // @[Main.scala 47:28:@83672.4]
  wire  SRFF_reset; // @[Main.scala 47:28:@83672.4]
  wire  SRFF_io_input_set; // @[Main.scala 47:28:@83672.4]
  wire  SRFF_io_input_reset; // @[Main.scala 47:28:@83672.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 47:28:@83672.4]
  wire  SRFF_io_output; // @[Main.scala 47:28:@83672.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@83721.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@83721.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@83721.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@83721.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@83721.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@83721.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@83721.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@83721.4]
  wire  RootController_sm_io_doneIn_1; // @[sm_RootController.scala 36:18:@83721.4]
  wire  RootController_sm_io_doneIn_2; // @[sm_RootController.scala 36:18:@83721.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@83721.4]
  wire  RootController_sm_io_enableOut_1; // @[sm_RootController.scala 36:18:@83721.4]
  wire  RootController_sm_io_enableOut_2; // @[sm_RootController.scala 36:18:@83721.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@83721.4]
  wire  RootController_sm_io_childAck_1; // @[sm_RootController.scala 36:18:@83721.4]
  wire  RootController_sm_io_childAck_2; // @[sm_RootController.scala 36:18:@83721.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@83763.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@83763.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@83763.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@83763.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@83763.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x468_A_dram_number; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_in_x670_ready; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_in_x670_valid; // @[sm_RootController.scala 125:24:@83837.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x670_bits_wdata_0; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_in_x670_bits_wstrb; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_in_x669_ready; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_in_x669_valid; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x669_bits_addr; // @[sm_RootController.scala 125:24:@83837.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x669_bits_size; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_in_x476_ready; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_in_x476_valid; // @[sm_RootController.scala 125:24:@83837.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x476_bits_rdata_0; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x470_out_host_number; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_in_x671_ready; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_in_x671_valid; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_in_x474_ready; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_in_x474_valid; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x474_bits_addr; // @[sm_RootController.scala 125:24:@83837.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x474_bits_size; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_0_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_0_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_1_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_1_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_2_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_2_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_2_stalls; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_2_idles; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_3_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_3_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_4_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_4_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_4_stalls; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_4_idles; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_5_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_5_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_5_stalls; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_5_idles; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_6_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_6_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_7_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_7_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_8_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_8_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_9_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_9_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_10_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_10_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_11_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_11_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_12_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_12_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_13_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_13_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_14_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_14_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_15_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_15_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_16_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_16_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_17_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_17_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_18_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_18_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_19_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_19_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_20_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_20_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_21_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_21_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_21_stalls; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_21_idles; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_22_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_22_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_22_stalls; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_22_idles; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_23_cycs; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_23_iters; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_23_stalls; // @[sm_RootController.scala 125:24:@83837.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_instrctrs_23_idles; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_done; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_baseEn; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_2; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_2; // @[sm_RootController.scala 125:24:@83837.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 125:24:@83837.4]
  wire  _T_1263; // @[package.scala 96:25:@83548.4 package.scala 96:25:@83549.4]
  wire  _T_1376; // @[Main.scala 49:50:@83759.4]
  wire  _T_1377; // @[Main.scala 49:59:@83760.4]
  wire  _T_1391; // @[package.scala 100:49:@83781.4]
  reg  _T_1394; // @[package.scala 48:56:@83782.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 42:32:@83525.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@83543.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 47:28:@83672.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@83721.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_doneIn_1(RootController_sm_io_doneIn_1),
    .io_doneIn_2(RootController_sm_io_doneIn_2),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_enableOut_1(RootController_sm_io_enableOut_1),
    .io_enableOut_2(RootController_sm_io_enableOut_2),
    .io_childAck_0(RootController_sm_io_childAck_0),
    .io_childAck_1(RootController_sm_io_childAck_1),
    .io_childAck_2(RootController_sm_io_childAck_2)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@83763.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 125:24:@83837.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x468_A_dram_number(RootController_kernelRootController_concrete1_io_in_x468_A_dram_number),
    .io_in_x670_ready(RootController_kernelRootController_concrete1_io_in_x670_ready),
    .io_in_x670_valid(RootController_kernelRootController_concrete1_io_in_x670_valid),
    .io_in_x670_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x670_bits_wdata_0),
    .io_in_x670_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x670_bits_wstrb),
    .io_in_x669_ready(RootController_kernelRootController_concrete1_io_in_x669_ready),
    .io_in_x669_valid(RootController_kernelRootController_concrete1_io_in_x669_valid),
    .io_in_x669_bits_addr(RootController_kernelRootController_concrete1_io_in_x669_bits_addr),
    .io_in_x669_bits_size(RootController_kernelRootController_concrete1_io_in_x669_bits_size),
    .io_in_x476_ready(RootController_kernelRootController_concrete1_io_in_x476_ready),
    .io_in_x476_valid(RootController_kernelRootController_concrete1_io_in_x476_valid),
    .io_in_x476_bits_rdata_0(RootController_kernelRootController_concrete1_io_in_x476_bits_rdata_0),
    .io_in_x470_out_host_number(RootController_kernelRootController_concrete1_io_in_x470_out_host_number),
    .io_in_x671_ready(RootController_kernelRootController_concrete1_io_in_x671_ready),
    .io_in_x671_valid(RootController_kernelRootController_concrete1_io_in_x671_valid),
    .io_in_x474_ready(RootController_kernelRootController_concrete1_io_in_x474_ready),
    .io_in_x474_valid(RootController_kernelRootController_concrete1_io_in_x474_valid),
    .io_in_x474_bits_addr(RootController_kernelRootController_concrete1_io_in_x474_bits_addr),
    .io_in_x474_bits_size(RootController_kernelRootController_concrete1_io_in_x474_bits_size),
    .io_in_instrctrs_0_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_0_cycs),
    .io_in_instrctrs_0_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_0_iters),
    .io_in_instrctrs_1_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_1_cycs),
    .io_in_instrctrs_1_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_1_iters),
    .io_in_instrctrs_2_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_2_cycs),
    .io_in_instrctrs_2_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_2_iters),
    .io_in_instrctrs_2_stalls(RootController_kernelRootController_concrete1_io_in_instrctrs_2_stalls),
    .io_in_instrctrs_2_idles(RootController_kernelRootController_concrete1_io_in_instrctrs_2_idles),
    .io_in_instrctrs_3_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_3_cycs),
    .io_in_instrctrs_3_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_3_iters),
    .io_in_instrctrs_4_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_4_cycs),
    .io_in_instrctrs_4_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_4_iters),
    .io_in_instrctrs_4_stalls(RootController_kernelRootController_concrete1_io_in_instrctrs_4_stalls),
    .io_in_instrctrs_4_idles(RootController_kernelRootController_concrete1_io_in_instrctrs_4_idles),
    .io_in_instrctrs_5_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_5_cycs),
    .io_in_instrctrs_5_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_5_iters),
    .io_in_instrctrs_5_stalls(RootController_kernelRootController_concrete1_io_in_instrctrs_5_stalls),
    .io_in_instrctrs_5_idles(RootController_kernelRootController_concrete1_io_in_instrctrs_5_idles),
    .io_in_instrctrs_6_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_6_cycs),
    .io_in_instrctrs_6_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_6_iters),
    .io_in_instrctrs_7_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_7_cycs),
    .io_in_instrctrs_7_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_7_iters),
    .io_in_instrctrs_8_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_8_cycs),
    .io_in_instrctrs_8_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_8_iters),
    .io_in_instrctrs_9_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_9_cycs),
    .io_in_instrctrs_9_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_9_iters),
    .io_in_instrctrs_10_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_10_cycs),
    .io_in_instrctrs_10_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_10_iters),
    .io_in_instrctrs_11_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_11_cycs),
    .io_in_instrctrs_11_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_11_iters),
    .io_in_instrctrs_12_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_12_cycs),
    .io_in_instrctrs_12_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_12_iters),
    .io_in_instrctrs_13_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_13_cycs),
    .io_in_instrctrs_13_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_13_iters),
    .io_in_instrctrs_14_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_14_cycs),
    .io_in_instrctrs_14_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_14_iters),
    .io_in_instrctrs_15_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_15_cycs),
    .io_in_instrctrs_15_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_15_iters),
    .io_in_instrctrs_16_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_16_cycs),
    .io_in_instrctrs_16_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_16_iters),
    .io_in_instrctrs_17_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_17_cycs),
    .io_in_instrctrs_17_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_17_iters),
    .io_in_instrctrs_18_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_18_cycs),
    .io_in_instrctrs_18_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_18_iters),
    .io_in_instrctrs_19_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_19_cycs),
    .io_in_instrctrs_19_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_19_iters),
    .io_in_instrctrs_20_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_20_cycs),
    .io_in_instrctrs_20_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_20_iters),
    .io_in_instrctrs_21_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_21_cycs),
    .io_in_instrctrs_21_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_21_iters),
    .io_in_instrctrs_21_stalls(RootController_kernelRootController_concrete1_io_in_instrctrs_21_stalls),
    .io_in_instrctrs_21_idles(RootController_kernelRootController_concrete1_io_in_instrctrs_21_idles),
    .io_in_instrctrs_22_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_22_cycs),
    .io_in_instrctrs_22_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_22_iters),
    .io_in_instrctrs_22_stalls(RootController_kernelRootController_concrete1_io_in_instrctrs_22_stalls),
    .io_in_instrctrs_22_idles(RootController_kernelRootController_concrete1_io_in_instrctrs_22_idles),
    .io_in_instrctrs_23_cycs(RootController_kernelRootController_concrete1_io_in_instrctrs_23_cycs),
    .io_in_instrctrs_23_iters(RootController_kernelRootController_concrete1_io_in_instrctrs_23_iters),
    .io_in_instrctrs_23_stalls(RootController_kernelRootController_concrete1_io_in_instrctrs_23_stalls),
    .io_in_instrctrs_23_idles(RootController_kernelRootController_concrete1_io_in_instrctrs_23_idles),
    .io_sigsIn_done(RootController_kernelRootController_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(RootController_kernelRootController_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_2),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_1263 = RetimeWrapper_io_out; // @[package.scala 96:25:@83548.4 package.scala 96:25:@83549.4]
  assign _T_1376 = io_enable & _T_1263; // @[Main.scala 49:50:@83759.4]
  assign _T_1377 = ~ SRFF_io_output; // @[Main.scala 49:59:@83760.4]
  assign _T_1391 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@83781.4]
  assign io_done = SRFF_io_output; // @[Main.scala 56:23:@83780.4]
  assign io_memStreams_loads_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x474_valid; // @[sm_RootController.scala 69:23:@84012.4]
  assign io_memStreams_loads_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x474_bits_addr; // @[sm_RootController.scala 69:23:@84011.4]
  assign io_memStreams_loads_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x474_bits_size; // @[sm_RootController.scala 69:23:@84010.4]
  assign io_memStreams_loads_0_data_ready = RootController_kernelRootController_concrete1_io_in_x476_ready; // @[sm_RootController.scala 66:23:@84005.4]
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x669_valid; // @[sm_RootController.scala 65:23:@84001.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x669_bits_addr; // @[sm_RootController.scala 65:23:@84000.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x669_bits_size; // @[sm_RootController.scala 65:23:@83999.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x670_valid; // @[sm_RootController.scala 64:23:@83997.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x670_bits_wdata_0; // @[sm_RootController.scala 64:23:@83996.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x670_bits_wstrb; // @[sm_RootController.scala 64:23:@83995.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x671_ready; // @[sm_RootController.scala 68:23:@84009.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_16 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_17 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_18 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_19 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_20 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_21 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_22 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_23 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_24 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_25 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_26 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_27 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_28 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_29 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_30 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_31 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_32 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_33 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_34 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_35 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_36 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_37 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_38 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_39 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_40 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_41 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_42 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_43 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_44 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_45 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_46 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_47 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_48 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_49 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_50 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_51 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_52 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_53 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_54 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_55 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_56 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_57 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_58 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_59 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_60 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_61 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_62 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_63 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_16 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_17 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_18 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_19 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_20 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_21 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_22 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_23 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_24 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_25 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_26 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_27 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_28 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_29 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_30 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_31 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_32 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_33 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_34 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_35 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_36 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_37 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_38 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_39 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_40 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_41 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_42 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_43 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_44 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_45 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_46 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_47 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_48 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_49 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_50 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_51 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_52 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_53 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_54 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_55 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_56 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_57 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_58 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_59 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_60 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_61 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_62 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_63 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_16 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_17 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_18 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_19 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_20 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_21 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_22 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_23 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_24 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_25 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_26 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_27 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_28 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_29 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_30 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_31 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_32 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_33 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_34 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_35 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_36 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_37 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_38 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_39 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_40 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_41 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_42 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_43 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_44 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_45 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_46 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_47 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_48 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_49 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_50 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_51 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_52 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_53 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_54 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_55 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_56 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_57 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_58 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_59 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_60 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_61 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_62 = 8'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_63 = 8'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = 1'h0;
  assign io_axiStreamsOut_0_TVALID = 1'h0;
  assign io_axiStreamsOut_0_TDATA = 256'h0;
  assign io_axiStreamsOut_0_TSTRB = 32'h0;
  assign io_axiStreamsOut_0_TKEEP = 32'h0;
  assign io_axiStreamsOut_0_TLAST = 1'h0;
  assign io_axiStreamsOut_0_TID = 8'h0;
  assign io_axiStreamsOut_0_TDEST = 8'h0;
  assign io_axiStreamsOut_0_TUSER = 32'h0;
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = io_enable; // @[Instrument.scala 29:62:@84149.4]
  assign io_argOuts_0_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_0_cycs; // @[Instrument.scala 28:61:@84148.4]
  assign io_argOuts_1_port_valid = io_enable; // @[Instrument.scala 31:61:@84151.4]
  assign io_argOuts_1_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_0_iters; // @[Instrument.scala 30:60:@84150.4]
  assign io_argOuts_2_port_valid = io_enable; // @[Instrument.scala 33:62:@84153.4]
  assign io_argOuts_2_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_1_cycs; // @[Instrument.scala 32:61:@84152.4]
  assign io_argOuts_3_port_valid = io_enable; // @[Instrument.scala 35:61:@84155.4]
  assign io_argOuts_3_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_1_iters; // @[Instrument.scala 34:60:@84154.4]
  assign io_argOuts_4_port_valid = io_enable; // @[Instrument.scala 37:62:@84157.4]
  assign io_argOuts_4_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_2_cycs; // @[Instrument.scala 36:61:@84156.4]
  assign io_argOuts_5_port_valid = io_enable; // @[Instrument.scala 39:61:@84159.4]
  assign io_argOuts_5_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_2_iters; // @[Instrument.scala 38:60:@84158.4]
  assign io_argOuts_6_port_valid = io_enable; // @[Instrument.scala 41:63:@84161.4]
  assign io_argOuts_6_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_2_stalls; // @[Instrument.scala 40:62:@84160.4]
  assign io_argOuts_7_port_valid = io_enable; // @[Instrument.scala 43:60:@84163.4]
  assign io_argOuts_7_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_2_idles; // @[Instrument.scala 42:59:@84162.4]
  assign io_argOuts_8_port_valid = io_enable; // @[Instrument.scala 45:62:@84165.4]
  assign io_argOuts_8_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_3_cycs; // @[Instrument.scala 44:61:@84164.4]
  assign io_argOuts_9_port_valid = io_enable; // @[Instrument.scala 47:61:@84167.4]
  assign io_argOuts_9_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_3_iters; // @[Instrument.scala 46:60:@84166.4]
  assign io_argOuts_10_port_valid = io_enable; // @[Instrument.scala 49:62:@84169.4]
  assign io_argOuts_10_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_4_cycs; // @[Instrument.scala 48:61:@84168.4]
  assign io_argOuts_11_port_valid = io_enable; // @[Instrument.scala 51:61:@84171.4]
  assign io_argOuts_11_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_4_iters; // @[Instrument.scala 50:60:@84170.4]
  assign io_argOuts_12_port_valid = io_enable; // @[Instrument.scala 53:63:@84173.4]
  assign io_argOuts_12_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_4_stalls; // @[Instrument.scala 52:62:@84172.4]
  assign io_argOuts_13_port_valid = io_enable; // @[Instrument.scala 55:60:@84175.4]
  assign io_argOuts_13_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_4_idles; // @[Instrument.scala 54:59:@84174.4]
  assign io_argOuts_14_port_valid = io_enable; // @[Instrument.scala 57:62:@84177.4]
  assign io_argOuts_14_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_5_cycs; // @[Instrument.scala 56:61:@84176.4]
  assign io_argOuts_15_port_valid = io_enable; // @[Instrument.scala 59:61:@84179.4]
  assign io_argOuts_15_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_5_iters; // @[Instrument.scala 58:60:@84178.4]
  assign io_argOuts_16_port_valid = io_enable; // @[Instrument.scala 61:63:@84181.4]
  assign io_argOuts_16_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_5_stalls; // @[Instrument.scala 60:62:@84180.4]
  assign io_argOuts_17_port_valid = io_enable; // @[Instrument.scala 63:60:@84183.4]
  assign io_argOuts_17_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_5_idles; // @[Instrument.scala 62:59:@84182.4]
  assign io_argOuts_18_port_valid = io_enable; // @[Instrument.scala 65:62:@84185.4]
  assign io_argOuts_18_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_6_cycs; // @[Instrument.scala 64:61:@84184.4]
  assign io_argOuts_19_port_valid = io_enable; // @[Instrument.scala 67:61:@84187.4]
  assign io_argOuts_19_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_6_iters; // @[Instrument.scala 66:60:@84186.4]
  assign io_argOuts_20_port_valid = io_enable; // @[Instrument.scala 69:62:@84189.4]
  assign io_argOuts_20_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_7_cycs; // @[Instrument.scala 68:61:@84188.4]
  assign io_argOuts_21_port_valid = io_enable; // @[Instrument.scala 71:61:@84191.4]
  assign io_argOuts_21_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_7_iters; // @[Instrument.scala 70:60:@84190.4]
  assign io_argOuts_22_port_valid = io_enable; // @[Instrument.scala 73:62:@84193.4]
  assign io_argOuts_22_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_8_cycs; // @[Instrument.scala 72:61:@84192.4]
  assign io_argOuts_23_port_valid = io_enable; // @[Instrument.scala 75:61:@84195.4]
  assign io_argOuts_23_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_8_iters; // @[Instrument.scala 74:60:@84194.4]
  assign io_argOuts_24_port_valid = io_enable; // @[Instrument.scala 83:62:@84197.4]
  assign io_argOuts_24_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_9_cycs; // @[Instrument.scala 76:61:@84196.4]
  assign io_argOuts_25_port_valid = io_enable; // @[Instrument.scala 85:61:@84199.4]
  assign io_argOuts_25_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_9_iters; // @[Instrument.scala 84:60:@84198.4]
  assign io_argOuts_26_port_valid = io_enable; // @[Instrument.scala 87:62:@84201.4]
  assign io_argOuts_26_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_10_cycs; // @[Instrument.scala 86:61:@84200.4]
  assign io_argOuts_27_port_valid = io_enable; // @[Instrument.scala 89:61:@84203.4]
  assign io_argOuts_27_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_10_iters; // @[Instrument.scala 88:60:@84202.4]
  assign io_argOuts_28_port_valid = io_enable; // @[Instrument.scala 91:62:@84205.4]
  assign io_argOuts_28_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_11_cycs; // @[Instrument.scala 90:61:@84204.4]
  assign io_argOuts_29_port_valid = io_enable; // @[Instrument.scala 93:61:@84207.4]
  assign io_argOuts_29_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_11_iters; // @[Instrument.scala 92:60:@84206.4]
  assign io_argOuts_30_port_valid = io_enable; // @[Instrument.scala 95:62:@84209.4]
  assign io_argOuts_30_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_12_cycs; // @[Instrument.scala 94:61:@84208.4]
  assign io_argOuts_31_port_valid = io_enable; // @[Instrument.scala 97:61:@84211.4]
  assign io_argOuts_31_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_12_iters; // @[Instrument.scala 96:60:@84210.4]
  assign io_argOuts_32_port_valid = io_enable; // @[Instrument.scala 99:62:@84213.4]
  assign io_argOuts_32_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_13_cycs; // @[Instrument.scala 98:61:@84212.4]
  assign io_argOuts_33_port_valid = io_enable; // @[Instrument.scala 101:61:@84215.4]
  assign io_argOuts_33_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_13_iters; // @[Instrument.scala 100:60:@84214.4]
  assign io_argOuts_34_port_valid = io_enable; // @[Instrument.scala 103:62:@84217.4]
  assign io_argOuts_34_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_14_cycs; // @[Instrument.scala 102:61:@84216.4]
  assign io_argOuts_35_port_valid = io_enable; // @[Instrument.scala 105:61:@84219.4]
  assign io_argOuts_35_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_14_iters; // @[Instrument.scala 104:60:@84218.4]
  assign io_argOuts_36_port_valid = io_enable; // @[Instrument.scala 107:62:@84221.4]
  assign io_argOuts_36_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_15_cycs; // @[Instrument.scala 106:61:@84220.4]
  assign io_argOuts_37_port_valid = io_enable; // @[Instrument.scala 109:61:@84223.4]
  assign io_argOuts_37_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_15_iters; // @[Instrument.scala 108:60:@84222.4]
  assign io_argOuts_38_port_valid = io_enable; // @[Instrument.scala 111:62:@84225.4]
  assign io_argOuts_38_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_16_cycs; // @[Instrument.scala 110:61:@84224.4]
  assign io_argOuts_39_port_valid = io_enable; // @[Instrument.scala 113:61:@84227.4]
  assign io_argOuts_39_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_16_iters; // @[Instrument.scala 112:60:@84226.4]
  assign io_argOuts_40_port_valid = io_enable; // @[Instrument.scala 115:62:@84229.4]
  assign io_argOuts_40_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_17_cycs; // @[Instrument.scala 114:61:@84228.4]
  assign io_argOuts_41_port_valid = io_enable; // @[Instrument.scala 117:61:@84231.4]
  assign io_argOuts_41_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_17_iters; // @[Instrument.scala 116:60:@84230.4]
  assign io_argOuts_42_port_valid = io_enable; // @[Instrument.scala 119:62:@84233.4]
  assign io_argOuts_42_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_18_cycs; // @[Instrument.scala 118:61:@84232.4]
  assign io_argOuts_43_port_valid = io_enable; // @[Instrument.scala 121:61:@84235.4]
  assign io_argOuts_43_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_18_iters; // @[Instrument.scala 120:60:@84234.4]
  assign io_argOuts_44_port_valid = io_enable; // @[Instrument.scala 123:62:@84237.4]
  assign io_argOuts_44_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_19_cycs; // @[Instrument.scala 122:61:@84236.4]
  assign io_argOuts_45_port_valid = io_enable; // @[Instrument.scala 125:61:@84239.4]
  assign io_argOuts_45_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_19_iters; // @[Instrument.scala 124:60:@84238.4]
  assign io_argOuts_46_port_valid = io_enable; // @[Instrument.scala 127:62:@84241.4]
  assign io_argOuts_46_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_20_cycs; // @[Instrument.scala 126:61:@84240.4]
  assign io_argOuts_47_port_valid = io_enable; // @[Instrument.scala 129:61:@84243.4]
  assign io_argOuts_47_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_20_iters; // @[Instrument.scala 128:60:@84242.4]
  assign io_argOuts_48_port_valid = io_enable; // @[Instrument.scala 131:62:@84245.4]
  assign io_argOuts_48_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_21_cycs; // @[Instrument.scala 130:61:@84244.4]
  assign io_argOuts_49_port_valid = io_enable; // @[Instrument.scala 139:61:@84247.4]
  assign io_argOuts_49_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_21_iters; // @[Instrument.scala 138:60:@84246.4]
  assign io_argOuts_50_port_valid = io_enable; // @[Instrument.scala 141:63:@84249.4]
  assign io_argOuts_50_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_21_stalls; // @[Instrument.scala 140:62:@84248.4]
  assign io_argOuts_51_port_valid = io_enable; // @[Instrument.scala 143:60:@84251.4]
  assign io_argOuts_51_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_21_idles; // @[Instrument.scala 142:59:@84250.4]
  assign io_argOuts_52_port_valid = io_enable; // @[Instrument.scala 145:62:@84253.4]
  assign io_argOuts_52_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_22_cycs; // @[Instrument.scala 144:61:@84252.4]
  assign io_argOuts_53_port_valid = io_enable; // @[Instrument.scala 147:61:@84255.4]
  assign io_argOuts_53_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_22_iters; // @[Instrument.scala 146:60:@84254.4]
  assign io_argOuts_54_port_valid = io_enable; // @[Instrument.scala 149:63:@84257.4]
  assign io_argOuts_54_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_22_stalls; // @[Instrument.scala 148:62:@84256.4]
  assign io_argOuts_55_port_valid = io_enable; // @[Instrument.scala 151:60:@84259.4]
  assign io_argOuts_55_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_22_idles; // @[Instrument.scala 150:59:@84258.4]
  assign io_argOuts_56_port_valid = io_enable; // @[Instrument.scala 153:62:@84261.4]
  assign io_argOuts_56_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_23_cycs; // @[Instrument.scala 152:61:@84260.4]
  assign io_argOuts_57_port_valid = io_enable; // @[Instrument.scala 155:61:@84263.4]
  assign io_argOuts_57_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_23_iters; // @[Instrument.scala 154:60:@84262.4]
  assign io_argOuts_58_port_valid = io_enable; // @[Instrument.scala 157:63:@84265.4]
  assign io_argOuts_58_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_23_stalls; // @[Instrument.scala 156:62:@84264.4]
  assign io_argOuts_59_port_valid = io_enable; // @[Instrument.scala 159:60:@84267.4]
  assign io_argOuts_59_port_bits = RootController_kernelRootController_concrete1_io_in_instrctrs_23_idles; // @[Instrument.scala 158:59:@84266.4]
  assign SingleCounter_clock = clock; // @[:@83526.4]
  assign SingleCounter_reset = reset; // @[:@83527.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 43:79:@83541.4]
  assign RetimeWrapper_clock = clock; // @[:@83544.4]
  assign RetimeWrapper_reset = reset; // @[:@83545.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@83547.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@83546.4]
  assign SRFF_clock = clock; // @[:@83673.4]
  assign SRFF_reset = reset; // @[:@83674.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 65:29:@84147.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 54:31:@83778.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 55:36:@83779.4]
  assign RootController_sm_clock = clock; // @[:@83722.4]
  assign RootController_sm_reset = reset; // @[:@83723.4]
  assign RootController_sm_io_enable = _T_1376 & _T_1377; // @[Main.scala 53:33:@83777.4 SpatialBlocks.scala 139:18:@83822.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 133:15:@83816.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_1394; // @[Main.scala 57:34:@83785.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@83809.4]
  assign RootController_sm_io_doneIn_1 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:72:@83810.4]
  assign RootController_sm_io_doneIn_2 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:72:@83811.4]
  assign RetimeWrapper_1_clock = clock; // @[:@83764.4]
  assign RetimeWrapper_1_reset = reset; // @[:@83765.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@83767.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@83766.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@83838.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@83839.4]
  assign RootController_kernelRootController_concrete1_io_in_x468_A_dram_number = io_argIns_0; // @[sm_RootController.scala 63:30:@83994.4]
  assign RootController_kernelRootController_concrete1_io_in_x670_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 64:23:@83998.4]
  assign RootController_kernelRootController_concrete1_io_in_x669_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 65:23:@84002.4]
  assign RootController_kernelRootController_concrete1_io_in_x476_valid = io_memStreams_loads_0_data_valid; // @[sm_RootController.scala 66:23:@84004.4]
  assign RootController_kernelRootController_concrete1_io_in_x476_bits_rdata_0 = io_memStreams_loads_0_data_bits_rdata_0; // @[sm_RootController.scala 66:23:@84003.4]
  assign RootController_kernelRootController_concrete1_io_in_x470_out_host_number = io_argIns_1; // @[sm_RootController.scala 67:32:@84006.4]
  assign RootController_kernelRootController_concrete1_io_in_x671_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 68:23:@84008.4]
  assign RootController_kernelRootController_concrete1_io_in_x474_ready = io_memStreams_loads_0_cmd_ready; // @[sm_RootController.scala 69:23:@84013.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_done = RootController_sm_io_done; // @[sm_RootController.scala 131:22:@84135.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_baseEn = _T_1376 & _T_1377; // @[sm_RootController.scala 131:22:@84127.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 131:22:@84122.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1 = RootController_sm_io_enableOut_1; // @[sm_RootController.scala 131:22:@84123.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_2 = RootController_sm_io_enableOut_2; // @[sm_RootController.scala 131:22:@84124.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 131:22:@84116.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1 = RootController_sm_io_childAck_1; // @[sm_RootController.scala 131:22:@84117.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_2 = RootController_sm_io_childAck_2; // @[sm_RootController.scala 131:22:@84118.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 130:18:@84110.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1394 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1394 <= 1'h0;
    end else begin
      _T_1394 <= _T_1391;
    end
  end
endmodule
module Counter( // @[:@84269.2]
  input        clock, // @[:@84270.4]
  input        reset, // @[:@84271.4]
  input        io_reset, // @[:@84272.4]
  input        io_enable, // @[:@84272.4]
  input  [5:0] io_stride, // @[:@84272.4]
  output [5:0] io_out, // @[:@84272.4]
  output [5:0] io_next // @[:@84272.4]
);
  reg [5:0] count; // @[Counter.scala 15:22:@84274.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_17; // @[Counter.scala 17:24:@84275.4]
  wire [5:0] newCount; // @[Counter.scala 17:24:@84276.4]
  wire [5:0] _GEN_0; // @[Counter.scala 21:26:@84281.6]
  wire [5:0] _GEN_1; // @[Counter.scala 19:18:@84277.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@84275.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@84276.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@84281.6]
  assign _GEN_1 = io_reset ? 6'h0 : _GEN_0; // @[Counter.scala 19:18:@84277.4]
  assign io_out = count; // @[Counter.scala 25:10:@84284.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@84285.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 6'h0;
    end else begin
      if (io_reset) begin
        count <= 6'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_76( // @[:@84321.2]
  input         clock, // @[:@84322.4]
  input  [5:0]  io_raddr, // @[:@84324.4]
  input         io_wen, // @[:@84324.4]
  input  [5:0]  io_waddr, // @[:@84324.4]
  input  [63:0] io_wdata_addr, // @[:@84324.4]
  input  [31:0] io_wdata_size, // @[:@84324.4]
  output [63:0] io_rdata_addr, // @[:@84324.4]
  output [31:0] io_rdata_size, // @[:@84324.4]
  input         io_backpressure // @[:@84324.4]
);
  wire [95:0] SRAMVerilogSim_rdata; // @[SRAM.scala 187:23:@84326.4]
  wire [95:0] SRAMVerilogSim_wdata; // @[SRAM.scala 187:23:@84326.4]
  wire  SRAMVerilogSim_backpressure; // @[SRAM.scala 187:23:@84326.4]
  wire  SRAMVerilogSim_wen; // @[SRAM.scala 187:23:@84326.4]
  wire  SRAMVerilogSim_waddrEn; // @[SRAM.scala 187:23:@84326.4]
  wire  SRAMVerilogSim_raddrEn; // @[SRAM.scala 187:23:@84326.4]
  wire [5:0] SRAMVerilogSim_waddr; // @[SRAM.scala 187:23:@84326.4]
  wire [5:0] SRAMVerilogSim_raddr; // @[SRAM.scala 187:23:@84326.4]
  wire  SRAMVerilogSim_clk; // @[SRAM.scala 187:23:@84326.4]
  wire [95:0] _T_23; // @[:@84346.4 :@84347.4]
  SRAMVerilogSim #(.DWIDTH(96), .WORDS(64), .AWIDTH(6)) SRAMVerilogSim ( // @[SRAM.scala 187:23:@84326.4]
    .rdata(SRAMVerilogSim_rdata),
    .wdata(SRAMVerilogSim_wdata),
    .backpressure(SRAMVerilogSim_backpressure),
    .wen(SRAMVerilogSim_wen),
    .waddrEn(SRAMVerilogSim_waddrEn),
    .raddrEn(SRAMVerilogSim_raddrEn),
    .waddr(SRAMVerilogSim_waddr),
    .raddr(SRAMVerilogSim_raddr),
    .clk(SRAMVerilogSim_clk)
  );
  assign _T_23 = SRAMVerilogSim_rdata; // @[:@84346.4 :@84347.4]
  assign io_rdata_addr = _T_23[95:32]; // @[SRAM.scala 197:16:@84353.4]
  assign io_rdata_size = _T_23[31:0]; // @[SRAM.scala 197:16:@84352.4]
  assign SRAMVerilogSim_wdata = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 192:20:@84341.4]
  assign SRAMVerilogSim_backpressure = io_backpressure; // @[SRAM.scala 193:27:@84342.4]
  assign SRAMVerilogSim_wen = io_wen; // @[SRAM.scala 190:18:@84338.4]
  assign SRAMVerilogSim_waddrEn = 1'h1; // @[SRAM.scala 195:22:@84344.4]
  assign SRAMVerilogSim_raddrEn = 1'h1; // @[SRAM.scala 194:22:@84343.4]
  assign SRAMVerilogSim_waddr = io_waddr; // @[SRAM.scala 191:20:@84339.4]
  assign SRAMVerilogSim_raddr = io_raddr; // @[SRAM.scala 189:20:@84337.4]
  assign SRAMVerilogSim_clk = clock; // @[SRAM.scala 188:18:@84336.4]
endmodule
module FIFO( // @[:@84355.2]
  input         clock, // @[:@84356.4]
  input         reset, // @[:@84357.4]
  output        io_in_ready, // @[:@84358.4]
  input         io_in_valid, // @[:@84358.4]
  input  [63:0] io_in_bits_addr, // @[:@84358.4]
  input  [31:0] io_in_bits_size, // @[:@84358.4]
  input         io_out_ready, // @[:@84358.4]
  output        io_out_valid, // @[:@84358.4]
  output [63:0] io_out_bits_addr, // @[:@84358.4]
  output [31:0] io_out_bits_size // @[:@84358.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@84754.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@84754.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@84754.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@84754.4]
  wire [5:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@84754.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@84754.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@84754.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@84764.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@84764.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@84764.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@84764.4]
  wire [5:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@84764.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@84764.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@84764.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@84779.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@84779.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@84779.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@84779.4]
  wire [63:0] SRAM_io_wdata_addr; // @[FIFO.scala 73:19:@84779.4]
  wire [31:0] SRAM_io_wdata_size; // @[FIFO.scala 73:19:@84779.4]
  wire [63:0] SRAM_io_rdata_addr; // @[FIFO.scala 73:19:@84779.4]
  wire [31:0] SRAM_io_rdata_size; // @[FIFO.scala 73:19:@84779.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@84779.4]
  wire  writeEn; // @[FIFO.scala 30:29:@84752.4]
  wire  readEn; // @[FIFO.scala 31:29:@84753.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@84774.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@84775.4]
  wire  _T_824; // @[FIFO.scala 45:27:@84776.4]
  wire  empty; // @[FIFO.scala 45:24:@84777.4]
  wire  full; // @[FIFO.scala 46:23:@84778.4]
  wire  _T_827; // @[FIFO.scala 83:17:@84791.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@84792.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@84754.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@84764.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_76 SRAM ( // @[FIFO.scala 73:19:@84779.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata_addr(SRAM_io_wdata_addr),
    .io_wdata_size(SRAM_io_wdata_size),
    .io_rdata_addr(SRAM_io_rdata_addr),
    .io_rdata_size(SRAM_io_rdata_size),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@84752.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@84753.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@84775.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@84776.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@84777.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@84778.4]
  assign _T_827 = writeEn != readEn; // @[FIFO.scala 83:17:@84791.4]
  assign _GEN_0 = _T_827 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@84792.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@84798.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@84796.4]
  assign io_out_bits_addr = SRAM_io_rdata_addr; // @[FIFO.scala 79:17:@84789.4]
  assign io_out_bits_size = SRAM_io_rdata_size; // @[FIFO.scala 79:17:@84788.4]
  assign enqCounter_clock = clock; // @[:@84755.4]
  assign enqCounter_reset = reset; // @[:@84756.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@84762.4]
  assign enqCounter_io_stride = 6'h1; // @[FIFO.scala 37:24:@84763.4]
  assign deqCounter_clock = clock; // @[:@84765.4]
  assign deqCounter_reset = reset; // @[:@84766.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@84772.4]
  assign deqCounter_io_stride = 6'h1; // @[FIFO.scala 41:24:@84773.4]
  assign SRAM_clock = clock; // @[:@84780.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@84783.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@84784.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@84785.4]
  assign SRAM_io_wdata_addr = io_in_bits_addr; // @[FIFO.scala 78:16:@84787.4]
  assign SRAM_io_wdata_size = io_in_bits_size; // @[FIFO.scala 78:16:@84786.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@84790.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_827) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module Counter_2( // @[:@84800.2]
  input        clock, // @[:@84801.4]
  input        reset, // @[:@84802.4]
  input        io_reset, // @[:@84803.4]
  input        io_enable, // @[:@84803.4]
  input  [3:0] io_stride, // @[:@84803.4]
  output [3:0] io_out // @[:@84803.4]
);
  reg [3:0] count; // @[Counter.scala 15:22:@84805.4]
  reg [31:0] _RAND_0;
  wire [4:0] _T_17; // @[Counter.scala 17:24:@84806.4]
  wire [3:0] newCount; // @[Counter.scala 17:24:@84807.4]
  wire [3:0] _GEN_0; // @[Counter.scala 21:26:@84812.6]
  wire [3:0] _GEN_1; // @[Counter.scala 19:18:@84808.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@84806.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@84807.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@84812.6]
  assign _GEN_1 = io_reset ? 4'h0 : _GEN_0; // @[Counter.scala 19:18:@84808.4]
  assign io_out = count; // @[Counter.scala 25:10:@84815.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 4'h0;
    end else begin
      if (io_reset) begin
        count <= 4'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module Counter_4( // @[:@84836.2]
  input        clock, // @[:@84837.4]
  input        reset, // @[:@84838.4]
  input        io_reset, // @[:@84839.4]
  input        io_enable, // @[:@84839.4]
  input  [1:0] io_stride, // @[:@84839.4]
  output [1:0] io_out, // @[:@84839.4]
  output [1:0] io_next // @[:@84839.4]
);
  reg [1:0] count; // @[Counter.scala 15:22:@84841.4]
  reg [31:0] _RAND_0;
  wire [2:0] _T_17; // @[Counter.scala 17:24:@84842.4]
  wire [1:0] newCount; // @[Counter.scala 17:24:@84843.4]
  wire [1:0] _GEN_0; // @[Counter.scala 21:26:@84848.6]
  wire [1:0] _GEN_1; // @[Counter.scala 19:18:@84844.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@84842.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@84843.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@84848.6]
  assign _GEN_1 = io_reset ? 2'h0 : _GEN_0; // @[Counter.scala 19:18:@84844.4]
  assign io_out = count; // @[Counter.scala 25:10:@84851.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@84852.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 2'h0;
    end else begin
      if (io_reset) begin
        count <= 2'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_77( // @[:@84888.2]
  input         clock, // @[:@84889.4]
  input  [1:0]  io_raddr, // @[:@84891.4]
  input         io_wen, // @[:@84891.4]
  input  [1:0]  io_waddr, // @[:@84891.4]
  input  [31:0] io_wdata, // @[:@84891.4]
  output [31:0] io_rdata, // @[:@84891.4]
  input         io_backpressure // @[:@84891.4]
);
  wire [31:0] SRAMVerilogSim_rdata; // @[SRAM.scala 187:23:@84893.4]
  wire [31:0] SRAMVerilogSim_wdata; // @[SRAM.scala 187:23:@84893.4]
  wire  SRAMVerilogSim_backpressure; // @[SRAM.scala 187:23:@84893.4]
  wire  SRAMVerilogSim_wen; // @[SRAM.scala 187:23:@84893.4]
  wire  SRAMVerilogSim_waddrEn; // @[SRAM.scala 187:23:@84893.4]
  wire  SRAMVerilogSim_raddrEn; // @[SRAM.scala 187:23:@84893.4]
  wire [1:0] SRAMVerilogSim_waddr; // @[SRAM.scala 187:23:@84893.4]
  wire [1:0] SRAMVerilogSim_raddr; // @[SRAM.scala 187:23:@84893.4]
  wire  SRAMVerilogSim_clk; // @[SRAM.scala 187:23:@84893.4]
  SRAMVerilogSim #(.DWIDTH(32), .WORDS(4), .AWIDTH(2)) SRAMVerilogSim ( // @[SRAM.scala 187:23:@84893.4]
    .rdata(SRAMVerilogSim_rdata),
    .wdata(SRAMVerilogSim_wdata),
    .backpressure(SRAMVerilogSim_backpressure),
    .wen(SRAMVerilogSim_wen),
    .waddrEn(SRAMVerilogSim_waddrEn),
    .raddrEn(SRAMVerilogSim_raddrEn),
    .waddr(SRAMVerilogSim_waddr),
    .raddr(SRAMVerilogSim_raddr),
    .clk(SRAMVerilogSim_clk)
  );
  assign io_rdata = SRAMVerilogSim_rdata; // @[SRAM.scala 197:16:@84913.4]
  assign SRAMVerilogSim_wdata = io_wdata; // @[SRAM.scala 192:20:@84907.4]
  assign SRAMVerilogSim_backpressure = io_backpressure; // @[SRAM.scala 193:27:@84908.4]
  assign SRAMVerilogSim_wen = io_wen; // @[SRAM.scala 190:18:@84905.4]
  assign SRAMVerilogSim_waddrEn = 1'h1; // @[SRAM.scala 195:22:@84910.4]
  assign SRAMVerilogSim_raddrEn = 1'h1; // @[SRAM.scala 194:22:@84909.4]
  assign SRAMVerilogSim_waddr = io_waddr; // @[SRAM.scala 191:20:@84906.4]
  assign SRAMVerilogSim_raddr = io_raddr; // @[SRAM.scala 189:20:@84904.4]
  assign SRAMVerilogSim_clk = clock; // @[SRAM.scala 188:18:@84903.4]
endmodule
module FIFO_1( // @[:@84915.2]
  input         clock, // @[:@84916.4]
  input         reset, // @[:@84917.4]
  output        io_in_ready, // @[:@84918.4]
  input         io_in_valid, // @[:@84918.4]
  input  [31:0] io_in_bits, // @[:@84918.4]
  input         io_out_ready, // @[:@84918.4]
  output        io_out_valid, // @[:@84918.4]
  output [31:0] io_out_bits // @[:@84918.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@84944.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@84944.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@84944.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@84944.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@84944.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@84944.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@84944.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@84954.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@84954.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@84954.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@84954.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@84954.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@84954.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@84954.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@84969.4]
  wire [1:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@84969.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@84969.4]
  wire [1:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@84969.4]
  wire [31:0] SRAM_io_wdata; // @[FIFO.scala 73:19:@84969.4]
  wire [31:0] SRAM_io_rdata; // @[FIFO.scala 73:19:@84969.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@84969.4]
  wire  writeEn; // @[FIFO.scala 30:29:@84942.4]
  wire  readEn; // @[FIFO.scala 31:29:@84943.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@84964.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@84965.4]
  wire  _T_104; // @[FIFO.scala 45:27:@84966.4]
  wire  empty; // @[FIFO.scala 45:24:@84967.4]
  wire  full; // @[FIFO.scala 46:23:@84968.4]
  wire  _T_107; // @[FIFO.scala 83:17:@84979.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@84980.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@84944.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@84954.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_77 SRAM ( // @[FIFO.scala 73:19:@84969.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@84942.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@84943.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@84965.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@84966.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@84967.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@84968.4]
  assign _T_107 = writeEn != readEn; // @[FIFO.scala 83:17:@84979.4]
  assign _GEN_0 = _T_107 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@84980.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@84986.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@84984.4]
  assign io_out_bits = SRAM_io_rdata; // @[FIFO.scala 79:17:@84977.4]
  assign enqCounter_clock = clock; // @[:@84945.4]
  assign enqCounter_reset = reset; // @[:@84946.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@84952.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@84953.4]
  assign deqCounter_clock = clock; // @[:@84955.4]
  assign deqCounter_reset = reset; // @[:@84956.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@84962.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@84963.4]
  assign SRAM_clock = clock; // @[:@84970.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@84973.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@84974.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@84975.4]
  assign SRAM_io_wdata = io_in_bits; // @[FIFO.scala 78:16:@84976.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@84978.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_107) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec( // @[:@87268.2]
  input         clock, // @[:@87269.4]
  input         reset, // @[:@87270.4]
  output        io_in_ready, // @[:@87271.4]
  input         io_in_valid, // @[:@87271.4]
  input  [31:0] io_in_bits_0, // @[:@87271.4]
  input  [31:0] io_in_bits_1, // @[:@87271.4]
  input  [31:0] io_in_bits_2, // @[:@87271.4]
  input  [31:0] io_in_bits_3, // @[:@87271.4]
  input  [31:0] io_in_bits_4, // @[:@87271.4]
  input  [31:0] io_in_bits_5, // @[:@87271.4]
  input  [31:0] io_in_bits_6, // @[:@87271.4]
  input  [31:0] io_in_bits_7, // @[:@87271.4]
  input  [31:0] io_in_bits_8, // @[:@87271.4]
  input  [31:0] io_in_bits_9, // @[:@87271.4]
  input  [31:0] io_in_bits_10, // @[:@87271.4]
  input  [31:0] io_in_bits_11, // @[:@87271.4]
  input  [31:0] io_in_bits_12, // @[:@87271.4]
  input  [31:0] io_in_bits_13, // @[:@87271.4]
  input  [31:0] io_in_bits_14, // @[:@87271.4]
  input  [31:0] io_in_bits_15, // @[:@87271.4]
  input         io_out_ready, // @[:@87271.4]
  output        io_out_valid, // @[:@87271.4]
  output [31:0] io_out_bits_0, // @[:@87271.4]
  output [31:0] io_out_bits_1, // @[:@87271.4]
  output [31:0] io_out_bits_2, // @[:@87271.4]
  output [31:0] io_out_bits_3, // @[:@87271.4]
  output [31:0] io_out_bits_4, // @[:@87271.4]
  output [31:0] io_out_bits_5, // @[:@87271.4]
  output [31:0] io_out_bits_6, // @[:@87271.4]
  output [31:0] io_out_bits_7, // @[:@87271.4]
  output [31:0] io_out_bits_8, // @[:@87271.4]
  output [31:0] io_out_bits_9, // @[:@87271.4]
  output [31:0] io_out_bits_10, // @[:@87271.4]
  output [31:0] io_out_bits_11, // @[:@87271.4]
  output [31:0] io_out_bits_12, // @[:@87271.4]
  output [31:0] io_out_bits_13, // @[:@87271.4]
  output [31:0] io_out_bits_14, // @[:@87271.4]
  output [31:0] io_out_bits_15, // @[:@87271.4]
  input         io_chainEnq, // @[:@87271.4]
  input         io_chainDeq // @[:@87271.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@87275.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@87275.4]
  wire  enqCounter_io_reset; // @[FIFOVec.scala 24:26:@87275.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@87275.4]
  wire [3:0] enqCounter_io_stride; // @[FIFOVec.scala 24:26:@87275.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@87275.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@87286.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@87286.4]
  wire  deqCounter_io_reset; // @[FIFOVec.scala 28:26:@87286.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@87286.4]
  wire [3:0] deqCounter_io_stride; // @[FIFOVec.scala 28:26:@87286.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@87286.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@87299.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@87299.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@87299.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@87299.4]
  wire [31:0] fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@87299.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@87299.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@87299.4]
  wire [31:0] fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@87299.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@87334.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@87334.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@87334.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@87334.4]
  wire [31:0] fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@87334.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@87334.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@87334.4]
  wire [31:0] fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@87334.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@87369.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@87369.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@87369.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@87369.4]
  wire [31:0] fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@87369.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@87369.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@87369.4]
  wire [31:0] fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@87369.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@87404.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@87404.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@87404.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@87404.4]
  wire [31:0] fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@87404.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@87404.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@87404.4]
  wire [31:0] fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@87404.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@87439.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@87439.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@87439.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@87439.4]
  wire [31:0] fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@87439.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@87439.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@87439.4]
  wire [31:0] fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@87439.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@87474.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@87474.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@87474.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@87474.4]
  wire [31:0] fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@87474.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@87474.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@87474.4]
  wire [31:0] fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@87474.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@87509.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@87509.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@87509.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@87509.4]
  wire [31:0] fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@87509.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@87509.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@87509.4]
  wire [31:0] fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@87509.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@87544.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@87544.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@87544.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@87544.4]
  wire [31:0] fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@87544.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@87544.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@87544.4]
  wire [31:0] fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@87544.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@87579.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@87579.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@87579.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@87579.4]
  wire [31:0] fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@87579.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@87579.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@87579.4]
  wire [31:0] fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@87579.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@87614.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@87614.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@87614.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@87614.4]
  wire [31:0] fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@87614.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@87614.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@87614.4]
  wire [31:0] fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@87614.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@87649.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@87649.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@87649.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@87649.4]
  wire [31:0] fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@87649.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@87649.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@87649.4]
  wire [31:0] fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@87649.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@87684.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@87684.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@87684.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@87684.4]
  wire [31:0] fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@87684.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@87684.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@87684.4]
  wire [31:0] fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@87684.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@87719.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@87719.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@87719.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@87719.4]
  wire [31:0] fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@87719.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@87719.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@87719.4]
  wire [31:0] fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@87719.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@87754.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@87754.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@87754.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@87754.4]
  wire [31:0] fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@87754.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@87754.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@87754.4]
  wire [31:0] fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@87754.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@87789.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@87789.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@87789.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@87789.4]
  wire [31:0] fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@87789.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@87789.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@87789.4]
  wire [31:0] fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@87789.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@87824.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@87824.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@87824.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@87824.4]
  wire [31:0] fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@87824.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@87824.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@87824.4]
  wire [31:0] fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@87824.4]
  wire  readEn; // @[FIFOVec.scala 20:29:@87273.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@87274.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@87297.4]
  wire [15:0] deqDecoder; // @[OneHot.scala 45:35:@87298.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@87324.4]
  wire  _T_151; // @[FIFOVec.scala 42:25:@87325.4]
  wire  _T_154; // @[FIFOVec.scala 44:50:@87330.4]
  wire  _T_156; // @[FIFOVec.scala 44:26:@87331.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@87359.4]
  wire  _T_160; // @[FIFOVec.scala 42:25:@87360.4]
  wire  _T_163; // @[FIFOVec.scala 44:50:@87365.4]
  wire  _T_165; // @[FIFOVec.scala 44:26:@87366.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@87394.4]
  wire  _T_169; // @[FIFOVec.scala 42:25:@87395.4]
  wire  _T_172; // @[FIFOVec.scala 44:50:@87400.4]
  wire  _T_174; // @[FIFOVec.scala 44:26:@87401.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@87429.4]
  wire  _T_178; // @[FIFOVec.scala 42:25:@87430.4]
  wire  _T_181; // @[FIFOVec.scala 44:50:@87435.4]
  wire  _T_183; // @[FIFOVec.scala 44:26:@87436.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@87464.4]
  wire  _T_187; // @[FIFOVec.scala 42:25:@87465.4]
  wire  _T_190; // @[FIFOVec.scala 44:50:@87470.4]
  wire  _T_192; // @[FIFOVec.scala 44:26:@87471.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@87499.4]
  wire  _T_196; // @[FIFOVec.scala 42:25:@87500.4]
  wire  _T_199; // @[FIFOVec.scala 44:50:@87505.4]
  wire  _T_201; // @[FIFOVec.scala 44:26:@87506.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@87534.4]
  wire  _T_205; // @[FIFOVec.scala 42:25:@87535.4]
  wire  _T_208; // @[FIFOVec.scala 44:50:@87540.4]
  wire  _T_210; // @[FIFOVec.scala 44:26:@87541.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@87569.4]
  wire  _T_214; // @[FIFOVec.scala 42:25:@87570.4]
  wire  _T_217; // @[FIFOVec.scala 44:50:@87575.4]
  wire  _T_219; // @[FIFOVec.scala 44:26:@87576.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@87604.4]
  wire  _T_223; // @[FIFOVec.scala 42:25:@87605.4]
  wire  _T_226; // @[FIFOVec.scala 44:50:@87610.4]
  wire  _T_228; // @[FIFOVec.scala 44:26:@87611.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@87639.4]
  wire  _T_232; // @[FIFOVec.scala 42:25:@87640.4]
  wire  _T_235; // @[FIFOVec.scala 44:50:@87645.4]
  wire  _T_237; // @[FIFOVec.scala 44:26:@87646.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@87674.4]
  wire  _T_241; // @[FIFOVec.scala 42:25:@87675.4]
  wire  _T_244; // @[FIFOVec.scala 44:50:@87680.4]
  wire  _T_246; // @[FIFOVec.scala 44:26:@87681.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@87709.4]
  wire  _T_250; // @[FIFOVec.scala 42:25:@87710.4]
  wire  _T_253; // @[FIFOVec.scala 44:50:@87715.4]
  wire  _T_255; // @[FIFOVec.scala 44:26:@87716.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@87744.4]
  wire  _T_259; // @[FIFOVec.scala 42:25:@87745.4]
  wire  _T_262; // @[FIFOVec.scala 44:50:@87750.4]
  wire  _T_264; // @[FIFOVec.scala 44:26:@87751.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@87779.4]
  wire  _T_268; // @[FIFOVec.scala 42:25:@87780.4]
  wire  _T_271; // @[FIFOVec.scala 44:50:@87785.4]
  wire  _T_273; // @[FIFOVec.scala 44:26:@87786.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@87814.4]
  wire  _T_277; // @[FIFOVec.scala 42:25:@87815.4]
  wire  _T_280; // @[FIFOVec.scala 44:50:@87820.4]
  wire  _T_282; // @[FIFOVec.scala 44:26:@87821.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@87849.4]
  wire  _T_286; // @[FIFOVec.scala 42:25:@87850.4]
  wire  _T_289; // @[FIFOVec.scala 44:50:@87855.4]
  wire  _T_291; // @[FIFOVec.scala 44:26:@87856.4]
  wire  _T_316; // @[FIFOVec.scala 49:90:@87876.4]
  wire  _T_317; // @[FIFOVec.scala 49:90:@87877.4]
  wire  _T_318; // @[FIFOVec.scala 49:90:@87878.4]
  wire  _T_319; // @[FIFOVec.scala 49:90:@87879.4]
  wire  _T_320; // @[FIFOVec.scala 49:90:@87880.4]
  wire  _T_321; // @[FIFOVec.scala 49:90:@87881.4]
  wire  _T_322; // @[FIFOVec.scala 49:90:@87882.4]
  wire  _T_323; // @[FIFOVec.scala 49:90:@87883.4]
  wire  _T_324; // @[FIFOVec.scala 49:90:@87884.4]
  wire  _T_325; // @[FIFOVec.scala 49:90:@87885.4]
  wire  _T_326; // @[FIFOVec.scala 49:90:@87886.4]
  wire  _T_327; // @[FIFOVec.scala 49:90:@87887.4]
  wire  _T_328; // @[FIFOVec.scala 49:90:@87888.4]
  wire  _T_329; // @[FIFOVec.scala 49:90:@87889.4]
  wire  _T_330; // @[FIFOVec.scala 49:90:@87890.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87860.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87861.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@87891.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87862.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@87891.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87863.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@87891.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87864.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@87891.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87865.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@87891.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87866.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@87891.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87867.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@87891.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87868.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@87891.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87869.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@87891.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87870.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@87891.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87871.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@87891.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87872.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@87891.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87873.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@87891.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87874.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@87891.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87875.4]
  wire  _GEN_15; // @[FIFOVec.scala 49:21:@87891.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@87910.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@87911.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@87912.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@87913.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@87914.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@87915.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@87916.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@87917.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@87918.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@87919.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@87920.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@87921.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@87922.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@87923.4]
  wire  _T_369; // @[FIFOVec.scala 51:93:@87924.4]
  wire  _T_335_0; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87894.4]
  wire  _T_335_1; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87895.4]
  wire  _GEN_17; // @[FIFOVec.scala 51:22:@87925.4]
  wire  _T_335_2; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87896.4]
  wire  _GEN_18; // @[FIFOVec.scala 51:22:@87925.4]
  wire  _T_335_3; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87897.4]
  wire  _GEN_19; // @[FIFOVec.scala 51:22:@87925.4]
  wire  _T_335_4; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87898.4]
  wire  _GEN_20; // @[FIFOVec.scala 51:22:@87925.4]
  wire  _T_335_5; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87899.4]
  wire  _GEN_21; // @[FIFOVec.scala 51:22:@87925.4]
  wire  _T_335_6; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87900.4]
  wire  _GEN_22; // @[FIFOVec.scala 51:22:@87925.4]
  wire  _T_335_7; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87901.4]
  wire  _GEN_23; // @[FIFOVec.scala 51:22:@87925.4]
  wire  _T_335_8; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87902.4]
  wire  _GEN_24; // @[FIFOVec.scala 51:22:@87925.4]
  wire  _T_335_9; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87903.4]
  wire  _GEN_25; // @[FIFOVec.scala 51:22:@87925.4]
  wire  _T_335_10; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87904.4]
  wire  _GEN_26; // @[FIFOVec.scala 51:22:@87925.4]
  wire  _T_335_11; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87905.4]
  wire  _GEN_27; // @[FIFOVec.scala 51:22:@87925.4]
  wire  _T_335_12; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87906.4]
  wire  _GEN_28; // @[FIFOVec.scala 51:22:@87925.4]
  wire  _T_335_13; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87907.4]
  wire  _GEN_29; // @[FIFOVec.scala 51:22:@87925.4]
  wire  _T_335_14; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87908.4]
  wire  _GEN_30; // @[FIFOVec.scala 51:22:@87925.4]
  wire  _T_335_15; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87909.4]
  wire  _GEN_31; // @[FIFOVec.scala 51:22:@87925.4]
  wire [31:0] _T_374_0; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87928.4]
  wire [31:0] _T_374_1; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87929.4]
  wire [31:0] _GEN_33; // @[FIFOVec.scala 53:42:@88200.4]
  wire [31:0] _T_374_2; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87930.4]
  wire [31:0] _GEN_34; // @[FIFOVec.scala 53:42:@88200.4]
  wire [31:0] _T_374_3; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87931.4]
  wire [31:0] _GEN_35; // @[FIFOVec.scala 53:42:@88200.4]
  wire [31:0] _T_374_4; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87932.4]
  wire [31:0] _GEN_36; // @[FIFOVec.scala 53:42:@88200.4]
  wire [31:0] _T_374_5; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87933.4]
  wire [31:0] _GEN_37; // @[FIFOVec.scala 53:42:@88200.4]
  wire [31:0] _T_374_6; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87934.4]
  wire [31:0] _GEN_38; // @[FIFOVec.scala 53:42:@88200.4]
  wire [31:0] _T_374_7; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87935.4]
  wire [31:0] _GEN_39; // @[FIFOVec.scala 53:42:@88200.4]
  wire [31:0] _T_374_8; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87936.4]
  wire [31:0] _GEN_40; // @[FIFOVec.scala 53:42:@88200.4]
  wire [31:0] _T_374_9; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87937.4]
  wire [31:0] _GEN_41; // @[FIFOVec.scala 53:42:@88200.4]
  wire [31:0] _T_374_10; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87938.4]
  wire [31:0] _GEN_42; // @[FIFOVec.scala 53:42:@88200.4]
  wire [31:0] _T_374_11; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87939.4]
  wire [31:0] _GEN_43; // @[FIFOVec.scala 53:42:@88200.4]
  wire [31:0] _T_374_12; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87940.4]
  wire [31:0] _GEN_44; // @[FIFOVec.scala 53:42:@88200.4]
  wire [31:0] _T_374_13; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87941.4]
  wire [31:0] _GEN_45; // @[FIFOVec.scala 53:42:@88200.4]
  wire [31:0] _T_374_14; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87942.4]
  wire [31:0] _GEN_46; // @[FIFOVec.scala 53:42:@88200.4]
  wire [31:0] _T_374_15; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87943.4]
  wire [31:0] _GEN_47; // @[FIFOVec.scala 53:42:@88200.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@87275.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@87286.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out)
  );
  FIFO_1 fifos_0 ( // @[FIFOVec.scala 40:19:@87299.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_1 fifos_1 ( // @[FIFOVec.scala 40:19:@87334.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_1 fifos_2 ( // @[FIFOVec.scala 40:19:@87369.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_1 fifos_3 ( // @[FIFOVec.scala 40:19:@87404.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_1 fifos_4 ( // @[FIFOVec.scala 40:19:@87439.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_1 fifos_5 ( // @[FIFOVec.scala 40:19:@87474.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_1 fifos_6 ( // @[FIFOVec.scala 40:19:@87509.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_1 fifos_7 ( // @[FIFOVec.scala 40:19:@87544.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_1 fifos_8 ( // @[FIFOVec.scala 40:19:@87579.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_1 fifos_9 ( // @[FIFOVec.scala 40:19:@87614.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_1 fifos_10 ( // @[FIFOVec.scala 40:19:@87649.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_1 fifos_11 ( // @[FIFOVec.scala 40:19:@87684.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_1 fifos_12 ( // @[FIFOVec.scala 40:19:@87719.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_1 fifos_13 ( // @[FIFOVec.scala 40:19:@87754.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_1 fifos_14 ( // @[FIFOVec.scala 40:19:@87789.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_1 fifos_15 ( // @[FIFOVec.scala 40:19:@87824.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign readEn = io_out_valid & io_out_ready; // @[FIFOVec.scala 20:29:@87273.4]
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@87274.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@87297.4]
  assign deqDecoder = 16'h1 << deqCounter_io_out; // @[OneHot.scala 45:35:@87298.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@87324.4]
  assign _T_151 = io_chainEnq ? _T_149 : 1'h1; // @[FIFOVec.scala 42:25:@87325.4]
  assign _T_154 = deqDecoder[0]; // @[FIFOVec.scala 44:50:@87330.4]
  assign _T_156 = io_chainDeq ? _T_154 : 1'h1; // @[FIFOVec.scala 44:26:@87331.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@87359.4]
  assign _T_160 = io_chainEnq ? _T_158 : 1'h1; // @[FIFOVec.scala 42:25:@87360.4]
  assign _T_163 = deqDecoder[1]; // @[FIFOVec.scala 44:50:@87365.4]
  assign _T_165 = io_chainDeq ? _T_163 : 1'h1; // @[FIFOVec.scala 44:26:@87366.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@87394.4]
  assign _T_169 = io_chainEnq ? _T_167 : 1'h1; // @[FIFOVec.scala 42:25:@87395.4]
  assign _T_172 = deqDecoder[2]; // @[FIFOVec.scala 44:50:@87400.4]
  assign _T_174 = io_chainDeq ? _T_172 : 1'h1; // @[FIFOVec.scala 44:26:@87401.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@87429.4]
  assign _T_178 = io_chainEnq ? _T_176 : 1'h1; // @[FIFOVec.scala 42:25:@87430.4]
  assign _T_181 = deqDecoder[3]; // @[FIFOVec.scala 44:50:@87435.4]
  assign _T_183 = io_chainDeq ? _T_181 : 1'h1; // @[FIFOVec.scala 44:26:@87436.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@87464.4]
  assign _T_187 = io_chainEnq ? _T_185 : 1'h1; // @[FIFOVec.scala 42:25:@87465.4]
  assign _T_190 = deqDecoder[4]; // @[FIFOVec.scala 44:50:@87470.4]
  assign _T_192 = io_chainDeq ? _T_190 : 1'h1; // @[FIFOVec.scala 44:26:@87471.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@87499.4]
  assign _T_196 = io_chainEnq ? _T_194 : 1'h1; // @[FIFOVec.scala 42:25:@87500.4]
  assign _T_199 = deqDecoder[5]; // @[FIFOVec.scala 44:50:@87505.4]
  assign _T_201 = io_chainDeq ? _T_199 : 1'h1; // @[FIFOVec.scala 44:26:@87506.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@87534.4]
  assign _T_205 = io_chainEnq ? _T_203 : 1'h1; // @[FIFOVec.scala 42:25:@87535.4]
  assign _T_208 = deqDecoder[6]; // @[FIFOVec.scala 44:50:@87540.4]
  assign _T_210 = io_chainDeq ? _T_208 : 1'h1; // @[FIFOVec.scala 44:26:@87541.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@87569.4]
  assign _T_214 = io_chainEnq ? _T_212 : 1'h1; // @[FIFOVec.scala 42:25:@87570.4]
  assign _T_217 = deqDecoder[7]; // @[FIFOVec.scala 44:50:@87575.4]
  assign _T_219 = io_chainDeq ? _T_217 : 1'h1; // @[FIFOVec.scala 44:26:@87576.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@87604.4]
  assign _T_223 = io_chainEnq ? _T_221 : 1'h1; // @[FIFOVec.scala 42:25:@87605.4]
  assign _T_226 = deqDecoder[8]; // @[FIFOVec.scala 44:50:@87610.4]
  assign _T_228 = io_chainDeq ? _T_226 : 1'h1; // @[FIFOVec.scala 44:26:@87611.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@87639.4]
  assign _T_232 = io_chainEnq ? _T_230 : 1'h1; // @[FIFOVec.scala 42:25:@87640.4]
  assign _T_235 = deqDecoder[9]; // @[FIFOVec.scala 44:50:@87645.4]
  assign _T_237 = io_chainDeq ? _T_235 : 1'h1; // @[FIFOVec.scala 44:26:@87646.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@87674.4]
  assign _T_241 = io_chainEnq ? _T_239 : 1'h1; // @[FIFOVec.scala 42:25:@87675.4]
  assign _T_244 = deqDecoder[10]; // @[FIFOVec.scala 44:50:@87680.4]
  assign _T_246 = io_chainDeq ? _T_244 : 1'h1; // @[FIFOVec.scala 44:26:@87681.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@87709.4]
  assign _T_250 = io_chainEnq ? _T_248 : 1'h1; // @[FIFOVec.scala 42:25:@87710.4]
  assign _T_253 = deqDecoder[11]; // @[FIFOVec.scala 44:50:@87715.4]
  assign _T_255 = io_chainDeq ? _T_253 : 1'h1; // @[FIFOVec.scala 44:26:@87716.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@87744.4]
  assign _T_259 = io_chainEnq ? _T_257 : 1'h1; // @[FIFOVec.scala 42:25:@87745.4]
  assign _T_262 = deqDecoder[12]; // @[FIFOVec.scala 44:50:@87750.4]
  assign _T_264 = io_chainDeq ? _T_262 : 1'h1; // @[FIFOVec.scala 44:26:@87751.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@87779.4]
  assign _T_268 = io_chainEnq ? _T_266 : 1'h1; // @[FIFOVec.scala 42:25:@87780.4]
  assign _T_271 = deqDecoder[13]; // @[FIFOVec.scala 44:50:@87785.4]
  assign _T_273 = io_chainDeq ? _T_271 : 1'h1; // @[FIFOVec.scala 44:26:@87786.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@87814.4]
  assign _T_277 = io_chainEnq ? _T_275 : 1'h1; // @[FIFOVec.scala 42:25:@87815.4]
  assign _T_280 = deqDecoder[14]; // @[FIFOVec.scala 44:50:@87820.4]
  assign _T_282 = io_chainDeq ? _T_280 : 1'h1; // @[FIFOVec.scala 44:26:@87821.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@87849.4]
  assign _T_286 = io_chainEnq ? _T_284 : 1'h1; // @[FIFOVec.scala 42:25:@87850.4]
  assign _T_289 = deqDecoder[15]; // @[FIFOVec.scala 44:50:@87855.4]
  assign _T_291 = io_chainDeq ? _T_289 : 1'h1; // @[FIFOVec.scala 44:26:@87856.4]
  assign _T_316 = fifos_0_io_in_ready & fifos_1_io_in_ready; // @[FIFOVec.scala 49:90:@87876.4]
  assign _T_317 = _T_316 & fifos_2_io_in_ready; // @[FIFOVec.scala 49:90:@87877.4]
  assign _T_318 = _T_317 & fifos_3_io_in_ready; // @[FIFOVec.scala 49:90:@87878.4]
  assign _T_319 = _T_318 & fifos_4_io_in_ready; // @[FIFOVec.scala 49:90:@87879.4]
  assign _T_320 = _T_319 & fifos_5_io_in_ready; // @[FIFOVec.scala 49:90:@87880.4]
  assign _T_321 = _T_320 & fifos_6_io_in_ready; // @[FIFOVec.scala 49:90:@87881.4]
  assign _T_322 = _T_321 & fifos_7_io_in_ready; // @[FIFOVec.scala 49:90:@87882.4]
  assign _T_323 = _T_322 & fifos_8_io_in_ready; // @[FIFOVec.scala 49:90:@87883.4]
  assign _T_324 = _T_323 & fifos_9_io_in_ready; // @[FIFOVec.scala 49:90:@87884.4]
  assign _T_325 = _T_324 & fifos_10_io_in_ready; // @[FIFOVec.scala 49:90:@87885.4]
  assign _T_326 = _T_325 & fifos_11_io_in_ready; // @[FIFOVec.scala 49:90:@87886.4]
  assign _T_327 = _T_326 & fifos_12_io_in_ready; // @[FIFOVec.scala 49:90:@87887.4]
  assign _T_328 = _T_327 & fifos_13_io_in_ready; // @[FIFOVec.scala 49:90:@87888.4]
  assign _T_329 = _T_328 & fifos_14_io_in_ready; // @[FIFOVec.scala 49:90:@87889.4]
  assign _T_330 = _T_329 & fifos_15_io_in_ready; // @[FIFOVec.scala 49:90:@87890.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87860.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87861.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@87891.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87862.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@87891.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87863.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@87891.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87864.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@87891.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87865.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@87891.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87866.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@87891.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87867.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@87891.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87868.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@87891.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87869.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@87891.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87870.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@87891.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87871.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@87891.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87872.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@87891.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87873.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@87891.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87874.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@87891.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@87859.4 FIFOVec.scala 49:42:@87875.4]
  assign _GEN_15 = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:21:@87891.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@87910.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@87911.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@87912.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@87913.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@87914.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@87915.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@87916.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@87917.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@87918.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@87919.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@87920.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@87921.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@87922.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@87923.4]
  assign _T_369 = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:93:@87924.4]
  assign _T_335_0 = fifos_0_io_out_valid; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87894.4]
  assign _T_335_1 = fifos_1_io_out_valid; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87895.4]
  assign _GEN_17 = 4'h1 == deqCounter_io_out ? _T_335_1 : _T_335_0; // @[FIFOVec.scala 51:22:@87925.4]
  assign _T_335_2 = fifos_2_io_out_valid; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87896.4]
  assign _GEN_18 = 4'h2 == deqCounter_io_out ? _T_335_2 : _GEN_17; // @[FIFOVec.scala 51:22:@87925.4]
  assign _T_335_3 = fifos_3_io_out_valid; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87897.4]
  assign _GEN_19 = 4'h3 == deqCounter_io_out ? _T_335_3 : _GEN_18; // @[FIFOVec.scala 51:22:@87925.4]
  assign _T_335_4 = fifos_4_io_out_valid; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87898.4]
  assign _GEN_20 = 4'h4 == deqCounter_io_out ? _T_335_4 : _GEN_19; // @[FIFOVec.scala 51:22:@87925.4]
  assign _T_335_5 = fifos_5_io_out_valid; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87899.4]
  assign _GEN_21 = 4'h5 == deqCounter_io_out ? _T_335_5 : _GEN_20; // @[FIFOVec.scala 51:22:@87925.4]
  assign _T_335_6 = fifos_6_io_out_valid; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87900.4]
  assign _GEN_22 = 4'h6 == deqCounter_io_out ? _T_335_6 : _GEN_21; // @[FIFOVec.scala 51:22:@87925.4]
  assign _T_335_7 = fifos_7_io_out_valid; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87901.4]
  assign _GEN_23 = 4'h7 == deqCounter_io_out ? _T_335_7 : _GEN_22; // @[FIFOVec.scala 51:22:@87925.4]
  assign _T_335_8 = fifos_8_io_out_valid; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87902.4]
  assign _GEN_24 = 4'h8 == deqCounter_io_out ? _T_335_8 : _GEN_23; // @[FIFOVec.scala 51:22:@87925.4]
  assign _T_335_9 = fifos_9_io_out_valid; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87903.4]
  assign _GEN_25 = 4'h9 == deqCounter_io_out ? _T_335_9 : _GEN_24; // @[FIFOVec.scala 51:22:@87925.4]
  assign _T_335_10 = fifos_10_io_out_valid; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87904.4]
  assign _GEN_26 = 4'ha == deqCounter_io_out ? _T_335_10 : _GEN_25; // @[FIFOVec.scala 51:22:@87925.4]
  assign _T_335_11 = fifos_11_io_out_valid; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87905.4]
  assign _GEN_27 = 4'hb == deqCounter_io_out ? _T_335_11 : _GEN_26; // @[FIFOVec.scala 51:22:@87925.4]
  assign _T_335_12 = fifos_12_io_out_valid; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87906.4]
  assign _GEN_28 = 4'hc == deqCounter_io_out ? _T_335_12 : _GEN_27; // @[FIFOVec.scala 51:22:@87925.4]
  assign _T_335_13 = fifos_13_io_out_valid; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87907.4]
  assign _GEN_29 = 4'hd == deqCounter_io_out ? _T_335_13 : _GEN_28; // @[FIFOVec.scala 51:22:@87925.4]
  assign _T_335_14 = fifos_14_io_out_valid; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87908.4]
  assign _GEN_30 = 4'he == deqCounter_io_out ? _T_335_14 : _GEN_29; // @[FIFOVec.scala 51:22:@87925.4]
  assign _T_335_15 = fifos_15_io_out_valid; // @[FIFOVec.scala 51:43:@87893.4 FIFOVec.scala 51:43:@87909.4]
  assign _GEN_31 = 4'hf == deqCounter_io_out ? _T_335_15 : _GEN_30; // @[FIFOVec.scala 51:22:@87925.4]
  assign _T_374_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87928.4]
  assign _T_374_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87929.4]
  assign _GEN_33 = 4'h1 == deqCounter_io_out ? _T_374_1 : _T_374_0; // @[FIFOVec.scala 53:42:@88200.4]
  assign _T_374_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87930.4]
  assign _GEN_34 = 4'h2 == deqCounter_io_out ? _T_374_2 : _GEN_33; // @[FIFOVec.scala 53:42:@88200.4]
  assign _T_374_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87931.4]
  assign _GEN_35 = 4'h3 == deqCounter_io_out ? _T_374_3 : _GEN_34; // @[FIFOVec.scala 53:42:@88200.4]
  assign _T_374_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87932.4]
  assign _GEN_36 = 4'h4 == deqCounter_io_out ? _T_374_4 : _GEN_35; // @[FIFOVec.scala 53:42:@88200.4]
  assign _T_374_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87933.4]
  assign _GEN_37 = 4'h5 == deqCounter_io_out ? _T_374_5 : _GEN_36; // @[FIFOVec.scala 53:42:@88200.4]
  assign _T_374_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87934.4]
  assign _GEN_38 = 4'h6 == deqCounter_io_out ? _T_374_6 : _GEN_37; // @[FIFOVec.scala 53:42:@88200.4]
  assign _T_374_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87935.4]
  assign _GEN_39 = 4'h7 == deqCounter_io_out ? _T_374_7 : _GEN_38; // @[FIFOVec.scala 53:42:@88200.4]
  assign _T_374_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87936.4]
  assign _GEN_40 = 4'h8 == deqCounter_io_out ? _T_374_8 : _GEN_39; // @[FIFOVec.scala 53:42:@88200.4]
  assign _T_374_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87937.4]
  assign _GEN_41 = 4'h9 == deqCounter_io_out ? _T_374_9 : _GEN_40; // @[FIFOVec.scala 53:42:@88200.4]
  assign _T_374_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87938.4]
  assign _GEN_42 = 4'ha == deqCounter_io_out ? _T_374_10 : _GEN_41; // @[FIFOVec.scala 53:42:@88200.4]
  assign _T_374_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87939.4]
  assign _GEN_43 = 4'hb == deqCounter_io_out ? _T_374_11 : _GEN_42; // @[FIFOVec.scala 53:42:@88200.4]
  assign _T_374_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87940.4]
  assign _GEN_44 = 4'hc == deqCounter_io_out ? _T_374_12 : _GEN_43; // @[FIFOVec.scala 53:42:@88200.4]
  assign _T_374_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87941.4]
  assign _GEN_45 = 4'hd == deqCounter_io_out ? _T_374_13 : _GEN_44; // @[FIFOVec.scala 53:42:@88200.4]
  assign _T_374_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87942.4]
  assign _GEN_46 = 4'he == deqCounter_io_out ? _T_374_14 : _GEN_45; // @[FIFOVec.scala 53:42:@88200.4]
  assign _T_374_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:65:@87927.4 FIFOVec.scala 53:65:@87943.4]
  assign _GEN_47 = 4'hf == deqCounter_io_out ? _T_374_15 : _GEN_46; // @[FIFOVec.scala 53:42:@88200.4]
  assign io_in_ready = io_chainEnq ? _GEN_15 : _T_330; // @[FIFOVec.scala 49:15:@87892.4]
  assign io_out_valid = io_chainDeq ? _GEN_31 : _T_369; // @[FIFOVec.scala 51:16:@87926.4]
  assign io_out_bits_0 = io_chainDeq ? _GEN_47 : _T_374_0; // @[FIFOVec.scala 53:15:@88234.4]
  assign io_out_bits_1 = io_chainDeq ? _GEN_47 : _T_374_1; // @[FIFOVec.scala 53:15:@88235.4]
  assign io_out_bits_2 = io_chainDeq ? _GEN_47 : _T_374_2; // @[FIFOVec.scala 53:15:@88236.4]
  assign io_out_bits_3 = io_chainDeq ? _GEN_47 : _T_374_3; // @[FIFOVec.scala 53:15:@88237.4]
  assign io_out_bits_4 = io_chainDeq ? _GEN_47 : _T_374_4; // @[FIFOVec.scala 53:15:@88238.4]
  assign io_out_bits_5 = io_chainDeq ? _GEN_47 : _T_374_5; // @[FIFOVec.scala 53:15:@88239.4]
  assign io_out_bits_6 = io_chainDeq ? _GEN_47 : _T_374_6; // @[FIFOVec.scala 53:15:@88240.4]
  assign io_out_bits_7 = io_chainDeq ? _GEN_47 : _T_374_7; // @[FIFOVec.scala 53:15:@88241.4]
  assign io_out_bits_8 = io_chainDeq ? _GEN_47 : _T_374_8; // @[FIFOVec.scala 53:15:@88242.4]
  assign io_out_bits_9 = io_chainDeq ? _GEN_47 : _T_374_9; // @[FIFOVec.scala 53:15:@88243.4]
  assign io_out_bits_10 = io_chainDeq ? _GEN_47 : _T_374_10; // @[FIFOVec.scala 53:15:@88244.4]
  assign io_out_bits_11 = io_chainDeq ? _GEN_47 : _T_374_11; // @[FIFOVec.scala 53:15:@88245.4]
  assign io_out_bits_12 = io_chainDeq ? _GEN_47 : _T_374_12; // @[FIFOVec.scala 53:15:@88246.4]
  assign io_out_bits_13 = io_chainDeq ? _GEN_47 : _T_374_13; // @[FIFOVec.scala 53:15:@88247.4]
  assign io_out_bits_14 = io_chainDeq ? _GEN_47 : _T_374_14; // @[FIFOVec.scala 53:15:@88248.4]
  assign io_out_bits_15 = io_chainDeq ? _GEN_47 : _T_374_15; // @[FIFOVec.scala 53:15:@88249.4]
  assign enqCounter_clock = clock; // @[:@87276.4]
  assign enqCounter_reset = reset; // @[:@87277.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = writeEn & io_chainEnq; // @[FIFOVec.scala 26:24:@87284.4]
  assign enqCounter_io_stride = 4'h1; // @[FIFOVec.scala 27:24:@87285.4]
  assign deqCounter_clock = clock; // @[:@87287.4]
  assign deqCounter_reset = reset; // @[:@87288.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = readEn & io_chainDeq; // @[FIFOVec.scala 30:24:@87295.4]
  assign deqCounter_io_stride = 4'h1; // @[FIFOVec.scala 31:24:@87296.4]
  assign fifos_0_clock = clock; // @[:@87300.4]
  assign fifos_0_reset = reset; // @[:@87301.4]
  assign fifos_0_io_in_valid = _T_151 & writeEn; // @[FIFOVec.scala 42:19:@87327.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@87329.4]
  assign fifos_0_io_out_ready = _T_156 & readEn; // @[FIFOVec.scala 44:20:@87333.4]
  assign fifos_1_clock = clock; // @[:@87335.4]
  assign fifos_1_reset = reset; // @[:@87336.4]
  assign fifos_1_io_in_valid = _T_160 & writeEn; // @[FIFOVec.scala 42:19:@87362.4]
  assign fifos_1_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_1; // @[FIFOVec.scala 43:18:@87364.4]
  assign fifos_1_io_out_ready = _T_165 & readEn; // @[FIFOVec.scala 44:20:@87368.4]
  assign fifos_2_clock = clock; // @[:@87370.4]
  assign fifos_2_reset = reset; // @[:@87371.4]
  assign fifos_2_io_in_valid = _T_169 & writeEn; // @[FIFOVec.scala 42:19:@87397.4]
  assign fifos_2_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_2; // @[FIFOVec.scala 43:18:@87399.4]
  assign fifos_2_io_out_ready = _T_174 & readEn; // @[FIFOVec.scala 44:20:@87403.4]
  assign fifos_3_clock = clock; // @[:@87405.4]
  assign fifos_3_reset = reset; // @[:@87406.4]
  assign fifos_3_io_in_valid = _T_178 & writeEn; // @[FIFOVec.scala 42:19:@87432.4]
  assign fifos_3_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_3; // @[FIFOVec.scala 43:18:@87434.4]
  assign fifos_3_io_out_ready = _T_183 & readEn; // @[FIFOVec.scala 44:20:@87438.4]
  assign fifos_4_clock = clock; // @[:@87440.4]
  assign fifos_4_reset = reset; // @[:@87441.4]
  assign fifos_4_io_in_valid = _T_187 & writeEn; // @[FIFOVec.scala 42:19:@87467.4]
  assign fifos_4_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_4; // @[FIFOVec.scala 43:18:@87469.4]
  assign fifos_4_io_out_ready = _T_192 & readEn; // @[FIFOVec.scala 44:20:@87473.4]
  assign fifos_5_clock = clock; // @[:@87475.4]
  assign fifos_5_reset = reset; // @[:@87476.4]
  assign fifos_5_io_in_valid = _T_196 & writeEn; // @[FIFOVec.scala 42:19:@87502.4]
  assign fifos_5_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_5; // @[FIFOVec.scala 43:18:@87504.4]
  assign fifos_5_io_out_ready = _T_201 & readEn; // @[FIFOVec.scala 44:20:@87508.4]
  assign fifos_6_clock = clock; // @[:@87510.4]
  assign fifos_6_reset = reset; // @[:@87511.4]
  assign fifos_6_io_in_valid = _T_205 & writeEn; // @[FIFOVec.scala 42:19:@87537.4]
  assign fifos_6_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_6; // @[FIFOVec.scala 43:18:@87539.4]
  assign fifos_6_io_out_ready = _T_210 & readEn; // @[FIFOVec.scala 44:20:@87543.4]
  assign fifos_7_clock = clock; // @[:@87545.4]
  assign fifos_7_reset = reset; // @[:@87546.4]
  assign fifos_7_io_in_valid = _T_214 & writeEn; // @[FIFOVec.scala 42:19:@87572.4]
  assign fifos_7_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_7; // @[FIFOVec.scala 43:18:@87574.4]
  assign fifos_7_io_out_ready = _T_219 & readEn; // @[FIFOVec.scala 44:20:@87578.4]
  assign fifos_8_clock = clock; // @[:@87580.4]
  assign fifos_8_reset = reset; // @[:@87581.4]
  assign fifos_8_io_in_valid = _T_223 & writeEn; // @[FIFOVec.scala 42:19:@87607.4]
  assign fifos_8_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_8; // @[FIFOVec.scala 43:18:@87609.4]
  assign fifos_8_io_out_ready = _T_228 & readEn; // @[FIFOVec.scala 44:20:@87613.4]
  assign fifos_9_clock = clock; // @[:@87615.4]
  assign fifos_9_reset = reset; // @[:@87616.4]
  assign fifos_9_io_in_valid = _T_232 & writeEn; // @[FIFOVec.scala 42:19:@87642.4]
  assign fifos_9_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_9; // @[FIFOVec.scala 43:18:@87644.4]
  assign fifos_9_io_out_ready = _T_237 & readEn; // @[FIFOVec.scala 44:20:@87648.4]
  assign fifos_10_clock = clock; // @[:@87650.4]
  assign fifos_10_reset = reset; // @[:@87651.4]
  assign fifos_10_io_in_valid = _T_241 & writeEn; // @[FIFOVec.scala 42:19:@87677.4]
  assign fifos_10_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_10; // @[FIFOVec.scala 43:18:@87679.4]
  assign fifos_10_io_out_ready = _T_246 & readEn; // @[FIFOVec.scala 44:20:@87683.4]
  assign fifos_11_clock = clock; // @[:@87685.4]
  assign fifos_11_reset = reset; // @[:@87686.4]
  assign fifos_11_io_in_valid = _T_250 & writeEn; // @[FIFOVec.scala 42:19:@87712.4]
  assign fifos_11_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_11; // @[FIFOVec.scala 43:18:@87714.4]
  assign fifos_11_io_out_ready = _T_255 & readEn; // @[FIFOVec.scala 44:20:@87718.4]
  assign fifos_12_clock = clock; // @[:@87720.4]
  assign fifos_12_reset = reset; // @[:@87721.4]
  assign fifos_12_io_in_valid = _T_259 & writeEn; // @[FIFOVec.scala 42:19:@87747.4]
  assign fifos_12_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_12; // @[FIFOVec.scala 43:18:@87749.4]
  assign fifos_12_io_out_ready = _T_264 & readEn; // @[FIFOVec.scala 44:20:@87753.4]
  assign fifos_13_clock = clock; // @[:@87755.4]
  assign fifos_13_reset = reset; // @[:@87756.4]
  assign fifos_13_io_in_valid = _T_268 & writeEn; // @[FIFOVec.scala 42:19:@87782.4]
  assign fifos_13_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_13; // @[FIFOVec.scala 43:18:@87784.4]
  assign fifos_13_io_out_ready = _T_273 & readEn; // @[FIFOVec.scala 44:20:@87788.4]
  assign fifos_14_clock = clock; // @[:@87790.4]
  assign fifos_14_reset = reset; // @[:@87791.4]
  assign fifos_14_io_in_valid = _T_277 & writeEn; // @[FIFOVec.scala 42:19:@87817.4]
  assign fifos_14_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_14; // @[FIFOVec.scala 43:18:@87819.4]
  assign fifos_14_io_out_ready = _T_282 & readEn; // @[FIFOVec.scala 44:20:@87823.4]
  assign fifos_15_clock = clock; // @[:@87825.4]
  assign fifos_15_reset = reset; // @[:@87826.4]
  assign fifos_15_io_in_valid = _T_286 & writeEn; // @[FIFOVec.scala 42:19:@87852.4]
  assign fifos_15_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_15; // @[FIFOVec.scala 43:18:@87854.4]
  assign fifos_15_io_out_ready = _T_291 & readEn; // @[FIFOVec.scala 44:20:@87858.4]
endmodule
module SRAM_93( // @[:@88339.2]
  input        clock, // @[:@88340.4]
  input  [5:0] io_raddr, // @[:@88342.4]
  input        io_wen, // @[:@88342.4]
  input  [5:0] io_waddr // @[:@88342.4]
);
  wire [63:0] SRAMVerilogSim_rdata; // @[SRAM.scala 187:23:@88344.4]
  wire [63:0] SRAMVerilogSim_wdata; // @[SRAM.scala 187:23:@88344.4]
  wire  SRAMVerilogSim_backpressure; // @[SRAM.scala 187:23:@88344.4]
  wire  SRAMVerilogSim_wen; // @[SRAM.scala 187:23:@88344.4]
  wire  SRAMVerilogSim_waddrEn; // @[SRAM.scala 187:23:@88344.4]
  wire  SRAMVerilogSim_raddrEn; // @[SRAM.scala 187:23:@88344.4]
  wire [5:0] SRAMVerilogSim_waddr; // @[SRAM.scala 187:23:@88344.4]
  wire [5:0] SRAMVerilogSim_raddr; // @[SRAM.scala 187:23:@88344.4]
  wire  SRAMVerilogSim_clk; // @[SRAM.scala 187:23:@88344.4]
  SRAMVerilogSim #(.DWIDTH(64), .WORDS(64), .AWIDTH(6)) SRAMVerilogSim ( // @[SRAM.scala 187:23:@88344.4]
    .rdata(SRAMVerilogSim_rdata),
    .wdata(SRAMVerilogSim_wdata),
    .backpressure(SRAMVerilogSim_backpressure),
    .wen(SRAMVerilogSim_wen),
    .waddrEn(SRAMVerilogSim_waddrEn),
    .raddrEn(SRAMVerilogSim_raddrEn),
    .waddr(SRAMVerilogSim_waddr),
    .raddr(SRAMVerilogSim_raddr),
    .clk(SRAMVerilogSim_clk)
  );
  assign SRAMVerilogSim_wdata = 64'h0; // @[SRAM.scala 192:20:@88358.4]
  assign SRAMVerilogSim_backpressure = 1'h1; // @[SRAM.scala 193:27:@88359.4]
  assign SRAMVerilogSim_wen = io_wen; // @[SRAM.scala 190:18:@88356.4]
  assign SRAMVerilogSim_waddrEn = 1'h1; // @[SRAM.scala 195:22:@88361.4]
  assign SRAMVerilogSim_raddrEn = 1'h1; // @[SRAM.scala 194:22:@88360.4]
  assign SRAMVerilogSim_waddr = io_waddr; // @[SRAM.scala 191:20:@88357.4]
  assign SRAMVerilogSim_raddr = io_raddr; // @[SRAM.scala 189:20:@88355.4]
  assign SRAMVerilogSim_clk = clock; // @[SRAM.scala 188:18:@88354.4]
endmodule
module FIFO_17( // @[:@88366.2]
  input   clock, // @[:@88367.4]
  input   reset, // @[:@88368.4]
  output  io_in_ready, // @[:@88369.4]
  input   io_in_valid // @[:@88369.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@88635.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@88635.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@88635.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@88635.4]
  wire [5:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@88635.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@88635.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@88635.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@88645.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@88645.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@88645.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@88645.4]
  wire [5:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@88645.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@88645.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@88645.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@88660.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@88660.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@88660.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@88660.4]
  wire  writeEn; // @[FIFO.scala 30:29:@88633.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@88655.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@88656.4]
  wire  full; // @[FIFO.scala 46:23:@88659.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@88671.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@88635.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@88645.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_93 SRAM ( // @[FIFO.scala 73:19:@88660.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@88633.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@88656.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@88659.4]
  assign _GEN_0 = writeEn ? writeEn : maybeFull; // @[FIFO.scala 83:29:@88671.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@88677.4]
  assign enqCounter_clock = clock; // @[:@88636.4]
  assign enqCounter_reset = reset; // @[:@88637.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@88643.4]
  assign enqCounter_io_stride = 6'h1; // @[FIFO.scala 37:24:@88644.4]
  assign deqCounter_clock = clock; // @[:@88646.4]
  assign deqCounter_reset = reset; // @[:@88647.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = 1'h0; // @[FIFO.scala 40:24:@88653.4]
  assign deqCounter_io_stride = 6'h1; // @[FIFO.scala 41:24:@88654.4]
  assign SRAM_clock = clock; // @[:@88661.4]
  assign SRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 75:16:@88664.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@88665.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@88666.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (writeEn) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_1( // @[:@88679.2]
  input   clock, // @[:@88680.4]
  input   reset, // @[:@88681.4]
  output  io_in_ready, // @[:@88682.4]
  input   io_in_valid // @[:@88682.4]
);
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@88710.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@88710.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@88710.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@88710.4]
  FIFO_17 fifos_0 ( // @[FIFOVec.scala 40:19:@88710.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid)
  );
  assign io_in_ready = fifos_0_io_in_ready; // @[FIFOVec.scala 49:15:@88988.4]
  assign fifos_0_clock = clock; // @[:@88711.4]
  assign fifos_0_reset = reset; // @[:@88712.4]
  assign fifos_0_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@88978.4]
endmodule
module FIFOWidthConvert( // @[:@89002.2]
  input         clock, // @[:@89003.4]
  input         reset, // @[:@89004.4]
  output        io_in_ready, // @[:@89005.4]
  input         io_in_valid, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_0, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_1, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_2, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_3, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_4, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_5, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_6, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_7, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_8, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_9, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_10, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_11, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_12, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_13, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_14, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_15, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_16, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_17, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_18, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_19, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_20, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_21, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_22, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_23, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_24, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_25, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_26, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_27, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_28, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_29, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_30, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_31, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_32, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_33, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_34, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_35, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_36, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_37, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_38, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_39, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_40, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_41, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_42, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_43, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_44, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_45, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_46, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_47, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_48, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_49, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_50, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_51, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_52, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_53, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_54, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_55, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_56, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_57, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_58, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_59, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_60, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_61, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_62, // @[:@89005.4]
  input  [7:0]  io_in_bits_data_63, // @[:@89005.4]
  input         io_out_ready, // @[:@89005.4]
  output        io_out_valid, // @[:@89005.4]
  output [31:0] io_out_bits_data_0 // @[:@89005.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_in_bits_1; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_in_bits_2; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_in_bits_3; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_in_bits_4; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_in_bits_5; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_in_bits_6; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_in_bits_7; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_in_bits_8; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_in_bits_9; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_in_bits_10; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_in_bits_11; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_in_bits_12; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_in_bits_13; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_in_bits_14; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_in_bits_15; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_out_bits_1; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_out_bits_2; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_out_bits_3; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_out_bits_4; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_out_bits_5; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_out_bits_6; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_out_bits_7; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_out_bits_8; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_out_bits_9; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_out_bits_10; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_out_bits_11; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_out_bits_12; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_out_bits_13; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_out_bits_14; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire [31:0] FIFOVec_io_out_bits_15; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire  FIFOVec_io_chainEnq; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire  FIFOVec_io_chainDeq; // @[FIFOWidthConvert.scala 82:22:@89007.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 83:26:@89048.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 83:26:@89048.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 83:26:@89048.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 83:26:@89048.4]
  wire [79:0] _T_55; // @[Cat.scala 30:58:@89073.4]
  wire [151:0] _T_64; // @[Cat.scala 30:58:@89082.4]
  wire [223:0] _T_73; // @[Cat.scala 30:58:@89091.4]
  wire [295:0] _T_82; // @[Cat.scala 30:58:@89100.4]
  wire [367:0] _T_91; // @[Cat.scala 30:58:@89109.4]
  wire [439:0] _T_100; // @[Cat.scala 30:58:@89118.4]
  wire [511:0] _T_109; // @[Cat.scala 30:58:@89127.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 82:22:@89007.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_in_bits_1(FIFOVec_io_in_bits_1),
    .io_in_bits_2(FIFOVec_io_in_bits_2),
    .io_in_bits_3(FIFOVec_io_in_bits_3),
    .io_in_bits_4(FIFOVec_io_in_bits_4),
    .io_in_bits_5(FIFOVec_io_in_bits_5),
    .io_in_bits_6(FIFOVec_io_in_bits_6),
    .io_in_bits_7(FIFOVec_io_in_bits_7),
    .io_in_bits_8(FIFOVec_io_in_bits_8),
    .io_in_bits_9(FIFOVec_io_in_bits_9),
    .io_in_bits_10(FIFOVec_io_in_bits_10),
    .io_in_bits_11(FIFOVec_io_in_bits_11),
    .io_in_bits_12(FIFOVec_io_in_bits_12),
    .io_in_bits_13(FIFOVec_io_in_bits_13),
    .io_in_bits_14(FIFOVec_io_in_bits_14),
    .io_in_bits_15(FIFOVec_io_in_bits_15),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0),
    .io_out_bits_1(FIFOVec_io_out_bits_1),
    .io_out_bits_2(FIFOVec_io_out_bits_2),
    .io_out_bits_3(FIFOVec_io_out_bits_3),
    .io_out_bits_4(FIFOVec_io_out_bits_4),
    .io_out_bits_5(FIFOVec_io_out_bits_5),
    .io_out_bits_6(FIFOVec_io_out_bits_6),
    .io_out_bits_7(FIFOVec_io_out_bits_7),
    .io_out_bits_8(FIFOVec_io_out_bits_8),
    .io_out_bits_9(FIFOVec_io_out_bits_9),
    .io_out_bits_10(FIFOVec_io_out_bits_10),
    .io_out_bits_11(FIFOVec_io_out_bits_11),
    .io_out_bits_12(FIFOVec_io_out_bits_12),
    .io_out_bits_13(FIFOVec_io_out_bits_13),
    .io_out_bits_14(FIFOVec_io_out_bits_14),
    .io_out_bits_15(FIFOVec_io_out_bits_15),
    .io_chainEnq(FIFOVec_io_chainEnq),
    .io_chainDeq(FIFOVec_io_chainDeq)
  );
  FIFOVec_1 FIFOVec_1 ( // @[FIFOWidthConvert.scala 83:26:@89048.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid)
  );
  assign _T_55 = {io_in_bits_data_63,io_in_bits_data_62,io_in_bits_data_61,io_in_bits_data_60,io_in_bits_data_59,io_in_bits_data_58,io_in_bits_data_57,io_in_bits_data_56,io_in_bits_data_55,io_in_bits_data_54}; // @[Cat.scala 30:58:@89073.4]
  assign _T_64 = {_T_55,io_in_bits_data_53,io_in_bits_data_52,io_in_bits_data_51,io_in_bits_data_50,io_in_bits_data_49,io_in_bits_data_48,io_in_bits_data_47,io_in_bits_data_46,io_in_bits_data_45}; // @[Cat.scala 30:58:@89082.4]
  assign _T_73 = {_T_64,io_in_bits_data_44,io_in_bits_data_43,io_in_bits_data_42,io_in_bits_data_41,io_in_bits_data_40,io_in_bits_data_39,io_in_bits_data_38,io_in_bits_data_37,io_in_bits_data_36}; // @[Cat.scala 30:58:@89091.4]
  assign _T_82 = {_T_73,io_in_bits_data_35,io_in_bits_data_34,io_in_bits_data_33,io_in_bits_data_32,io_in_bits_data_31,io_in_bits_data_30,io_in_bits_data_29,io_in_bits_data_28,io_in_bits_data_27}; // @[Cat.scala 30:58:@89100.4]
  assign _T_91 = {_T_82,io_in_bits_data_26,io_in_bits_data_25,io_in_bits_data_24,io_in_bits_data_23,io_in_bits_data_22,io_in_bits_data_21,io_in_bits_data_20,io_in_bits_data_19,io_in_bits_data_18}; // @[Cat.scala 30:58:@89109.4]
  assign _T_100 = {_T_91,io_in_bits_data_17,io_in_bits_data_16,io_in_bits_data_15,io_in_bits_data_14,io_in_bits_data_13,io_in_bits_data_12,io_in_bits_data_11,io_in_bits_data_10,io_in_bits_data_9}; // @[Cat.scala 30:58:@89118.4]
  assign _T_109 = {_T_100,io_in_bits_data_8,io_in_bits_data_7,io_in_bits_data_6,io_in_bits_data_5,io_in_bits_data_4,io_in_bits_data_3,io_in_bits_data_2,io_in_bits_data_1,io_in_bits_data_0}; // @[Cat.scala 30:58:@89127.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 88:17:@89063.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 89:18:@89064.4]
  assign io_out_bits_data_0 = FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 96:22:@89185.4]
  assign FIFOVec_clock = clock; // @[:@89008.4]
  assign FIFOVec_reset = reset; // @[:@89009.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 92:22:@89177.4]
  assign FIFOVec_io_in_bits_0 = _T_109[31:0]; // @[FIFOWidthConvert.scala 91:21:@89161.4]
  assign FIFOVec_io_in_bits_1 = _T_109[63:32]; // @[FIFOWidthConvert.scala 91:21:@89162.4]
  assign FIFOVec_io_in_bits_2 = _T_109[95:64]; // @[FIFOWidthConvert.scala 91:21:@89163.4]
  assign FIFOVec_io_in_bits_3 = _T_109[127:96]; // @[FIFOWidthConvert.scala 91:21:@89164.4]
  assign FIFOVec_io_in_bits_4 = _T_109[159:128]; // @[FIFOWidthConvert.scala 91:21:@89165.4]
  assign FIFOVec_io_in_bits_5 = _T_109[191:160]; // @[FIFOWidthConvert.scala 91:21:@89166.4]
  assign FIFOVec_io_in_bits_6 = _T_109[223:192]; // @[FIFOWidthConvert.scala 91:21:@89167.4]
  assign FIFOVec_io_in_bits_7 = _T_109[255:224]; // @[FIFOWidthConvert.scala 91:21:@89168.4]
  assign FIFOVec_io_in_bits_8 = _T_109[287:256]; // @[FIFOWidthConvert.scala 91:21:@89169.4]
  assign FIFOVec_io_in_bits_9 = _T_109[319:288]; // @[FIFOWidthConvert.scala 91:21:@89170.4]
  assign FIFOVec_io_in_bits_10 = _T_109[351:320]; // @[FIFOWidthConvert.scala 91:21:@89171.4]
  assign FIFOVec_io_in_bits_11 = _T_109[383:352]; // @[FIFOWidthConvert.scala 91:21:@89172.4]
  assign FIFOVec_io_in_bits_12 = _T_109[415:384]; // @[FIFOWidthConvert.scala 91:21:@89173.4]
  assign FIFOVec_io_in_bits_13 = _T_109[447:416]; // @[FIFOWidthConvert.scala 91:21:@89174.4]
  assign FIFOVec_io_in_bits_14 = _T_109[479:448]; // @[FIFOWidthConvert.scala 91:21:@89175.4]
  assign FIFOVec_io_in_bits_15 = _T_109[511:480]; // @[FIFOWidthConvert.scala 91:21:@89176.4]
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 98:23:@89199.4]
  assign FIFOVec_io_chainEnq = 1'h0; // @[FIFOWidthConvert.scala 84:22:@89059.4]
  assign FIFOVec_io_chainDeq = 1'h1; // @[FIFOWidthConvert.scala 85:22:@89060.4]
  assign FIFOVec_1_clock = clock; // @[:@89049.4]
  assign FIFOVec_1_reset = reset; // @[:@89050.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 94:26:@89179.4]
endmodule
module StreamControllerLoad( // @[:@89201.2]
  input         clock, // @[:@89202.4]
  input         reset, // @[:@89203.4]
  input         io_dram_cmd_ready, // @[:@89204.4]
  output        io_dram_cmd_valid, // @[:@89204.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@89204.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@89204.4]
  output        io_dram_rresp_ready, // @[:@89204.4]
  input         io_dram_rresp_valid, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_0, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_1, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_2, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_3, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_4, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_5, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_6, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_7, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_8, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_9, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_10, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_11, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_12, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_13, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_14, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_15, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_16, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_17, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_18, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_19, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_20, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_21, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_22, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_23, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_24, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_25, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_26, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_27, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_28, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_29, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_30, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_31, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_32, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_33, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_34, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_35, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_36, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_37, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_38, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_39, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_40, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_41, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_42, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_43, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_44, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_45, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_46, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_47, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_48, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_49, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_50, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_51, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_52, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_53, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_54, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_55, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_56, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_57, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_58, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_59, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_60, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_61, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_62, // @[:@89204.4]
  input  [7:0]  io_dram_rresp_bits_rdata_63, // @[:@89204.4]
  output        io_load_cmd_ready, // @[:@89204.4]
  input         io_load_cmd_valid, // @[:@89204.4]
  input  [63:0] io_load_cmd_bits_addr, // @[:@89204.4]
  input  [31:0] io_load_cmd_bits_size, // @[:@89204.4]
  input         io_load_data_ready, // @[:@89204.4]
  output        io_load_data_valid, // @[:@89204.4]
  output [31:0] io_load_data_bits_rdata_0 // @[:@89204.4]
);
  wire  cmd_clock; // @[StreamController.scala 38:19:@89421.4]
  wire  cmd_reset; // @[StreamController.scala 38:19:@89421.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 38:19:@89421.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 38:19:@89421.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 38:19:@89421.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 38:19:@89421.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 38:19:@89421.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 38:19:@89421.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 38:19:@89421.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 38:19:@89421.4]
  wire  rdata_clock; // @[StreamController.scala 51:21:@89827.4]
  wire  rdata_reset; // @[StreamController.scala 51:21:@89827.4]
  wire  rdata_io_in_ready; // @[StreamController.scala 51:21:@89827.4]
  wire  rdata_io_in_valid; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_0; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_1; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_2; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_3; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_4; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_5; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_6; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_7; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_8; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_9; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_10; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_11; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_12; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_13; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_14; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_15; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_16; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_17; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_18; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_19; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_20; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_21; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_22; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_23; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_24; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_25; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_26; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_27; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_28; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_29; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_30; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_31; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_32; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_33; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_34; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_35; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_36; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_37; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_38; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_39; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_40; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_41; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_42; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_43; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_44; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_45; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_46; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_47; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_48; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_49; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_50; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_51; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_52; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_53; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_54; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_55; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_56; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_57; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_58; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_59; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_60; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_61; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_62; // @[StreamController.scala 51:21:@89827.4]
  wire [7:0] rdata_io_in_bits_data_63; // @[StreamController.scala 51:21:@89827.4]
  wire  rdata_io_out_ready; // @[StreamController.scala 51:21:@89827.4]
  wire  rdata_io_out_valid; // @[StreamController.scala 51:21:@89827.4]
  wire [31:0] rdata_io_out_bits_data_0; // @[StreamController.scala 51:21:@89827.4]
  wire [25:0] _T_95; // @[StreamController.scala 21:10:@89824.4]
  FIFO cmd ( // @[StreamController.scala 38:19:@89421.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert rdata ( // @[StreamController.scala 51:21:@89827.4]
    .clock(rdata_clock),
    .reset(rdata_reset),
    .io_in_ready(rdata_io_in_ready),
    .io_in_valid(rdata_io_in_valid),
    .io_in_bits_data_0(rdata_io_in_bits_data_0),
    .io_in_bits_data_1(rdata_io_in_bits_data_1),
    .io_in_bits_data_2(rdata_io_in_bits_data_2),
    .io_in_bits_data_3(rdata_io_in_bits_data_3),
    .io_in_bits_data_4(rdata_io_in_bits_data_4),
    .io_in_bits_data_5(rdata_io_in_bits_data_5),
    .io_in_bits_data_6(rdata_io_in_bits_data_6),
    .io_in_bits_data_7(rdata_io_in_bits_data_7),
    .io_in_bits_data_8(rdata_io_in_bits_data_8),
    .io_in_bits_data_9(rdata_io_in_bits_data_9),
    .io_in_bits_data_10(rdata_io_in_bits_data_10),
    .io_in_bits_data_11(rdata_io_in_bits_data_11),
    .io_in_bits_data_12(rdata_io_in_bits_data_12),
    .io_in_bits_data_13(rdata_io_in_bits_data_13),
    .io_in_bits_data_14(rdata_io_in_bits_data_14),
    .io_in_bits_data_15(rdata_io_in_bits_data_15),
    .io_in_bits_data_16(rdata_io_in_bits_data_16),
    .io_in_bits_data_17(rdata_io_in_bits_data_17),
    .io_in_bits_data_18(rdata_io_in_bits_data_18),
    .io_in_bits_data_19(rdata_io_in_bits_data_19),
    .io_in_bits_data_20(rdata_io_in_bits_data_20),
    .io_in_bits_data_21(rdata_io_in_bits_data_21),
    .io_in_bits_data_22(rdata_io_in_bits_data_22),
    .io_in_bits_data_23(rdata_io_in_bits_data_23),
    .io_in_bits_data_24(rdata_io_in_bits_data_24),
    .io_in_bits_data_25(rdata_io_in_bits_data_25),
    .io_in_bits_data_26(rdata_io_in_bits_data_26),
    .io_in_bits_data_27(rdata_io_in_bits_data_27),
    .io_in_bits_data_28(rdata_io_in_bits_data_28),
    .io_in_bits_data_29(rdata_io_in_bits_data_29),
    .io_in_bits_data_30(rdata_io_in_bits_data_30),
    .io_in_bits_data_31(rdata_io_in_bits_data_31),
    .io_in_bits_data_32(rdata_io_in_bits_data_32),
    .io_in_bits_data_33(rdata_io_in_bits_data_33),
    .io_in_bits_data_34(rdata_io_in_bits_data_34),
    .io_in_bits_data_35(rdata_io_in_bits_data_35),
    .io_in_bits_data_36(rdata_io_in_bits_data_36),
    .io_in_bits_data_37(rdata_io_in_bits_data_37),
    .io_in_bits_data_38(rdata_io_in_bits_data_38),
    .io_in_bits_data_39(rdata_io_in_bits_data_39),
    .io_in_bits_data_40(rdata_io_in_bits_data_40),
    .io_in_bits_data_41(rdata_io_in_bits_data_41),
    .io_in_bits_data_42(rdata_io_in_bits_data_42),
    .io_in_bits_data_43(rdata_io_in_bits_data_43),
    .io_in_bits_data_44(rdata_io_in_bits_data_44),
    .io_in_bits_data_45(rdata_io_in_bits_data_45),
    .io_in_bits_data_46(rdata_io_in_bits_data_46),
    .io_in_bits_data_47(rdata_io_in_bits_data_47),
    .io_in_bits_data_48(rdata_io_in_bits_data_48),
    .io_in_bits_data_49(rdata_io_in_bits_data_49),
    .io_in_bits_data_50(rdata_io_in_bits_data_50),
    .io_in_bits_data_51(rdata_io_in_bits_data_51),
    .io_in_bits_data_52(rdata_io_in_bits_data_52),
    .io_in_bits_data_53(rdata_io_in_bits_data_53),
    .io_in_bits_data_54(rdata_io_in_bits_data_54),
    .io_in_bits_data_55(rdata_io_in_bits_data_55),
    .io_in_bits_data_56(rdata_io_in_bits_data_56),
    .io_in_bits_data_57(rdata_io_in_bits_data_57),
    .io_in_bits_data_58(rdata_io_in_bits_data_58),
    .io_in_bits_data_59(rdata_io_in_bits_data_59),
    .io_in_bits_data_60(rdata_io_in_bits_data_60),
    .io_in_bits_data_61(rdata_io_in_bits_data_61),
    .io_in_bits_data_62(rdata_io_in_bits_data_62),
    .io_in_bits_data_63(rdata_io_in_bits_data_63),
    .io_out_ready(rdata_io_out_ready),
    .io_out_valid(rdata_io_out_valid),
    .io_out_bits_data_0(rdata_io_out_bits_data_0)
  );
  assign _T_95 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@89824.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 44:21:@89821.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 46:25:@89822.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_95}; // @[StreamController.scala 48:25:@89825.4]
  assign io_dram_rresp_ready = rdata_io_in_ready; // @[StreamController.scala 55:23:@89966.4]
  assign io_load_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 42:21:@89819.4]
  assign io_load_data_valid = rdata_io_out_valid; // @[StreamController.scala 57:22:@89967.4]
  assign io_load_data_bits_rdata_0 = rdata_io_out_bits_data_0; // @[StreamController.scala 58:27:@89968.4]
  assign cmd_clock = clock; // @[:@89422.4]
  assign cmd_reset = reset; // @[:@89423.4]
  assign cmd_io_in_valid = io_load_cmd_valid; // @[StreamController.scala 40:19:@89816.4]
  assign cmd_io_in_bits_addr = io_load_cmd_bits_addr; // @[StreamController.scala 41:18:@89818.4]
  assign cmd_io_in_bits_size = io_load_cmd_bits_size; // @[StreamController.scala 41:18:@89817.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 43:20:@89820.4]
  assign rdata_clock = clock; // @[:@89828.4]
  assign rdata_reset = reset; // @[:@89829.4]
  assign rdata_io_in_valid = io_dram_rresp_valid; // @[StreamController.scala 54:21:@89965.4]
  assign rdata_io_in_bits_data_0 = io_dram_rresp_bits_rdata_0; // @[StreamController.scala 53:25:@89901.4]
  assign rdata_io_in_bits_data_1 = io_dram_rresp_bits_rdata_1; // @[StreamController.scala 53:25:@89902.4]
  assign rdata_io_in_bits_data_2 = io_dram_rresp_bits_rdata_2; // @[StreamController.scala 53:25:@89903.4]
  assign rdata_io_in_bits_data_3 = io_dram_rresp_bits_rdata_3; // @[StreamController.scala 53:25:@89904.4]
  assign rdata_io_in_bits_data_4 = io_dram_rresp_bits_rdata_4; // @[StreamController.scala 53:25:@89905.4]
  assign rdata_io_in_bits_data_5 = io_dram_rresp_bits_rdata_5; // @[StreamController.scala 53:25:@89906.4]
  assign rdata_io_in_bits_data_6 = io_dram_rresp_bits_rdata_6; // @[StreamController.scala 53:25:@89907.4]
  assign rdata_io_in_bits_data_7 = io_dram_rresp_bits_rdata_7; // @[StreamController.scala 53:25:@89908.4]
  assign rdata_io_in_bits_data_8 = io_dram_rresp_bits_rdata_8; // @[StreamController.scala 53:25:@89909.4]
  assign rdata_io_in_bits_data_9 = io_dram_rresp_bits_rdata_9; // @[StreamController.scala 53:25:@89910.4]
  assign rdata_io_in_bits_data_10 = io_dram_rresp_bits_rdata_10; // @[StreamController.scala 53:25:@89911.4]
  assign rdata_io_in_bits_data_11 = io_dram_rresp_bits_rdata_11; // @[StreamController.scala 53:25:@89912.4]
  assign rdata_io_in_bits_data_12 = io_dram_rresp_bits_rdata_12; // @[StreamController.scala 53:25:@89913.4]
  assign rdata_io_in_bits_data_13 = io_dram_rresp_bits_rdata_13; // @[StreamController.scala 53:25:@89914.4]
  assign rdata_io_in_bits_data_14 = io_dram_rresp_bits_rdata_14; // @[StreamController.scala 53:25:@89915.4]
  assign rdata_io_in_bits_data_15 = io_dram_rresp_bits_rdata_15; // @[StreamController.scala 53:25:@89916.4]
  assign rdata_io_in_bits_data_16 = io_dram_rresp_bits_rdata_16; // @[StreamController.scala 53:25:@89917.4]
  assign rdata_io_in_bits_data_17 = io_dram_rresp_bits_rdata_17; // @[StreamController.scala 53:25:@89918.4]
  assign rdata_io_in_bits_data_18 = io_dram_rresp_bits_rdata_18; // @[StreamController.scala 53:25:@89919.4]
  assign rdata_io_in_bits_data_19 = io_dram_rresp_bits_rdata_19; // @[StreamController.scala 53:25:@89920.4]
  assign rdata_io_in_bits_data_20 = io_dram_rresp_bits_rdata_20; // @[StreamController.scala 53:25:@89921.4]
  assign rdata_io_in_bits_data_21 = io_dram_rresp_bits_rdata_21; // @[StreamController.scala 53:25:@89922.4]
  assign rdata_io_in_bits_data_22 = io_dram_rresp_bits_rdata_22; // @[StreamController.scala 53:25:@89923.4]
  assign rdata_io_in_bits_data_23 = io_dram_rresp_bits_rdata_23; // @[StreamController.scala 53:25:@89924.4]
  assign rdata_io_in_bits_data_24 = io_dram_rresp_bits_rdata_24; // @[StreamController.scala 53:25:@89925.4]
  assign rdata_io_in_bits_data_25 = io_dram_rresp_bits_rdata_25; // @[StreamController.scala 53:25:@89926.4]
  assign rdata_io_in_bits_data_26 = io_dram_rresp_bits_rdata_26; // @[StreamController.scala 53:25:@89927.4]
  assign rdata_io_in_bits_data_27 = io_dram_rresp_bits_rdata_27; // @[StreamController.scala 53:25:@89928.4]
  assign rdata_io_in_bits_data_28 = io_dram_rresp_bits_rdata_28; // @[StreamController.scala 53:25:@89929.4]
  assign rdata_io_in_bits_data_29 = io_dram_rresp_bits_rdata_29; // @[StreamController.scala 53:25:@89930.4]
  assign rdata_io_in_bits_data_30 = io_dram_rresp_bits_rdata_30; // @[StreamController.scala 53:25:@89931.4]
  assign rdata_io_in_bits_data_31 = io_dram_rresp_bits_rdata_31; // @[StreamController.scala 53:25:@89932.4]
  assign rdata_io_in_bits_data_32 = io_dram_rresp_bits_rdata_32; // @[StreamController.scala 53:25:@89933.4]
  assign rdata_io_in_bits_data_33 = io_dram_rresp_bits_rdata_33; // @[StreamController.scala 53:25:@89934.4]
  assign rdata_io_in_bits_data_34 = io_dram_rresp_bits_rdata_34; // @[StreamController.scala 53:25:@89935.4]
  assign rdata_io_in_bits_data_35 = io_dram_rresp_bits_rdata_35; // @[StreamController.scala 53:25:@89936.4]
  assign rdata_io_in_bits_data_36 = io_dram_rresp_bits_rdata_36; // @[StreamController.scala 53:25:@89937.4]
  assign rdata_io_in_bits_data_37 = io_dram_rresp_bits_rdata_37; // @[StreamController.scala 53:25:@89938.4]
  assign rdata_io_in_bits_data_38 = io_dram_rresp_bits_rdata_38; // @[StreamController.scala 53:25:@89939.4]
  assign rdata_io_in_bits_data_39 = io_dram_rresp_bits_rdata_39; // @[StreamController.scala 53:25:@89940.4]
  assign rdata_io_in_bits_data_40 = io_dram_rresp_bits_rdata_40; // @[StreamController.scala 53:25:@89941.4]
  assign rdata_io_in_bits_data_41 = io_dram_rresp_bits_rdata_41; // @[StreamController.scala 53:25:@89942.4]
  assign rdata_io_in_bits_data_42 = io_dram_rresp_bits_rdata_42; // @[StreamController.scala 53:25:@89943.4]
  assign rdata_io_in_bits_data_43 = io_dram_rresp_bits_rdata_43; // @[StreamController.scala 53:25:@89944.4]
  assign rdata_io_in_bits_data_44 = io_dram_rresp_bits_rdata_44; // @[StreamController.scala 53:25:@89945.4]
  assign rdata_io_in_bits_data_45 = io_dram_rresp_bits_rdata_45; // @[StreamController.scala 53:25:@89946.4]
  assign rdata_io_in_bits_data_46 = io_dram_rresp_bits_rdata_46; // @[StreamController.scala 53:25:@89947.4]
  assign rdata_io_in_bits_data_47 = io_dram_rresp_bits_rdata_47; // @[StreamController.scala 53:25:@89948.4]
  assign rdata_io_in_bits_data_48 = io_dram_rresp_bits_rdata_48; // @[StreamController.scala 53:25:@89949.4]
  assign rdata_io_in_bits_data_49 = io_dram_rresp_bits_rdata_49; // @[StreamController.scala 53:25:@89950.4]
  assign rdata_io_in_bits_data_50 = io_dram_rresp_bits_rdata_50; // @[StreamController.scala 53:25:@89951.4]
  assign rdata_io_in_bits_data_51 = io_dram_rresp_bits_rdata_51; // @[StreamController.scala 53:25:@89952.4]
  assign rdata_io_in_bits_data_52 = io_dram_rresp_bits_rdata_52; // @[StreamController.scala 53:25:@89953.4]
  assign rdata_io_in_bits_data_53 = io_dram_rresp_bits_rdata_53; // @[StreamController.scala 53:25:@89954.4]
  assign rdata_io_in_bits_data_54 = io_dram_rresp_bits_rdata_54; // @[StreamController.scala 53:25:@89955.4]
  assign rdata_io_in_bits_data_55 = io_dram_rresp_bits_rdata_55; // @[StreamController.scala 53:25:@89956.4]
  assign rdata_io_in_bits_data_56 = io_dram_rresp_bits_rdata_56; // @[StreamController.scala 53:25:@89957.4]
  assign rdata_io_in_bits_data_57 = io_dram_rresp_bits_rdata_57; // @[StreamController.scala 53:25:@89958.4]
  assign rdata_io_in_bits_data_58 = io_dram_rresp_bits_rdata_58; // @[StreamController.scala 53:25:@89959.4]
  assign rdata_io_in_bits_data_59 = io_dram_rresp_bits_rdata_59; // @[StreamController.scala 53:25:@89960.4]
  assign rdata_io_in_bits_data_60 = io_dram_rresp_bits_rdata_60; // @[StreamController.scala 53:25:@89961.4]
  assign rdata_io_in_bits_data_61 = io_dram_rresp_bits_rdata_61; // @[StreamController.scala 53:25:@89962.4]
  assign rdata_io_in_bits_data_62 = io_dram_rresp_bits_rdata_62; // @[StreamController.scala 53:25:@89963.4]
  assign rdata_io_in_bits_data_63 = io_dram_rresp_bits_rdata_63; // @[StreamController.scala 53:25:@89964.4]
  assign rdata_io_out_ready = io_load_data_ready; // @[StreamController.scala 59:22:@89969.4]
endmodule
module FFRAM( // @[:@94025.2]
  input        clock, // @[:@94026.4]
  input        reset, // @[:@94027.4]
  input  [1:0] io_raddr, // @[:@94028.4]
  input        io_wen, // @[:@94028.4]
  input  [1:0] io_waddr, // @[:@94028.4]
  input        io_wdata, // @[:@94028.4]
  output       io_rdata, // @[:@94028.4]
  input        io_banks_0_wdata_valid, // @[:@94028.4]
  input        io_banks_0_wdata_bits, // @[:@94028.4]
  input        io_banks_1_wdata_valid, // @[:@94028.4]
  input        io_banks_1_wdata_bits, // @[:@94028.4]
  input        io_banks_2_wdata_valid, // @[:@94028.4]
  input        io_banks_2_wdata_bits, // @[:@94028.4]
  input        io_banks_3_wdata_valid, // @[:@94028.4]
  input        io_banks_3_wdata_bits // @[:@94028.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@94032.4]
  reg [31:0] _RAND_0;
  wire  _T_88; // @[SRAM.scala 148:37:@94033.4]
  wire  _T_89; // @[SRAM.scala 148:25:@94034.4]
  wire  _T_90; // @[SRAM.scala 148:15:@94035.4]
  wire  _T_91; // @[SRAM.scala 149:15:@94037.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@94036.4]
  reg  regs_1; // @[SRAM.scala 145:20:@94043.4]
  reg [31:0] _RAND_1;
  wire  _T_97; // @[SRAM.scala 148:37:@94044.4]
  wire  _T_98; // @[SRAM.scala 148:25:@94045.4]
  wire  _T_99; // @[SRAM.scala 148:15:@94046.4]
  wire  _T_100; // @[SRAM.scala 149:15:@94048.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@94047.4]
  reg  regs_2; // @[SRAM.scala 145:20:@94054.4]
  reg [31:0] _RAND_2;
  wire  _T_106; // @[SRAM.scala 148:37:@94055.4]
  wire  _T_107; // @[SRAM.scala 148:25:@94056.4]
  wire  _T_108; // @[SRAM.scala 148:15:@94057.4]
  wire  _T_109; // @[SRAM.scala 149:15:@94059.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@94058.4]
  reg  regs_3; // @[SRAM.scala 145:20:@94065.4]
  reg [31:0] _RAND_3;
  wire  _T_115; // @[SRAM.scala 148:37:@94066.4]
  wire  _T_116; // @[SRAM.scala 148:25:@94067.4]
  wire  _T_117; // @[SRAM.scala 148:15:@94068.4]
  wire  _T_118; // @[SRAM.scala 149:15:@94070.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@94069.4]
  wire  _GEN_5; // @[SRAM.scala 155:12:@94079.4]
  wire  _GEN_6; // @[SRAM.scala 155:12:@94079.4]
  assign _T_88 = io_waddr == 2'h0; // @[SRAM.scala 148:37:@94033.4]
  assign _T_89 = io_wen & _T_88; // @[SRAM.scala 148:25:@94034.4]
  assign _T_90 = io_banks_0_wdata_valid | _T_89; // @[SRAM.scala 148:15:@94035.4]
  assign _T_91 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@94037.6]
  assign _GEN_0 = _T_90 ? _T_91 : regs_0; // @[SRAM.scala 148:48:@94036.4]
  assign _T_97 = io_waddr == 2'h1; // @[SRAM.scala 148:37:@94044.4]
  assign _T_98 = io_wen & _T_97; // @[SRAM.scala 148:25:@94045.4]
  assign _T_99 = io_banks_1_wdata_valid | _T_98; // @[SRAM.scala 148:15:@94046.4]
  assign _T_100 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@94048.6]
  assign _GEN_1 = _T_99 ? _T_100 : regs_1; // @[SRAM.scala 148:48:@94047.4]
  assign _T_106 = io_waddr == 2'h2; // @[SRAM.scala 148:37:@94055.4]
  assign _T_107 = io_wen & _T_106; // @[SRAM.scala 148:25:@94056.4]
  assign _T_108 = io_banks_2_wdata_valid | _T_107; // @[SRAM.scala 148:15:@94057.4]
  assign _T_109 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@94059.6]
  assign _GEN_2 = _T_108 ? _T_109 : regs_2; // @[SRAM.scala 148:48:@94058.4]
  assign _T_115 = io_waddr == 2'h3; // @[SRAM.scala 148:37:@94066.4]
  assign _T_116 = io_wen & _T_115; // @[SRAM.scala 148:25:@94067.4]
  assign _T_117 = io_banks_3_wdata_valid | _T_116; // @[SRAM.scala 148:15:@94068.4]
  assign _T_118 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@94070.6]
  assign _GEN_3 = _T_117 ? _T_118 : regs_3; // @[SRAM.scala 148:48:@94069.4]
  assign _GEN_5 = 2'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@94079.4]
  assign _GEN_6 = 2'h2 == io_raddr ? regs_2 : _GEN_5; // @[SRAM.scala 155:12:@94079.4]
  assign io_rdata = 2'h3 == io_raddr ? regs_3 : _GEN_6; // @[SRAM.scala 155:12:@94079.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_90) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_99) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_108) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_117) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_35( // @[:@94081.2]
  input   clock, // @[:@94082.4]
  input   reset, // @[:@94083.4]
  output  io_in_ready, // @[:@94084.4]
  input   io_in_valid, // @[:@94084.4]
  input   io_in_bits, // @[:@94084.4]
  input   io_out_ready, // @[:@94084.4]
  output  io_out_valid, // @[:@94084.4]
  output  io_out_bits // @[:@94084.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@94110.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@94110.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@94110.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@94110.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@94110.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@94110.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@94110.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@94120.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@94120.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@94120.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@94120.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@94120.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@94120.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@94120.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@94135.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@94135.4]
  wire [1:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@94135.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@94135.4]
  wire [1:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@94135.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@94135.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@94135.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@94135.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@94135.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@94135.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@94135.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@94135.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@94135.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@94135.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@94135.4]
  wire  writeEn; // @[FIFO.scala 30:29:@94108.4]
  wire  readEn; // @[FIFO.scala 31:29:@94109.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@94130.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@94131.4]
  wire  _T_104; // @[FIFO.scala 45:27:@94132.4]
  wire  empty; // @[FIFO.scala 45:24:@94133.4]
  wire  full; // @[FIFO.scala 46:23:@94134.4]
  wire  _T_157; // @[FIFO.scala 83:17:@94221.4]
  wire  _GEN_4; // @[FIFO.scala 83:29:@94222.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@94110.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@94120.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM FFRAM ( // @[FIFO.scala 49:19:@94135.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@94108.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@94109.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@94131.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@94132.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@94133.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@94134.4]
  assign _T_157 = writeEn != readEn; // @[FIFO.scala 83:17:@94221.4]
  assign _GEN_4 = _T_157 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@94222.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@94228.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@94226.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@94160.4]
  assign enqCounter_clock = clock; // @[:@94111.4]
  assign enqCounter_reset = reset; // @[:@94112.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@94118.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@94119.4]
  assign deqCounter_clock = clock; // @[:@94121.4]
  assign deqCounter_reset = reset; // @[:@94122.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@94128.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@94129.4]
  assign FFRAM_clock = clock; // @[:@94136.4]
  assign FFRAM_reset = reset; // @[:@94137.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@94156.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@94157.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@94158.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@94159.4]
  assign FFRAM_io_banks_0_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@94162.4]
  assign FFRAM_io_banks_0_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@94161.4]
  assign FFRAM_io_banks_1_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@94165.4]
  assign FFRAM_io_banks_1_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@94164.4]
  assign FFRAM_io_banks_2_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@94168.4]
  assign FFRAM_io_banks_2_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@94167.4]
  assign FFRAM_io_banks_3_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@94171.4]
  assign FFRAM_io_banks_3_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@94170.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_157) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_3( // @[:@97845.2]
  input   clock, // @[:@97846.4]
  input   reset, // @[:@97847.4]
  output  io_in_ready, // @[:@97848.4]
  input   io_in_valid, // @[:@97848.4]
  input   io_in_bits_0, // @[:@97848.4]
  input   io_out_ready, // @[:@97848.4]
  output  io_out_valid, // @[:@97848.4]
  output  io_out_bits_0, // @[:@97848.4]
  output  io_out_bits_1, // @[:@97848.4]
  output  io_out_bits_2, // @[:@97848.4]
  output  io_out_bits_3, // @[:@97848.4]
  output  io_out_bits_4, // @[:@97848.4]
  output  io_out_bits_5, // @[:@97848.4]
  output  io_out_bits_6, // @[:@97848.4]
  output  io_out_bits_7, // @[:@97848.4]
  output  io_out_bits_8, // @[:@97848.4]
  output  io_out_bits_9, // @[:@97848.4]
  output  io_out_bits_10, // @[:@97848.4]
  output  io_out_bits_11, // @[:@97848.4]
  output  io_out_bits_12, // @[:@97848.4]
  output  io_out_bits_13, // @[:@97848.4]
  output  io_out_bits_14, // @[:@97848.4]
  output  io_out_bits_15 // @[:@97848.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@97852.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@97852.4]
  wire  enqCounter_io_reset; // @[FIFOVec.scala 24:26:@97852.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@97852.4]
  wire [3:0] enqCounter_io_stride; // @[FIFOVec.scala 24:26:@97852.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@97852.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@97863.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@97863.4]
  wire  deqCounter_io_reset; // @[FIFOVec.scala 28:26:@97863.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@97863.4]
  wire [3:0] deqCounter_io_stride; // @[FIFOVec.scala 28:26:@97863.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@97863.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@97876.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@97876.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@97876.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@97876.4]
  wire  fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@97876.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@97876.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@97876.4]
  wire  fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@97876.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@97911.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@97911.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@97911.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@97911.4]
  wire  fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@97911.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@97911.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@97911.4]
  wire  fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@97911.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@97946.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@97946.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@97946.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@97946.4]
  wire  fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@97946.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@97946.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@97946.4]
  wire  fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@97946.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@97981.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@97981.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@97981.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@97981.4]
  wire  fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@97981.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@97981.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@97981.4]
  wire  fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@97981.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@98016.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@98016.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@98016.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@98016.4]
  wire  fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@98016.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@98016.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@98016.4]
  wire  fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@98016.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@98051.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@98051.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@98051.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@98051.4]
  wire  fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@98051.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@98051.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@98051.4]
  wire  fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@98051.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@98086.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@98086.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@98086.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@98086.4]
  wire  fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@98086.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@98086.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@98086.4]
  wire  fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@98086.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@98121.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@98121.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@98121.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@98121.4]
  wire  fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@98121.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@98121.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@98121.4]
  wire  fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@98121.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@98156.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@98156.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@98156.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@98156.4]
  wire  fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@98156.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@98156.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@98156.4]
  wire  fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@98156.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@98191.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@98191.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@98191.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@98191.4]
  wire  fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@98191.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@98191.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@98191.4]
  wire  fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@98191.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@98226.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@98226.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@98226.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@98226.4]
  wire  fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@98226.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@98226.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@98226.4]
  wire  fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@98226.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@98261.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@98261.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@98261.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@98261.4]
  wire  fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@98261.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@98261.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@98261.4]
  wire  fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@98261.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@98296.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@98296.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@98296.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@98296.4]
  wire  fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@98296.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@98296.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@98296.4]
  wire  fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@98296.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@98331.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@98331.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@98331.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@98331.4]
  wire  fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@98331.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@98331.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@98331.4]
  wire  fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@98331.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@98366.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@98366.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@98366.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@98366.4]
  wire  fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@98366.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@98366.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@98366.4]
  wire  fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@98366.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@98401.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@98401.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@98401.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@98401.4]
  wire  fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@98401.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@98401.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@98401.4]
  wire  fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@98401.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@97851.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@97874.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@97901.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@97936.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@97971.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@98006.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@98041.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@98076.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@98111.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@98146.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@98181.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@98216.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@98251.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@98286.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@98321.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@98356.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@98391.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@98426.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98437.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98438.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@98468.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98439.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@98468.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98440.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@98468.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98441.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@98468.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98442.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@98468.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98443.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@98468.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98444.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@98468.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98445.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@98468.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98446.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@98468.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98447.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@98468.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98448.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@98468.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98449.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@98468.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98450.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@98468.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98451.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@98468.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98452.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@98487.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@98488.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@98489.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@98490.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@98491.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@98492.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@98493.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@98494.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@98495.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@98496.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@98497.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@98498.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@98499.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@98500.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@97852.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@97863.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out)
  );
  FIFO_35 fifos_0 ( // @[FIFOVec.scala 40:19:@97876.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_35 fifos_1 ( // @[FIFOVec.scala 40:19:@97911.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_35 fifos_2 ( // @[FIFOVec.scala 40:19:@97946.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_35 fifos_3 ( // @[FIFOVec.scala 40:19:@97981.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_35 fifos_4 ( // @[FIFOVec.scala 40:19:@98016.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_35 fifos_5 ( // @[FIFOVec.scala 40:19:@98051.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_35 fifos_6 ( // @[FIFOVec.scala 40:19:@98086.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_35 fifos_7 ( // @[FIFOVec.scala 40:19:@98121.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_35 fifos_8 ( // @[FIFOVec.scala 40:19:@98156.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_35 fifos_9 ( // @[FIFOVec.scala 40:19:@98191.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_35 fifos_10 ( // @[FIFOVec.scala 40:19:@98226.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_35 fifos_11 ( // @[FIFOVec.scala 40:19:@98261.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_35 fifos_12 ( // @[FIFOVec.scala 40:19:@98296.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_35 fifos_13 ( // @[FIFOVec.scala 40:19:@98331.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_35 fifos_14 ( // @[FIFOVec.scala 40:19:@98366.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_35 fifos_15 ( // @[FIFOVec.scala 40:19:@98401.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@97851.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@97874.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@97901.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@97936.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@97971.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@98006.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@98041.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@98076.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@98111.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@98146.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@98181.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@98216.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@98251.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@98286.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@98321.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@98356.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@98391.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@98426.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98437.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98438.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@98468.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98439.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@98468.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98440.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@98468.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98441.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@98468.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98442.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@98468.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98443.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@98468.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98444.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@98468.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98445.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@98468.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98446.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@98468.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98447.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@98468.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98448.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@98468.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98449.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@98468.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98450.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@98468.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98451.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@98468.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@98436.4 FIFOVec.scala 49:42:@98452.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@98487.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@98488.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@98489.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@98490.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@98491.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@98492.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@98493.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@98494.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@98495.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@98496.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@98497.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@98498.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@98499.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@98500.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@98469.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@98503.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@98811.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@98812.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@98813.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@98814.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@98815.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@98816.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@98817.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@98818.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@98819.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@98820.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@98821.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@98822.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@98823.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@98824.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@98825.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@98826.4]
  assign enqCounter_clock = clock; // @[:@97853.4]
  assign enqCounter_reset = reset; // @[:@97854.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@97861.4]
  assign enqCounter_io_stride = 4'h1; // @[FIFOVec.scala 27:24:@97862.4]
  assign deqCounter_clock = clock; // @[:@97864.4]
  assign deqCounter_reset = reset; // @[:@97865.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@97872.4]
  assign deqCounter_io_stride = 4'h1; // @[FIFOVec.scala 31:24:@97873.4]
  assign fifos_0_clock = clock; // @[:@97877.4]
  assign fifos_0_reset = reset; // @[:@97878.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@97904.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@97906.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@97910.4]
  assign fifos_1_clock = clock; // @[:@97912.4]
  assign fifos_1_reset = reset; // @[:@97913.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@97939.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@97941.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@97945.4]
  assign fifos_2_clock = clock; // @[:@97947.4]
  assign fifos_2_reset = reset; // @[:@97948.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@97974.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@97976.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@97980.4]
  assign fifos_3_clock = clock; // @[:@97982.4]
  assign fifos_3_reset = reset; // @[:@97983.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@98009.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@98011.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@98015.4]
  assign fifos_4_clock = clock; // @[:@98017.4]
  assign fifos_4_reset = reset; // @[:@98018.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@98044.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@98046.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@98050.4]
  assign fifos_5_clock = clock; // @[:@98052.4]
  assign fifos_5_reset = reset; // @[:@98053.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@98079.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@98081.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@98085.4]
  assign fifos_6_clock = clock; // @[:@98087.4]
  assign fifos_6_reset = reset; // @[:@98088.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@98114.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@98116.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@98120.4]
  assign fifos_7_clock = clock; // @[:@98122.4]
  assign fifos_7_reset = reset; // @[:@98123.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@98149.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@98151.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@98155.4]
  assign fifos_8_clock = clock; // @[:@98157.4]
  assign fifos_8_reset = reset; // @[:@98158.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@98184.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@98186.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@98190.4]
  assign fifos_9_clock = clock; // @[:@98192.4]
  assign fifos_9_reset = reset; // @[:@98193.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@98219.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@98221.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@98225.4]
  assign fifos_10_clock = clock; // @[:@98227.4]
  assign fifos_10_reset = reset; // @[:@98228.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@98254.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@98256.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@98260.4]
  assign fifos_11_clock = clock; // @[:@98262.4]
  assign fifos_11_reset = reset; // @[:@98263.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@98289.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@98291.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@98295.4]
  assign fifos_12_clock = clock; // @[:@98297.4]
  assign fifos_12_reset = reset; // @[:@98298.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@98324.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@98326.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@98330.4]
  assign fifos_13_clock = clock; // @[:@98332.4]
  assign fifos_13_reset = reset; // @[:@98333.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@98359.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@98361.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@98365.4]
  assign fifos_14_clock = clock; // @[:@98367.4]
  assign fifos_14_reset = reset; // @[:@98368.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@98394.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@98396.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@98400.4]
  assign fifos_15_clock = clock; // @[:@98402.4]
  assign fifos_15_reset = reset; // @[:@98403.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@98429.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@98431.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@98435.4]
endmodule
module FIFOWidthConvert_1( // @[:@98828.2]
  input         clock, // @[:@98829.4]
  input         reset, // @[:@98830.4]
  output        io_in_ready, // @[:@98831.4]
  input         io_in_valid, // @[:@98831.4]
  input  [31:0] io_in_bits_data_0, // @[:@98831.4]
  input         io_in_bits_strobe, // @[:@98831.4]
  input         io_out_ready, // @[:@98831.4]
  output        io_out_valid, // @[:@98831.4]
  output [7:0]  io_out_bits_data_0, // @[:@98831.4]
  output [7:0]  io_out_bits_data_1, // @[:@98831.4]
  output [7:0]  io_out_bits_data_2, // @[:@98831.4]
  output [7:0]  io_out_bits_data_3, // @[:@98831.4]
  output [7:0]  io_out_bits_data_4, // @[:@98831.4]
  output [7:0]  io_out_bits_data_5, // @[:@98831.4]
  output [7:0]  io_out_bits_data_6, // @[:@98831.4]
  output [7:0]  io_out_bits_data_7, // @[:@98831.4]
  output [7:0]  io_out_bits_data_8, // @[:@98831.4]
  output [7:0]  io_out_bits_data_9, // @[:@98831.4]
  output [7:0]  io_out_bits_data_10, // @[:@98831.4]
  output [7:0]  io_out_bits_data_11, // @[:@98831.4]
  output [7:0]  io_out_bits_data_12, // @[:@98831.4]
  output [7:0]  io_out_bits_data_13, // @[:@98831.4]
  output [7:0]  io_out_bits_data_14, // @[:@98831.4]
  output [7:0]  io_out_bits_data_15, // @[:@98831.4]
  output [7:0]  io_out_bits_data_16, // @[:@98831.4]
  output [7:0]  io_out_bits_data_17, // @[:@98831.4]
  output [7:0]  io_out_bits_data_18, // @[:@98831.4]
  output [7:0]  io_out_bits_data_19, // @[:@98831.4]
  output [7:0]  io_out_bits_data_20, // @[:@98831.4]
  output [7:0]  io_out_bits_data_21, // @[:@98831.4]
  output [7:0]  io_out_bits_data_22, // @[:@98831.4]
  output [7:0]  io_out_bits_data_23, // @[:@98831.4]
  output [7:0]  io_out_bits_data_24, // @[:@98831.4]
  output [7:0]  io_out_bits_data_25, // @[:@98831.4]
  output [7:0]  io_out_bits_data_26, // @[:@98831.4]
  output [7:0]  io_out_bits_data_27, // @[:@98831.4]
  output [7:0]  io_out_bits_data_28, // @[:@98831.4]
  output [7:0]  io_out_bits_data_29, // @[:@98831.4]
  output [7:0]  io_out_bits_data_30, // @[:@98831.4]
  output [7:0]  io_out_bits_data_31, // @[:@98831.4]
  output [7:0]  io_out_bits_data_32, // @[:@98831.4]
  output [7:0]  io_out_bits_data_33, // @[:@98831.4]
  output [7:0]  io_out_bits_data_34, // @[:@98831.4]
  output [7:0]  io_out_bits_data_35, // @[:@98831.4]
  output [7:0]  io_out_bits_data_36, // @[:@98831.4]
  output [7:0]  io_out_bits_data_37, // @[:@98831.4]
  output [7:0]  io_out_bits_data_38, // @[:@98831.4]
  output [7:0]  io_out_bits_data_39, // @[:@98831.4]
  output [7:0]  io_out_bits_data_40, // @[:@98831.4]
  output [7:0]  io_out_bits_data_41, // @[:@98831.4]
  output [7:0]  io_out_bits_data_42, // @[:@98831.4]
  output [7:0]  io_out_bits_data_43, // @[:@98831.4]
  output [7:0]  io_out_bits_data_44, // @[:@98831.4]
  output [7:0]  io_out_bits_data_45, // @[:@98831.4]
  output [7:0]  io_out_bits_data_46, // @[:@98831.4]
  output [7:0]  io_out_bits_data_47, // @[:@98831.4]
  output [7:0]  io_out_bits_data_48, // @[:@98831.4]
  output [7:0]  io_out_bits_data_49, // @[:@98831.4]
  output [7:0]  io_out_bits_data_50, // @[:@98831.4]
  output [7:0]  io_out_bits_data_51, // @[:@98831.4]
  output [7:0]  io_out_bits_data_52, // @[:@98831.4]
  output [7:0]  io_out_bits_data_53, // @[:@98831.4]
  output [7:0]  io_out_bits_data_54, // @[:@98831.4]
  output [7:0]  io_out_bits_data_55, // @[:@98831.4]
  output [7:0]  io_out_bits_data_56, // @[:@98831.4]
  output [7:0]  io_out_bits_data_57, // @[:@98831.4]
  output [7:0]  io_out_bits_data_58, // @[:@98831.4]
  output [7:0]  io_out_bits_data_59, // @[:@98831.4]
  output [7:0]  io_out_bits_data_60, // @[:@98831.4]
  output [7:0]  io_out_bits_data_61, // @[:@98831.4]
  output [7:0]  io_out_bits_data_62, // @[:@98831.4]
  output [7:0]  io_out_bits_data_63, // @[:@98831.4]
  output [63:0] io_out_bits_strobe // @[:@98831.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_in_bits_1; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_in_bits_2; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_in_bits_3; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_in_bits_4; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_in_bits_5; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_in_bits_6; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_in_bits_7; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_in_bits_8; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_in_bits_9; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_in_bits_10; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_in_bits_11; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_in_bits_12; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_in_bits_13; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_in_bits_14; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_in_bits_15; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_out_bits_1; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_out_bits_2; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_out_bits_3; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_out_bits_4; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_out_bits_5; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_out_bits_6; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_out_bits_7; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_out_bits_8; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_out_bits_9; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_out_bits_10; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_out_bits_11; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_out_bits_12; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_out_bits_13; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_out_bits_14; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire [31:0] FIFOVec_io_out_bits_15; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire  FIFOVec_io_chainEnq; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire  FIFOVec_io_chainDeq; // @[FIFOWidthConvert.scala 61:22:@98833.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_in_bits_0; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_ready; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_valid; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_bits_0; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_bits_1; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_bits_2; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_bits_3; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_bits_4; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_bits_5; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_bits_6; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_bits_7; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_bits_8; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_bits_9; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_bits_10; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_bits_11; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_bits_12; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_bits_13; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_bits_14; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire  FIFOVec_1_io_out_bits_15; // @[FIFOWidthConvert.scala 62:26:@98874.4]
  wire [319:0] _T_55; // @[Cat.scala 30:58:@98933.4]
  wire [511:0] _T_61; // @[Cat.scala 30:58:@98939.4]
  wire [9:0] _T_204; // @[Cat.scala 30:58:@99141.4]
  wire [15:0] _T_210; // @[Cat.scala 30:58:@99147.4]
  wire  _T_211; // @[FIFOWidthConvert.scala 36:14:@99148.4]
  wire  _T_215; // @[FIFOWidthConvert.scala 36:14:@99152.4]
  wire  _T_219; // @[FIFOWidthConvert.scala 36:14:@99156.4]
  wire  _T_223; // @[FIFOWidthConvert.scala 36:14:@99160.4]
  wire  _T_227; // @[FIFOWidthConvert.scala 36:14:@99164.4]
  wire  _T_231; // @[FIFOWidthConvert.scala 36:14:@99168.4]
  wire  _T_235; // @[FIFOWidthConvert.scala 36:14:@99172.4]
  wire  _T_239; // @[FIFOWidthConvert.scala 36:14:@99176.4]
  wire  _T_243; // @[FIFOWidthConvert.scala 36:14:@99180.4]
  wire  _T_247; // @[FIFOWidthConvert.scala 36:14:@99184.4]
  wire  _T_251; // @[FIFOWidthConvert.scala 36:14:@99188.4]
  wire  _T_255; // @[FIFOWidthConvert.scala 36:14:@99192.4]
  wire  _T_259; // @[FIFOWidthConvert.scala 36:14:@99196.4]
  wire  _T_263; // @[FIFOWidthConvert.scala 36:14:@99200.4]
  wire  _T_267; // @[FIFOWidthConvert.scala 36:14:@99204.4]
  wire  _T_271; // @[FIFOWidthConvert.scala 36:14:@99208.4]
  wire [9:0] _T_353; // @[Cat.scala 30:58:@99285.4]
  wire [18:0] _T_362; // @[Cat.scala 30:58:@99294.4]
  wire [27:0] _T_371; // @[Cat.scala 30:58:@99303.4]
  wire [36:0] _T_380; // @[Cat.scala 30:58:@99312.4]
  wire [45:0] _T_389; // @[Cat.scala 30:58:@99321.4]
  wire [54:0] _T_398; // @[Cat.scala 30:58:@99330.4]
  wire [62:0] _T_406; // @[Cat.scala 30:58:@99338.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 61:22:@98833.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_in_bits_1(FIFOVec_io_in_bits_1),
    .io_in_bits_2(FIFOVec_io_in_bits_2),
    .io_in_bits_3(FIFOVec_io_in_bits_3),
    .io_in_bits_4(FIFOVec_io_in_bits_4),
    .io_in_bits_5(FIFOVec_io_in_bits_5),
    .io_in_bits_6(FIFOVec_io_in_bits_6),
    .io_in_bits_7(FIFOVec_io_in_bits_7),
    .io_in_bits_8(FIFOVec_io_in_bits_8),
    .io_in_bits_9(FIFOVec_io_in_bits_9),
    .io_in_bits_10(FIFOVec_io_in_bits_10),
    .io_in_bits_11(FIFOVec_io_in_bits_11),
    .io_in_bits_12(FIFOVec_io_in_bits_12),
    .io_in_bits_13(FIFOVec_io_in_bits_13),
    .io_in_bits_14(FIFOVec_io_in_bits_14),
    .io_in_bits_15(FIFOVec_io_in_bits_15),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0),
    .io_out_bits_1(FIFOVec_io_out_bits_1),
    .io_out_bits_2(FIFOVec_io_out_bits_2),
    .io_out_bits_3(FIFOVec_io_out_bits_3),
    .io_out_bits_4(FIFOVec_io_out_bits_4),
    .io_out_bits_5(FIFOVec_io_out_bits_5),
    .io_out_bits_6(FIFOVec_io_out_bits_6),
    .io_out_bits_7(FIFOVec_io_out_bits_7),
    .io_out_bits_8(FIFOVec_io_out_bits_8),
    .io_out_bits_9(FIFOVec_io_out_bits_9),
    .io_out_bits_10(FIFOVec_io_out_bits_10),
    .io_out_bits_11(FIFOVec_io_out_bits_11),
    .io_out_bits_12(FIFOVec_io_out_bits_12),
    .io_out_bits_13(FIFOVec_io_out_bits_13),
    .io_out_bits_14(FIFOVec_io_out_bits_14),
    .io_out_bits_15(FIFOVec_io_out_bits_15),
    .io_chainEnq(FIFOVec_io_chainEnq),
    .io_chainDeq(FIFOVec_io_chainDeq)
  );
  FIFOVec_3 FIFOVec_1 ( // @[FIFOWidthConvert.scala 62:26:@98874.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid),
    .io_in_bits_0(FIFOVec_1_io_in_bits_0),
    .io_out_ready(FIFOVec_1_io_out_ready),
    .io_out_valid(FIFOVec_1_io_out_valid),
    .io_out_bits_0(FIFOVec_1_io_out_bits_0),
    .io_out_bits_1(FIFOVec_1_io_out_bits_1),
    .io_out_bits_2(FIFOVec_1_io_out_bits_2),
    .io_out_bits_3(FIFOVec_1_io_out_bits_3),
    .io_out_bits_4(FIFOVec_1_io_out_bits_4),
    .io_out_bits_5(FIFOVec_1_io_out_bits_5),
    .io_out_bits_6(FIFOVec_1_io_out_bits_6),
    .io_out_bits_7(FIFOVec_1_io_out_bits_7),
    .io_out_bits_8(FIFOVec_1_io_out_bits_8),
    .io_out_bits_9(FIFOVec_1_io_out_bits_9),
    .io_out_bits_10(FIFOVec_1_io_out_bits_10),
    .io_out_bits_11(FIFOVec_1_io_out_bits_11),
    .io_out_bits_12(FIFOVec_1_io_out_bits_12),
    .io_out_bits_13(FIFOVec_1_io_out_bits_13),
    .io_out_bits_14(FIFOVec_1_io_out_bits_14),
    .io_out_bits_15(FIFOVec_1_io_out_bits_15)
  );
  assign _T_55 = {FIFOVec_io_out_bits_15,FIFOVec_io_out_bits_14,FIFOVec_io_out_bits_13,FIFOVec_io_out_bits_12,FIFOVec_io_out_bits_11,FIFOVec_io_out_bits_10,FIFOVec_io_out_bits_9,FIFOVec_io_out_bits_8,FIFOVec_io_out_bits_7,FIFOVec_io_out_bits_6}; // @[Cat.scala 30:58:@98933.4]
  assign _T_61 = {_T_55,FIFOVec_io_out_bits_5,FIFOVec_io_out_bits_4,FIFOVec_io_out_bits_3,FIFOVec_io_out_bits_2,FIFOVec_io_out_bits_1,FIFOVec_io_out_bits_0}; // @[Cat.scala 30:58:@98939.4]
  assign _T_204 = {FIFOVec_1_io_out_bits_0,FIFOVec_1_io_out_bits_1,FIFOVec_1_io_out_bits_2,FIFOVec_1_io_out_bits_3,FIFOVec_1_io_out_bits_4,FIFOVec_1_io_out_bits_5,FIFOVec_1_io_out_bits_6,FIFOVec_1_io_out_bits_7,FIFOVec_1_io_out_bits_8,FIFOVec_1_io_out_bits_9}; // @[Cat.scala 30:58:@99141.4]
  assign _T_210 = {_T_204,FIFOVec_1_io_out_bits_10,FIFOVec_1_io_out_bits_11,FIFOVec_1_io_out_bits_12,FIFOVec_1_io_out_bits_13,FIFOVec_1_io_out_bits_14,FIFOVec_1_io_out_bits_15}; // @[Cat.scala 30:58:@99147.4]
  assign _T_211 = _T_210[0]; // @[FIFOWidthConvert.scala 36:14:@99148.4]
  assign _T_215 = _T_210[1]; // @[FIFOWidthConvert.scala 36:14:@99152.4]
  assign _T_219 = _T_210[2]; // @[FIFOWidthConvert.scala 36:14:@99156.4]
  assign _T_223 = _T_210[3]; // @[FIFOWidthConvert.scala 36:14:@99160.4]
  assign _T_227 = _T_210[4]; // @[FIFOWidthConvert.scala 36:14:@99164.4]
  assign _T_231 = _T_210[5]; // @[FIFOWidthConvert.scala 36:14:@99168.4]
  assign _T_235 = _T_210[6]; // @[FIFOWidthConvert.scala 36:14:@99172.4]
  assign _T_239 = _T_210[7]; // @[FIFOWidthConvert.scala 36:14:@99176.4]
  assign _T_243 = _T_210[8]; // @[FIFOWidthConvert.scala 36:14:@99180.4]
  assign _T_247 = _T_210[9]; // @[FIFOWidthConvert.scala 36:14:@99184.4]
  assign _T_251 = _T_210[10]; // @[FIFOWidthConvert.scala 36:14:@99188.4]
  assign _T_255 = _T_210[11]; // @[FIFOWidthConvert.scala 36:14:@99192.4]
  assign _T_259 = _T_210[12]; // @[FIFOWidthConvert.scala 36:14:@99196.4]
  assign _T_263 = _T_210[13]; // @[FIFOWidthConvert.scala 36:14:@99200.4]
  assign _T_267 = _T_210[14]; // @[FIFOWidthConvert.scala 36:14:@99204.4]
  assign _T_271 = _T_210[15]; // @[FIFOWidthConvert.scala 36:14:@99208.4]
  assign _T_353 = {_T_271,_T_271,_T_271,_T_271,_T_267,_T_267,_T_267,_T_267,_T_263,_T_263}; // @[Cat.scala 30:58:@99285.4]
  assign _T_362 = {_T_353,_T_263,_T_263,_T_259,_T_259,_T_259,_T_259,_T_255,_T_255,_T_255}; // @[Cat.scala 30:58:@99294.4]
  assign _T_371 = {_T_362,_T_255,_T_251,_T_251,_T_251,_T_251,_T_247,_T_247,_T_247,_T_247}; // @[Cat.scala 30:58:@99303.4]
  assign _T_380 = {_T_371,_T_243,_T_243,_T_243,_T_243,_T_239,_T_239,_T_239,_T_239,_T_235}; // @[Cat.scala 30:58:@99312.4]
  assign _T_389 = {_T_380,_T_235,_T_235,_T_235,_T_231,_T_231,_T_231,_T_231,_T_227,_T_227}; // @[Cat.scala 30:58:@99321.4]
  assign _T_398 = {_T_389,_T_227,_T_227,_T_223,_T_223,_T_223,_T_223,_T_219,_T_219,_T_219}; // @[Cat.scala 30:58:@99330.4]
  assign _T_406 = {_T_398,_T_219,_T_215,_T_215,_T_215,_T_215,_T_211,_T_211,_T_211}; // @[Cat.scala 30:58:@99338.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 71:17:@98923.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 72:18:@98924.4]
  assign io_out_bits_data_0 = _T_61[7:0]; // @[FIFOWidthConvert.scala 73:22:@99069.4]
  assign io_out_bits_data_1 = _T_61[15:8]; // @[FIFOWidthConvert.scala 73:22:@99070.4]
  assign io_out_bits_data_2 = _T_61[23:16]; // @[FIFOWidthConvert.scala 73:22:@99071.4]
  assign io_out_bits_data_3 = _T_61[31:24]; // @[FIFOWidthConvert.scala 73:22:@99072.4]
  assign io_out_bits_data_4 = _T_61[39:32]; // @[FIFOWidthConvert.scala 73:22:@99073.4]
  assign io_out_bits_data_5 = _T_61[47:40]; // @[FIFOWidthConvert.scala 73:22:@99074.4]
  assign io_out_bits_data_6 = _T_61[55:48]; // @[FIFOWidthConvert.scala 73:22:@99075.4]
  assign io_out_bits_data_7 = _T_61[63:56]; // @[FIFOWidthConvert.scala 73:22:@99076.4]
  assign io_out_bits_data_8 = _T_61[71:64]; // @[FIFOWidthConvert.scala 73:22:@99077.4]
  assign io_out_bits_data_9 = _T_61[79:72]; // @[FIFOWidthConvert.scala 73:22:@99078.4]
  assign io_out_bits_data_10 = _T_61[87:80]; // @[FIFOWidthConvert.scala 73:22:@99079.4]
  assign io_out_bits_data_11 = _T_61[95:88]; // @[FIFOWidthConvert.scala 73:22:@99080.4]
  assign io_out_bits_data_12 = _T_61[103:96]; // @[FIFOWidthConvert.scala 73:22:@99081.4]
  assign io_out_bits_data_13 = _T_61[111:104]; // @[FIFOWidthConvert.scala 73:22:@99082.4]
  assign io_out_bits_data_14 = _T_61[119:112]; // @[FIFOWidthConvert.scala 73:22:@99083.4]
  assign io_out_bits_data_15 = _T_61[127:120]; // @[FIFOWidthConvert.scala 73:22:@99084.4]
  assign io_out_bits_data_16 = _T_61[135:128]; // @[FIFOWidthConvert.scala 73:22:@99085.4]
  assign io_out_bits_data_17 = _T_61[143:136]; // @[FIFOWidthConvert.scala 73:22:@99086.4]
  assign io_out_bits_data_18 = _T_61[151:144]; // @[FIFOWidthConvert.scala 73:22:@99087.4]
  assign io_out_bits_data_19 = _T_61[159:152]; // @[FIFOWidthConvert.scala 73:22:@99088.4]
  assign io_out_bits_data_20 = _T_61[167:160]; // @[FIFOWidthConvert.scala 73:22:@99089.4]
  assign io_out_bits_data_21 = _T_61[175:168]; // @[FIFOWidthConvert.scala 73:22:@99090.4]
  assign io_out_bits_data_22 = _T_61[183:176]; // @[FIFOWidthConvert.scala 73:22:@99091.4]
  assign io_out_bits_data_23 = _T_61[191:184]; // @[FIFOWidthConvert.scala 73:22:@99092.4]
  assign io_out_bits_data_24 = _T_61[199:192]; // @[FIFOWidthConvert.scala 73:22:@99093.4]
  assign io_out_bits_data_25 = _T_61[207:200]; // @[FIFOWidthConvert.scala 73:22:@99094.4]
  assign io_out_bits_data_26 = _T_61[215:208]; // @[FIFOWidthConvert.scala 73:22:@99095.4]
  assign io_out_bits_data_27 = _T_61[223:216]; // @[FIFOWidthConvert.scala 73:22:@99096.4]
  assign io_out_bits_data_28 = _T_61[231:224]; // @[FIFOWidthConvert.scala 73:22:@99097.4]
  assign io_out_bits_data_29 = _T_61[239:232]; // @[FIFOWidthConvert.scala 73:22:@99098.4]
  assign io_out_bits_data_30 = _T_61[247:240]; // @[FIFOWidthConvert.scala 73:22:@99099.4]
  assign io_out_bits_data_31 = _T_61[255:248]; // @[FIFOWidthConvert.scala 73:22:@99100.4]
  assign io_out_bits_data_32 = _T_61[263:256]; // @[FIFOWidthConvert.scala 73:22:@99101.4]
  assign io_out_bits_data_33 = _T_61[271:264]; // @[FIFOWidthConvert.scala 73:22:@99102.4]
  assign io_out_bits_data_34 = _T_61[279:272]; // @[FIFOWidthConvert.scala 73:22:@99103.4]
  assign io_out_bits_data_35 = _T_61[287:280]; // @[FIFOWidthConvert.scala 73:22:@99104.4]
  assign io_out_bits_data_36 = _T_61[295:288]; // @[FIFOWidthConvert.scala 73:22:@99105.4]
  assign io_out_bits_data_37 = _T_61[303:296]; // @[FIFOWidthConvert.scala 73:22:@99106.4]
  assign io_out_bits_data_38 = _T_61[311:304]; // @[FIFOWidthConvert.scala 73:22:@99107.4]
  assign io_out_bits_data_39 = _T_61[319:312]; // @[FIFOWidthConvert.scala 73:22:@99108.4]
  assign io_out_bits_data_40 = _T_61[327:320]; // @[FIFOWidthConvert.scala 73:22:@99109.4]
  assign io_out_bits_data_41 = _T_61[335:328]; // @[FIFOWidthConvert.scala 73:22:@99110.4]
  assign io_out_bits_data_42 = _T_61[343:336]; // @[FIFOWidthConvert.scala 73:22:@99111.4]
  assign io_out_bits_data_43 = _T_61[351:344]; // @[FIFOWidthConvert.scala 73:22:@99112.4]
  assign io_out_bits_data_44 = _T_61[359:352]; // @[FIFOWidthConvert.scala 73:22:@99113.4]
  assign io_out_bits_data_45 = _T_61[367:360]; // @[FIFOWidthConvert.scala 73:22:@99114.4]
  assign io_out_bits_data_46 = _T_61[375:368]; // @[FIFOWidthConvert.scala 73:22:@99115.4]
  assign io_out_bits_data_47 = _T_61[383:376]; // @[FIFOWidthConvert.scala 73:22:@99116.4]
  assign io_out_bits_data_48 = _T_61[391:384]; // @[FIFOWidthConvert.scala 73:22:@99117.4]
  assign io_out_bits_data_49 = _T_61[399:392]; // @[FIFOWidthConvert.scala 73:22:@99118.4]
  assign io_out_bits_data_50 = _T_61[407:400]; // @[FIFOWidthConvert.scala 73:22:@99119.4]
  assign io_out_bits_data_51 = _T_61[415:408]; // @[FIFOWidthConvert.scala 73:22:@99120.4]
  assign io_out_bits_data_52 = _T_61[423:416]; // @[FIFOWidthConvert.scala 73:22:@99121.4]
  assign io_out_bits_data_53 = _T_61[431:424]; // @[FIFOWidthConvert.scala 73:22:@99122.4]
  assign io_out_bits_data_54 = _T_61[439:432]; // @[FIFOWidthConvert.scala 73:22:@99123.4]
  assign io_out_bits_data_55 = _T_61[447:440]; // @[FIFOWidthConvert.scala 73:22:@99124.4]
  assign io_out_bits_data_56 = _T_61[455:448]; // @[FIFOWidthConvert.scala 73:22:@99125.4]
  assign io_out_bits_data_57 = _T_61[463:456]; // @[FIFOWidthConvert.scala 73:22:@99126.4]
  assign io_out_bits_data_58 = _T_61[471:464]; // @[FIFOWidthConvert.scala 73:22:@99127.4]
  assign io_out_bits_data_59 = _T_61[479:472]; // @[FIFOWidthConvert.scala 73:22:@99128.4]
  assign io_out_bits_data_60 = _T_61[487:480]; // @[FIFOWidthConvert.scala 73:22:@99129.4]
  assign io_out_bits_data_61 = _T_61[495:488]; // @[FIFOWidthConvert.scala 73:22:@99130.4]
  assign io_out_bits_data_62 = _T_61[503:496]; // @[FIFOWidthConvert.scala 73:22:@99131.4]
  assign io_out_bits_data_63 = _T_61[511:504]; // @[FIFOWidthConvert.scala 73:22:@99132.4]
  assign io_out_bits_strobe = {_T_406,_T_211}; // @[FIFOWidthConvert.scala 74:24:@99340.4]
  assign FIFOVec_clock = clock; // @[:@98834.4]
  assign FIFOVec_reset = reset; // @[:@98835.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 68:22:@98920.4]
  assign FIFOVec_io_in_bits_0 = io_in_bits_data_0; // @[FIFOWidthConvert.scala 67:24:@98919.4]
  assign FIFOVec_io_in_bits_1 = 32'h0;
  assign FIFOVec_io_in_bits_2 = 32'h0;
  assign FIFOVec_io_in_bits_3 = 32'h0;
  assign FIFOVec_io_in_bits_4 = 32'h0;
  assign FIFOVec_io_in_bits_5 = 32'h0;
  assign FIFOVec_io_in_bits_6 = 32'h0;
  assign FIFOVec_io_in_bits_7 = 32'h0;
  assign FIFOVec_io_in_bits_8 = 32'h0;
  assign FIFOVec_io_in_bits_9 = 32'h0;
  assign FIFOVec_io_in_bits_10 = 32'h0;
  assign FIFOVec_io_in_bits_11 = 32'h0;
  assign FIFOVec_io_in_bits_12 = 32'h0;
  assign FIFOVec_io_in_bits_13 = 32'h0;
  assign FIFOVec_io_in_bits_14 = 32'h0;
  assign FIFOVec_io_in_bits_15 = 32'h0;
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 75:23:@99341.4]
  assign FIFOVec_io_chainEnq = 1'h1; // @[FIFOWidthConvert.scala 63:22:@98915.4]
  assign FIFOVec_io_chainDeq = 1'h0; // @[FIFOWidthConvert.scala 64:22:@98916.4]
  assign FIFOVec_1_clock = clock; // @[:@98875.4]
  assign FIFOVec_1_reset = reset; // @[:@98876.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 70:26:@98922.4]
  assign FIFOVec_1_io_in_bits_0 = io_in_bits_strobe; // @[FIFOWidthConvert.scala 69:28:@98921.4]
  assign FIFOVec_1_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 76:27:@99342.4]
endmodule
module FFRAM_16( // @[:@99380.2]
  input        clock, // @[:@99381.4]
  input        reset, // @[:@99382.4]
  input  [5:0] io_raddr, // @[:@99383.4]
  input        io_wen, // @[:@99383.4]
  input  [5:0] io_waddr, // @[:@99383.4]
  output       io_rdata // @[:@99383.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@99387.4]
  reg [31:0] _RAND_0;
  wire  _T_688; // @[SRAM.scala 148:37:@99388.4]
  wire  _T_689; // @[SRAM.scala 148:25:@99389.4]
  wire  _GEN_0; // @[SRAM.scala 148:48:@99391.4]
  reg  regs_1; // @[SRAM.scala 145:20:@99398.4]
  reg [31:0] _RAND_1;
  wire  _T_697; // @[SRAM.scala 148:37:@99399.4]
  wire  _T_698; // @[SRAM.scala 148:25:@99400.4]
  wire  _GEN_1; // @[SRAM.scala 148:48:@99402.4]
  reg  regs_2; // @[SRAM.scala 145:20:@99409.4]
  reg [31:0] _RAND_2;
  wire  _T_706; // @[SRAM.scala 148:37:@99410.4]
  wire  _T_707; // @[SRAM.scala 148:25:@99411.4]
  wire  _GEN_2; // @[SRAM.scala 148:48:@99413.4]
  reg  regs_3; // @[SRAM.scala 145:20:@99420.4]
  reg [31:0] _RAND_3;
  wire  _T_715; // @[SRAM.scala 148:37:@99421.4]
  wire  _T_716; // @[SRAM.scala 148:25:@99422.4]
  wire  _GEN_3; // @[SRAM.scala 148:48:@99424.4]
  reg  regs_4; // @[SRAM.scala 145:20:@99431.4]
  reg [31:0] _RAND_4;
  wire  _T_724; // @[SRAM.scala 148:37:@99432.4]
  wire  _T_725; // @[SRAM.scala 148:25:@99433.4]
  wire  _GEN_4; // @[SRAM.scala 148:48:@99435.4]
  reg  regs_5; // @[SRAM.scala 145:20:@99442.4]
  reg [31:0] _RAND_5;
  wire  _T_733; // @[SRAM.scala 148:37:@99443.4]
  wire  _T_734; // @[SRAM.scala 148:25:@99444.4]
  wire  _GEN_5; // @[SRAM.scala 148:48:@99446.4]
  reg  regs_6; // @[SRAM.scala 145:20:@99453.4]
  reg [31:0] _RAND_6;
  wire  _T_742; // @[SRAM.scala 148:37:@99454.4]
  wire  _T_743; // @[SRAM.scala 148:25:@99455.4]
  wire  _GEN_6; // @[SRAM.scala 148:48:@99457.4]
  reg  regs_7; // @[SRAM.scala 145:20:@99464.4]
  reg [31:0] _RAND_7;
  wire  _T_751; // @[SRAM.scala 148:37:@99465.4]
  wire  _T_752; // @[SRAM.scala 148:25:@99466.4]
  wire  _GEN_7; // @[SRAM.scala 148:48:@99468.4]
  reg  regs_8; // @[SRAM.scala 145:20:@99475.4]
  reg [31:0] _RAND_8;
  wire  _T_760; // @[SRAM.scala 148:37:@99476.4]
  wire  _T_761; // @[SRAM.scala 148:25:@99477.4]
  wire  _GEN_8; // @[SRAM.scala 148:48:@99479.4]
  reg  regs_9; // @[SRAM.scala 145:20:@99486.4]
  reg [31:0] _RAND_9;
  wire  _T_769; // @[SRAM.scala 148:37:@99487.4]
  wire  _T_770; // @[SRAM.scala 148:25:@99488.4]
  wire  _GEN_9; // @[SRAM.scala 148:48:@99490.4]
  reg  regs_10; // @[SRAM.scala 145:20:@99497.4]
  reg [31:0] _RAND_10;
  wire  _T_778; // @[SRAM.scala 148:37:@99498.4]
  wire  _T_779; // @[SRAM.scala 148:25:@99499.4]
  wire  _GEN_10; // @[SRAM.scala 148:48:@99501.4]
  reg  regs_11; // @[SRAM.scala 145:20:@99508.4]
  reg [31:0] _RAND_11;
  wire  _T_787; // @[SRAM.scala 148:37:@99509.4]
  wire  _T_788; // @[SRAM.scala 148:25:@99510.4]
  wire  _GEN_11; // @[SRAM.scala 148:48:@99512.4]
  reg  regs_12; // @[SRAM.scala 145:20:@99519.4]
  reg [31:0] _RAND_12;
  wire  _T_796; // @[SRAM.scala 148:37:@99520.4]
  wire  _T_797; // @[SRAM.scala 148:25:@99521.4]
  wire  _GEN_12; // @[SRAM.scala 148:48:@99523.4]
  reg  regs_13; // @[SRAM.scala 145:20:@99530.4]
  reg [31:0] _RAND_13;
  wire  _T_805; // @[SRAM.scala 148:37:@99531.4]
  wire  _T_806; // @[SRAM.scala 148:25:@99532.4]
  wire  _GEN_13; // @[SRAM.scala 148:48:@99534.4]
  reg  regs_14; // @[SRAM.scala 145:20:@99541.4]
  reg [31:0] _RAND_14;
  wire  _T_814; // @[SRAM.scala 148:37:@99542.4]
  wire  _T_815; // @[SRAM.scala 148:25:@99543.4]
  wire  _GEN_14; // @[SRAM.scala 148:48:@99545.4]
  reg  regs_15; // @[SRAM.scala 145:20:@99552.4]
  reg [31:0] _RAND_15;
  wire  _T_823; // @[SRAM.scala 148:37:@99553.4]
  wire  _T_824; // @[SRAM.scala 148:25:@99554.4]
  wire  _GEN_15; // @[SRAM.scala 148:48:@99556.4]
  reg  regs_16; // @[SRAM.scala 145:20:@99563.4]
  reg [31:0] _RAND_16;
  wire  _T_832; // @[SRAM.scala 148:37:@99564.4]
  wire  _T_833; // @[SRAM.scala 148:25:@99565.4]
  wire  _GEN_16; // @[SRAM.scala 148:48:@99567.4]
  reg  regs_17; // @[SRAM.scala 145:20:@99574.4]
  reg [31:0] _RAND_17;
  wire  _T_841; // @[SRAM.scala 148:37:@99575.4]
  wire  _T_842; // @[SRAM.scala 148:25:@99576.4]
  wire  _GEN_17; // @[SRAM.scala 148:48:@99578.4]
  reg  regs_18; // @[SRAM.scala 145:20:@99585.4]
  reg [31:0] _RAND_18;
  wire  _T_850; // @[SRAM.scala 148:37:@99586.4]
  wire  _T_851; // @[SRAM.scala 148:25:@99587.4]
  wire  _GEN_18; // @[SRAM.scala 148:48:@99589.4]
  reg  regs_19; // @[SRAM.scala 145:20:@99596.4]
  reg [31:0] _RAND_19;
  wire  _T_859; // @[SRAM.scala 148:37:@99597.4]
  wire  _T_860; // @[SRAM.scala 148:25:@99598.4]
  wire  _GEN_19; // @[SRAM.scala 148:48:@99600.4]
  reg  regs_20; // @[SRAM.scala 145:20:@99607.4]
  reg [31:0] _RAND_20;
  wire  _T_868; // @[SRAM.scala 148:37:@99608.4]
  wire  _T_869; // @[SRAM.scala 148:25:@99609.4]
  wire  _GEN_20; // @[SRAM.scala 148:48:@99611.4]
  reg  regs_21; // @[SRAM.scala 145:20:@99618.4]
  reg [31:0] _RAND_21;
  wire  _T_877; // @[SRAM.scala 148:37:@99619.4]
  wire  _T_878; // @[SRAM.scala 148:25:@99620.4]
  wire  _GEN_21; // @[SRAM.scala 148:48:@99622.4]
  reg  regs_22; // @[SRAM.scala 145:20:@99629.4]
  reg [31:0] _RAND_22;
  wire  _T_886; // @[SRAM.scala 148:37:@99630.4]
  wire  _T_887; // @[SRAM.scala 148:25:@99631.4]
  wire  _GEN_22; // @[SRAM.scala 148:48:@99633.4]
  reg  regs_23; // @[SRAM.scala 145:20:@99640.4]
  reg [31:0] _RAND_23;
  wire  _T_895; // @[SRAM.scala 148:37:@99641.4]
  wire  _T_896; // @[SRAM.scala 148:25:@99642.4]
  wire  _GEN_23; // @[SRAM.scala 148:48:@99644.4]
  reg  regs_24; // @[SRAM.scala 145:20:@99651.4]
  reg [31:0] _RAND_24;
  wire  _T_904; // @[SRAM.scala 148:37:@99652.4]
  wire  _T_905; // @[SRAM.scala 148:25:@99653.4]
  wire  _GEN_24; // @[SRAM.scala 148:48:@99655.4]
  reg  regs_25; // @[SRAM.scala 145:20:@99662.4]
  reg [31:0] _RAND_25;
  wire  _T_913; // @[SRAM.scala 148:37:@99663.4]
  wire  _T_914; // @[SRAM.scala 148:25:@99664.4]
  wire  _GEN_25; // @[SRAM.scala 148:48:@99666.4]
  reg  regs_26; // @[SRAM.scala 145:20:@99673.4]
  reg [31:0] _RAND_26;
  wire  _T_922; // @[SRAM.scala 148:37:@99674.4]
  wire  _T_923; // @[SRAM.scala 148:25:@99675.4]
  wire  _GEN_26; // @[SRAM.scala 148:48:@99677.4]
  reg  regs_27; // @[SRAM.scala 145:20:@99684.4]
  reg [31:0] _RAND_27;
  wire  _T_931; // @[SRAM.scala 148:37:@99685.4]
  wire  _T_932; // @[SRAM.scala 148:25:@99686.4]
  wire  _GEN_27; // @[SRAM.scala 148:48:@99688.4]
  reg  regs_28; // @[SRAM.scala 145:20:@99695.4]
  reg [31:0] _RAND_28;
  wire  _T_940; // @[SRAM.scala 148:37:@99696.4]
  wire  _T_941; // @[SRAM.scala 148:25:@99697.4]
  wire  _GEN_28; // @[SRAM.scala 148:48:@99699.4]
  reg  regs_29; // @[SRAM.scala 145:20:@99706.4]
  reg [31:0] _RAND_29;
  wire  _T_949; // @[SRAM.scala 148:37:@99707.4]
  wire  _T_950; // @[SRAM.scala 148:25:@99708.4]
  wire  _GEN_29; // @[SRAM.scala 148:48:@99710.4]
  reg  regs_30; // @[SRAM.scala 145:20:@99717.4]
  reg [31:0] _RAND_30;
  wire  _T_958; // @[SRAM.scala 148:37:@99718.4]
  wire  _T_959; // @[SRAM.scala 148:25:@99719.4]
  wire  _GEN_30; // @[SRAM.scala 148:48:@99721.4]
  reg  regs_31; // @[SRAM.scala 145:20:@99728.4]
  reg [31:0] _RAND_31;
  wire  _T_967; // @[SRAM.scala 148:37:@99729.4]
  wire  _T_968; // @[SRAM.scala 148:25:@99730.4]
  wire  _GEN_31; // @[SRAM.scala 148:48:@99732.4]
  reg  regs_32; // @[SRAM.scala 145:20:@99739.4]
  reg [31:0] _RAND_32;
  wire  _T_976; // @[SRAM.scala 148:37:@99740.4]
  wire  _T_977; // @[SRAM.scala 148:25:@99741.4]
  wire  _GEN_32; // @[SRAM.scala 148:48:@99743.4]
  reg  regs_33; // @[SRAM.scala 145:20:@99750.4]
  reg [31:0] _RAND_33;
  wire  _T_985; // @[SRAM.scala 148:37:@99751.4]
  wire  _T_986; // @[SRAM.scala 148:25:@99752.4]
  wire  _GEN_33; // @[SRAM.scala 148:48:@99754.4]
  reg  regs_34; // @[SRAM.scala 145:20:@99761.4]
  reg [31:0] _RAND_34;
  wire  _T_994; // @[SRAM.scala 148:37:@99762.4]
  wire  _T_995; // @[SRAM.scala 148:25:@99763.4]
  wire  _GEN_34; // @[SRAM.scala 148:48:@99765.4]
  reg  regs_35; // @[SRAM.scala 145:20:@99772.4]
  reg [31:0] _RAND_35;
  wire  _T_1003; // @[SRAM.scala 148:37:@99773.4]
  wire  _T_1004; // @[SRAM.scala 148:25:@99774.4]
  wire  _GEN_35; // @[SRAM.scala 148:48:@99776.4]
  reg  regs_36; // @[SRAM.scala 145:20:@99783.4]
  reg [31:0] _RAND_36;
  wire  _T_1012; // @[SRAM.scala 148:37:@99784.4]
  wire  _T_1013; // @[SRAM.scala 148:25:@99785.4]
  wire  _GEN_36; // @[SRAM.scala 148:48:@99787.4]
  reg  regs_37; // @[SRAM.scala 145:20:@99794.4]
  reg [31:0] _RAND_37;
  wire  _T_1021; // @[SRAM.scala 148:37:@99795.4]
  wire  _T_1022; // @[SRAM.scala 148:25:@99796.4]
  wire  _GEN_37; // @[SRAM.scala 148:48:@99798.4]
  reg  regs_38; // @[SRAM.scala 145:20:@99805.4]
  reg [31:0] _RAND_38;
  wire  _T_1030; // @[SRAM.scala 148:37:@99806.4]
  wire  _T_1031; // @[SRAM.scala 148:25:@99807.4]
  wire  _GEN_38; // @[SRAM.scala 148:48:@99809.4]
  reg  regs_39; // @[SRAM.scala 145:20:@99816.4]
  reg [31:0] _RAND_39;
  wire  _T_1039; // @[SRAM.scala 148:37:@99817.4]
  wire  _T_1040; // @[SRAM.scala 148:25:@99818.4]
  wire  _GEN_39; // @[SRAM.scala 148:48:@99820.4]
  reg  regs_40; // @[SRAM.scala 145:20:@99827.4]
  reg [31:0] _RAND_40;
  wire  _T_1048; // @[SRAM.scala 148:37:@99828.4]
  wire  _T_1049; // @[SRAM.scala 148:25:@99829.4]
  wire  _GEN_40; // @[SRAM.scala 148:48:@99831.4]
  reg  regs_41; // @[SRAM.scala 145:20:@99838.4]
  reg [31:0] _RAND_41;
  wire  _T_1057; // @[SRAM.scala 148:37:@99839.4]
  wire  _T_1058; // @[SRAM.scala 148:25:@99840.4]
  wire  _GEN_41; // @[SRAM.scala 148:48:@99842.4]
  reg  regs_42; // @[SRAM.scala 145:20:@99849.4]
  reg [31:0] _RAND_42;
  wire  _T_1066; // @[SRAM.scala 148:37:@99850.4]
  wire  _T_1067; // @[SRAM.scala 148:25:@99851.4]
  wire  _GEN_42; // @[SRAM.scala 148:48:@99853.4]
  reg  regs_43; // @[SRAM.scala 145:20:@99860.4]
  reg [31:0] _RAND_43;
  wire  _T_1075; // @[SRAM.scala 148:37:@99861.4]
  wire  _T_1076; // @[SRAM.scala 148:25:@99862.4]
  wire  _GEN_43; // @[SRAM.scala 148:48:@99864.4]
  reg  regs_44; // @[SRAM.scala 145:20:@99871.4]
  reg [31:0] _RAND_44;
  wire  _T_1084; // @[SRAM.scala 148:37:@99872.4]
  wire  _T_1085; // @[SRAM.scala 148:25:@99873.4]
  wire  _GEN_44; // @[SRAM.scala 148:48:@99875.4]
  reg  regs_45; // @[SRAM.scala 145:20:@99882.4]
  reg [31:0] _RAND_45;
  wire  _T_1093; // @[SRAM.scala 148:37:@99883.4]
  wire  _T_1094; // @[SRAM.scala 148:25:@99884.4]
  wire  _GEN_45; // @[SRAM.scala 148:48:@99886.4]
  reg  regs_46; // @[SRAM.scala 145:20:@99893.4]
  reg [31:0] _RAND_46;
  wire  _T_1102; // @[SRAM.scala 148:37:@99894.4]
  wire  _T_1103; // @[SRAM.scala 148:25:@99895.4]
  wire  _GEN_46; // @[SRAM.scala 148:48:@99897.4]
  reg  regs_47; // @[SRAM.scala 145:20:@99904.4]
  reg [31:0] _RAND_47;
  wire  _T_1111; // @[SRAM.scala 148:37:@99905.4]
  wire  _T_1112; // @[SRAM.scala 148:25:@99906.4]
  wire  _GEN_47; // @[SRAM.scala 148:48:@99908.4]
  reg  regs_48; // @[SRAM.scala 145:20:@99915.4]
  reg [31:0] _RAND_48;
  wire  _T_1120; // @[SRAM.scala 148:37:@99916.4]
  wire  _T_1121; // @[SRAM.scala 148:25:@99917.4]
  wire  _GEN_48; // @[SRAM.scala 148:48:@99919.4]
  reg  regs_49; // @[SRAM.scala 145:20:@99926.4]
  reg [31:0] _RAND_49;
  wire  _T_1129; // @[SRAM.scala 148:37:@99927.4]
  wire  _T_1130; // @[SRAM.scala 148:25:@99928.4]
  wire  _GEN_49; // @[SRAM.scala 148:48:@99930.4]
  reg  regs_50; // @[SRAM.scala 145:20:@99937.4]
  reg [31:0] _RAND_50;
  wire  _T_1138; // @[SRAM.scala 148:37:@99938.4]
  wire  _T_1139; // @[SRAM.scala 148:25:@99939.4]
  wire  _GEN_50; // @[SRAM.scala 148:48:@99941.4]
  reg  regs_51; // @[SRAM.scala 145:20:@99948.4]
  reg [31:0] _RAND_51;
  wire  _T_1147; // @[SRAM.scala 148:37:@99949.4]
  wire  _T_1148; // @[SRAM.scala 148:25:@99950.4]
  wire  _GEN_51; // @[SRAM.scala 148:48:@99952.4]
  reg  regs_52; // @[SRAM.scala 145:20:@99959.4]
  reg [31:0] _RAND_52;
  wire  _T_1156; // @[SRAM.scala 148:37:@99960.4]
  wire  _T_1157; // @[SRAM.scala 148:25:@99961.4]
  wire  _GEN_52; // @[SRAM.scala 148:48:@99963.4]
  reg  regs_53; // @[SRAM.scala 145:20:@99970.4]
  reg [31:0] _RAND_53;
  wire  _T_1165; // @[SRAM.scala 148:37:@99971.4]
  wire  _T_1166; // @[SRAM.scala 148:25:@99972.4]
  wire  _GEN_53; // @[SRAM.scala 148:48:@99974.4]
  reg  regs_54; // @[SRAM.scala 145:20:@99981.4]
  reg [31:0] _RAND_54;
  wire  _T_1174; // @[SRAM.scala 148:37:@99982.4]
  wire  _T_1175; // @[SRAM.scala 148:25:@99983.4]
  wire  _GEN_54; // @[SRAM.scala 148:48:@99985.4]
  reg  regs_55; // @[SRAM.scala 145:20:@99992.4]
  reg [31:0] _RAND_55;
  wire  _T_1183; // @[SRAM.scala 148:37:@99993.4]
  wire  _T_1184; // @[SRAM.scala 148:25:@99994.4]
  wire  _GEN_55; // @[SRAM.scala 148:48:@99996.4]
  reg  regs_56; // @[SRAM.scala 145:20:@100003.4]
  reg [31:0] _RAND_56;
  wire  _T_1192; // @[SRAM.scala 148:37:@100004.4]
  wire  _T_1193; // @[SRAM.scala 148:25:@100005.4]
  wire  _GEN_56; // @[SRAM.scala 148:48:@100007.4]
  reg  regs_57; // @[SRAM.scala 145:20:@100014.4]
  reg [31:0] _RAND_57;
  wire  _T_1201; // @[SRAM.scala 148:37:@100015.4]
  wire  _T_1202; // @[SRAM.scala 148:25:@100016.4]
  wire  _GEN_57; // @[SRAM.scala 148:48:@100018.4]
  reg  regs_58; // @[SRAM.scala 145:20:@100025.4]
  reg [31:0] _RAND_58;
  wire  _T_1210; // @[SRAM.scala 148:37:@100026.4]
  wire  _T_1211; // @[SRAM.scala 148:25:@100027.4]
  wire  _GEN_58; // @[SRAM.scala 148:48:@100029.4]
  reg  regs_59; // @[SRAM.scala 145:20:@100036.4]
  reg [31:0] _RAND_59;
  wire  _T_1219; // @[SRAM.scala 148:37:@100037.4]
  wire  _T_1220; // @[SRAM.scala 148:25:@100038.4]
  wire  _GEN_59; // @[SRAM.scala 148:48:@100040.4]
  reg  regs_60; // @[SRAM.scala 145:20:@100047.4]
  reg [31:0] _RAND_60;
  wire  _T_1228; // @[SRAM.scala 148:37:@100048.4]
  wire  _T_1229; // @[SRAM.scala 148:25:@100049.4]
  wire  _GEN_60; // @[SRAM.scala 148:48:@100051.4]
  reg  regs_61; // @[SRAM.scala 145:20:@100058.4]
  reg [31:0] _RAND_61;
  wire  _T_1237; // @[SRAM.scala 148:37:@100059.4]
  wire  _T_1238; // @[SRAM.scala 148:25:@100060.4]
  wire  _GEN_61; // @[SRAM.scala 148:48:@100062.4]
  reg  regs_62; // @[SRAM.scala 145:20:@100069.4]
  reg [31:0] _RAND_62;
  wire  _T_1246; // @[SRAM.scala 148:37:@100070.4]
  wire  _T_1247; // @[SRAM.scala 148:25:@100071.4]
  wire  _GEN_62; // @[SRAM.scala 148:48:@100073.4]
  reg  regs_63; // @[SRAM.scala 145:20:@100080.4]
  reg [31:0] _RAND_63;
  wire  _T_1255; // @[SRAM.scala 148:37:@100081.4]
  wire  _T_1256; // @[SRAM.scala 148:25:@100082.4]
  wire  _GEN_63; // @[SRAM.scala 148:48:@100084.4]
  wire  _GEN_65; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_66; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_67; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_68; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_69; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_70; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_71; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_72; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_73; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_74; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_75; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_76; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_77; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_78; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_79; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_80; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_81; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_82; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_83; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_84; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_85; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_86; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_87; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_88; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_89; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_90; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_91; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_92; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_93; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_94; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_95; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_96; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_97; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_98; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_99; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_100; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_101; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_102; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_103; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_104; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_105; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_106; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_107; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_108; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_109; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_110; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_111; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_112; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_113; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_114; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_115; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_116; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_117; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_118; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_119; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_120; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_121; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_122; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_123; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_124; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_125; // @[SRAM.scala 155:12:@100154.4]
  wire  _GEN_126; // @[SRAM.scala 155:12:@100154.4]
  assign _T_688 = io_waddr == 6'h0; // @[SRAM.scala 148:37:@99388.4]
  assign _T_689 = io_wen & _T_688; // @[SRAM.scala 148:25:@99389.4]
  assign _GEN_0 = _T_689 ? 1'h1 : regs_0; // @[SRAM.scala 148:48:@99391.4]
  assign _T_697 = io_waddr == 6'h1; // @[SRAM.scala 148:37:@99399.4]
  assign _T_698 = io_wen & _T_697; // @[SRAM.scala 148:25:@99400.4]
  assign _GEN_1 = _T_698 ? 1'h1 : regs_1; // @[SRAM.scala 148:48:@99402.4]
  assign _T_706 = io_waddr == 6'h2; // @[SRAM.scala 148:37:@99410.4]
  assign _T_707 = io_wen & _T_706; // @[SRAM.scala 148:25:@99411.4]
  assign _GEN_2 = _T_707 ? 1'h1 : regs_2; // @[SRAM.scala 148:48:@99413.4]
  assign _T_715 = io_waddr == 6'h3; // @[SRAM.scala 148:37:@99421.4]
  assign _T_716 = io_wen & _T_715; // @[SRAM.scala 148:25:@99422.4]
  assign _GEN_3 = _T_716 ? 1'h1 : regs_3; // @[SRAM.scala 148:48:@99424.4]
  assign _T_724 = io_waddr == 6'h4; // @[SRAM.scala 148:37:@99432.4]
  assign _T_725 = io_wen & _T_724; // @[SRAM.scala 148:25:@99433.4]
  assign _GEN_4 = _T_725 ? 1'h1 : regs_4; // @[SRAM.scala 148:48:@99435.4]
  assign _T_733 = io_waddr == 6'h5; // @[SRAM.scala 148:37:@99443.4]
  assign _T_734 = io_wen & _T_733; // @[SRAM.scala 148:25:@99444.4]
  assign _GEN_5 = _T_734 ? 1'h1 : regs_5; // @[SRAM.scala 148:48:@99446.4]
  assign _T_742 = io_waddr == 6'h6; // @[SRAM.scala 148:37:@99454.4]
  assign _T_743 = io_wen & _T_742; // @[SRAM.scala 148:25:@99455.4]
  assign _GEN_6 = _T_743 ? 1'h1 : regs_6; // @[SRAM.scala 148:48:@99457.4]
  assign _T_751 = io_waddr == 6'h7; // @[SRAM.scala 148:37:@99465.4]
  assign _T_752 = io_wen & _T_751; // @[SRAM.scala 148:25:@99466.4]
  assign _GEN_7 = _T_752 ? 1'h1 : regs_7; // @[SRAM.scala 148:48:@99468.4]
  assign _T_760 = io_waddr == 6'h8; // @[SRAM.scala 148:37:@99476.4]
  assign _T_761 = io_wen & _T_760; // @[SRAM.scala 148:25:@99477.4]
  assign _GEN_8 = _T_761 ? 1'h1 : regs_8; // @[SRAM.scala 148:48:@99479.4]
  assign _T_769 = io_waddr == 6'h9; // @[SRAM.scala 148:37:@99487.4]
  assign _T_770 = io_wen & _T_769; // @[SRAM.scala 148:25:@99488.4]
  assign _GEN_9 = _T_770 ? 1'h1 : regs_9; // @[SRAM.scala 148:48:@99490.4]
  assign _T_778 = io_waddr == 6'ha; // @[SRAM.scala 148:37:@99498.4]
  assign _T_779 = io_wen & _T_778; // @[SRAM.scala 148:25:@99499.4]
  assign _GEN_10 = _T_779 ? 1'h1 : regs_10; // @[SRAM.scala 148:48:@99501.4]
  assign _T_787 = io_waddr == 6'hb; // @[SRAM.scala 148:37:@99509.4]
  assign _T_788 = io_wen & _T_787; // @[SRAM.scala 148:25:@99510.4]
  assign _GEN_11 = _T_788 ? 1'h1 : regs_11; // @[SRAM.scala 148:48:@99512.4]
  assign _T_796 = io_waddr == 6'hc; // @[SRAM.scala 148:37:@99520.4]
  assign _T_797 = io_wen & _T_796; // @[SRAM.scala 148:25:@99521.4]
  assign _GEN_12 = _T_797 ? 1'h1 : regs_12; // @[SRAM.scala 148:48:@99523.4]
  assign _T_805 = io_waddr == 6'hd; // @[SRAM.scala 148:37:@99531.4]
  assign _T_806 = io_wen & _T_805; // @[SRAM.scala 148:25:@99532.4]
  assign _GEN_13 = _T_806 ? 1'h1 : regs_13; // @[SRAM.scala 148:48:@99534.4]
  assign _T_814 = io_waddr == 6'he; // @[SRAM.scala 148:37:@99542.4]
  assign _T_815 = io_wen & _T_814; // @[SRAM.scala 148:25:@99543.4]
  assign _GEN_14 = _T_815 ? 1'h1 : regs_14; // @[SRAM.scala 148:48:@99545.4]
  assign _T_823 = io_waddr == 6'hf; // @[SRAM.scala 148:37:@99553.4]
  assign _T_824 = io_wen & _T_823; // @[SRAM.scala 148:25:@99554.4]
  assign _GEN_15 = _T_824 ? 1'h1 : regs_15; // @[SRAM.scala 148:48:@99556.4]
  assign _T_832 = io_waddr == 6'h10; // @[SRAM.scala 148:37:@99564.4]
  assign _T_833 = io_wen & _T_832; // @[SRAM.scala 148:25:@99565.4]
  assign _GEN_16 = _T_833 ? 1'h1 : regs_16; // @[SRAM.scala 148:48:@99567.4]
  assign _T_841 = io_waddr == 6'h11; // @[SRAM.scala 148:37:@99575.4]
  assign _T_842 = io_wen & _T_841; // @[SRAM.scala 148:25:@99576.4]
  assign _GEN_17 = _T_842 ? 1'h1 : regs_17; // @[SRAM.scala 148:48:@99578.4]
  assign _T_850 = io_waddr == 6'h12; // @[SRAM.scala 148:37:@99586.4]
  assign _T_851 = io_wen & _T_850; // @[SRAM.scala 148:25:@99587.4]
  assign _GEN_18 = _T_851 ? 1'h1 : regs_18; // @[SRAM.scala 148:48:@99589.4]
  assign _T_859 = io_waddr == 6'h13; // @[SRAM.scala 148:37:@99597.4]
  assign _T_860 = io_wen & _T_859; // @[SRAM.scala 148:25:@99598.4]
  assign _GEN_19 = _T_860 ? 1'h1 : regs_19; // @[SRAM.scala 148:48:@99600.4]
  assign _T_868 = io_waddr == 6'h14; // @[SRAM.scala 148:37:@99608.4]
  assign _T_869 = io_wen & _T_868; // @[SRAM.scala 148:25:@99609.4]
  assign _GEN_20 = _T_869 ? 1'h1 : regs_20; // @[SRAM.scala 148:48:@99611.4]
  assign _T_877 = io_waddr == 6'h15; // @[SRAM.scala 148:37:@99619.4]
  assign _T_878 = io_wen & _T_877; // @[SRAM.scala 148:25:@99620.4]
  assign _GEN_21 = _T_878 ? 1'h1 : regs_21; // @[SRAM.scala 148:48:@99622.4]
  assign _T_886 = io_waddr == 6'h16; // @[SRAM.scala 148:37:@99630.4]
  assign _T_887 = io_wen & _T_886; // @[SRAM.scala 148:25:@99631.4]
  assign _GEN_22 = _T_887 ? 1'h1 : regs_22; // @[SRAM.scala 148:48:@99633.4]
  assign _T_895 = io_waddr == 6'h17; // @[SRAM.scala 148:37:@99641.4]
  assign _T_896 = io_wen & _T_895; // @[SRAM.scala 148:25:@99642.4]
  assign _GEN_23 = _T_896 ? 1'h1 : regs_23; // @[SRAM.scala 148:48:@99644.4]
  assign _T_904 = io_waddr == 6'h18; // @[SRAM.scala 148:37:@99652.4]
  assign _T_905 = io_wen & _T_904; // @[SRAM.scala 148:25:@99653.4]
  assign _GEN_24 = _T_905 ? 1'h1 : regs_24; // @[SRAM.scala 148:48:@99655.4]
  assign _T_913 = io_waddr == 6'h19; // @[SRAM.scala 148:37:@99663.4]
  assign _T_914 = io_wen & _T_913; // @[SRAM.scala 148:25:@99664.4]
  assign _GEN_25 = _T_914 ? 1'h1 : regs_25; // @[SRAM.scala 148:48:@99666.4]
  assign _T_922 = io_waddr == 6'h1a; // @[SRAM.scala 148:37:@99674.4]
  assign _T_923 = io_wen & _T_922; // @[SRAM.scala 148:25:@99675.4]
  assign _GEN_26 = _T_923 ? 1'h1 : regs_26; // @[SRAM.scala 148:48:@99677.4]
  assign _T_931 = io_waddr == 6'h1b; // @[SRAM.scala 148:37:@99685.4]
  assign _T_932 = io_wen & _T_931; // @[SRAM.scala 148:25:@99686.4]
  assign _GEN_27 = _T_932 ? 1'h1 : regs_27; // @[SRAM.scala 148:48:@99688.4]
  assign _T_940 = io_waddr == 6'h1c; // @[SRAM.scala 148:37:@99696.4]
  assign _T_941 = io_wen & _T_940; // @[SRAM.scala 148:25:@99697.4]
  assign _GEN_28 = _T_941 ? 1'h1 : regs_28; // @[SRAM.scala 148:48:@99699.4]
  assign _T_949 = io_waddr == 6'h1d; // @[SRAM.scala 148:37:@99707.4]
  assign _T_950 = io_wen & _T_949; // @[SRAM.scala 148:25:@99708.4]
  assign _GEN_29 = _T_950 ? 1'h1 : regs_29; // @[SRAM.scala 148:48:@99710.4]
  assign _T_958 = io_waddr == 6'h1e; // @[SRAM.scala 148:37:@99718.4]
  assign _T_959 = io_wen & _T_958; // @[SRAM.scala 148:25:@99719.4]
  assign _GEN_30 = _T_959 ? 1'h1 : regs_30; // @[SRAM.scala 148:48:@99721.4]
  assign _T_967 = io_waddr == 6'h1f; // @[SRAM.scala 148:37:@99729.4]
  assign _T_968 = io_wen & _T_967; // @[SRAM.scala 148:25:@99730.4]
  assign _GEN_31 = _T_968 ? 1'h1 : regs_31; // @[SRAM.scala 148:48:@99732.4]
  assign _T_976 = io_waddr == 6'h20; // @[SRAM.scala 148:37:@99740.4]
  assign _T_977 = io_wen & _T_976; // @[SRAM.scala 148:25:@99741.4]
  assign _GEN_32 = _T_977 ? 1'h1 : regs_32; // @[SRAM.scala 148:48:@99743.4]
  assign _T_985 = io_waddr == 6'h21; // @[SRAM.scala 148:37:@99751.4]
  assign _T_986 = io_wen & _T_985; // @[SRAM.scala 148:25:@99752.4]
  assign _GEN_33 = _T_986 ? 1'h1 : regs_33; // @[SRAM.scala 148:48:@99754.4]
  assign _T_994 = io_waddr == 6'h22; // @[SRAM.scala 148:37:@99762.4]
  assign _T_995 = io_wen & _T_994; // @[SRAM.scala 148:25:@99763.4]
  assign _GEN_34 = _T_995 ? 1'h1 : regs_34; // @[SRAM.scala 148:48:@99765.4]
  assign _T_1003 = io_waddr == 6'h23; // @[SRAM.scala 148:37:@99773.4]
  assign _T_1004 = io_wen & _T_1003; // @[SRAM.scala 148:25:@99774.4]
  assign _GEN_35 = _T_1004 ? 1'h1 : regs_35; // @[SRAM.scala 148:48:@99776.4]
  assign _T_1012 = io_waddr == 6'h24; // @[SRAM.scala 148:37:@99784.4]
  assign _T_1013 = io_wen & _T_1012; // @[SRAM.scala 148:25:@99785.4]
  assign _GEN_36 = _T_1013 ? 1'h1 : regs_36; // @[SRAM.scala 148:48:@99787.4]
  assign _T_1021 = io_waddr == 6'h25; // @[SRAM.scala 148:37:@99795.4]
  assign _T_1022 = io_wen & _T_1021; // @[SRAM.scala 148:25:@99796.4]
  assign _GEN_37 = _T_1022 ? 1'h1 : regs_37; // @[SRAM.scala 148:48:@99798.4]
  assign _T_1030 = io_waddr == 6'h26; // @[SRAM.scala 148:37:@99806.4]
  assign _T_1031 = io_wen & _T_1030; // @[SRAM.scala 148:25:@99807.4]
  assign _GEN_38 = _T_1031 ? 1'h1 : regs_38; // @[SRAM.scala 148:48:@99809.4]
  assign _T_1039 = io_waddr == 6'h27; // @[SRAM.scala 148:37:@99817.4]
  assign _T_1040 = io_wen & _T_1039; // @[SRAM.scala 148:25:@99818.4]
  assign _GEN_39 = _T_1040 ? 1'h1 : regs_39; // @[SRAM.scala 148:48:@99820.4]
  assign _T_1048 = io_waddr == 6'h28; // @[SRAM.scala 148:37:@99828.4]
  assign _T_1049 = io_wen & _T_1048; // @[SRAM.scala 148:25:@99829.4]
  assign _GEN_40 = _T_1049 ? 1'h1 : regs_40; // @[SRAM.scala 148:48:@99831.4]
  assign _T_1057 = io_waddr == 6'h29; // @[SRAM.scala 148:37:@99839.4]
  assign _T_1058 = io_wen & _T_1057; // @[SRAM.scala 148:25:@99840.4]
  assign _GEN_41 = _T_1058 ? 1'h1 : regs_41; // @[SRAM.scala 148:48:@99842.4]
  assign _T_1066 = io_waddr == 6'h2a; // @[SRAM.scala 148:37:@99850.4]
  assign _T_1067 = io_wen & _T_1066; // @[SRAM.scala 148:25:@99851.4]
  assign _GEN_42 = _T_1067 ? 1'h1 : regs_42; // @[SRAM.scala 148:48:@99853.4]
  assign _T_1075 = io_waddr == 6'h2b; // @[SRAM.scala 148:37:@99861.4]
  assign _T_1076 = io_wen & _T_1075; // @[SRAM.scala 148:25:@99862.4]
  assign _GEN_43 = _T_1076 ? 1'h1 : regs_43; // @[SRAM.scala 148:48:@99864.4]
  assign _T_1084 = io_waddr == 6'h2c; // @[SRAM.scala 148:37:@99872.4]
  assign _T_1085 = io_wen & _T_1084; // @[SRAM.scala 148:25:@99873.4]
  assign _GEN_44 = _T_1085 ? 1'h1 : regs_44; // @[SRAM.scala 148:48:@99875.4]
  assign _T_1093 = io_waddr == 6'h2d; // @[SRAM.scala 148:37:@99883.4]
  assign _T_1094 = io_wen & _T_1093; // @[SRAM.scala 148:25:@99884.4]
  assign _GEN_45 = _T_1094 ? 1'h1 : regs_45; // @[SRAM.scala 148:48:@99886.4]
  assign _T_1102 = io_waddr == 6'h2e; // @[SRAM.scala 148:37:@99894.4]
  assign _T_1103 = io_wen & _T_1102; // @[SRAM.scala 148:25:@99895.4]
  assign _GEN_46 = _T_1103 ? 1'h1 : regs_46; // @[SRAM.scala 148:48:@99897.4]
  assign _T_1111 = io_waddr == 6'h2f; // @[SRAM.scala 148:37:@99905.4]
  assign _T_1112 = io_wen & _T_1111; // @[SRAM.scala 148:25:@99906.4]
  assign _GEN_47 = _T_1112 ? 1'h1 : regs_47; // @[SRAM.scala 148:48:@99908.4]
  assign _T_1120 = io_waddr == 6'h30; // @[SRAM.scala 148:37:@99916.4]
  assign _T_1121 = io_wen & _T_1120; // @[SRAM.scala 148:25:@99917.4]
  assign _GEN_48 = _T_1121 ? 1'h1 : regs_48; // @[SRAM.scala 148:48:@99919.4]
  assign _T_1129 = io_waddr == 6'h31; // @[SRAM.scala 148:37:@99927.4]
  assign _T_1130 = io_wen & _T_1129; // @[SRAM.scala 148:25:@99928.4]
  assign _GEN_49 = _T_1130 ? 1'h1 : regs_49; // @[SRAM.scala 148:48:@99930.4]
  assign _T_1138 = io_waddr == 6'h32; // @[SRAM.scala 148:37:@99938.4]
  assign _T_1139 = io_wen & _T_1138; // @[SRAM.scala 148:25:@99939.4]
  assign _GEN_50 = _T_1139 ? 1'h1 : regs_50; // @[SRAM.scala 148:48:@99941.4]
  assign _T_1147 = io_waddr == 6'h33; // @[SRAM.scala 148:37:@99949.4]
  assign _T_1148 = io_wen & _T_1147; // @[SRAM.scala 148:25:@99950.4]
  assign _GEN_51 = _T_1148 ? 1'h1 : regs_51; // @[SRAM.scala 148:48:@99952.4]
  assign _T_1156 = io_waddr == 6'h34; // @[SRAM.scala 148:37:@99960.4]
  assign _T_1157 = io_wen & _T_1156; // @[SRAM.scala 148:25:@99961.4]
  assign _GEN_52 = _T_1157 ? 1'h1 : regs_52; // @[SRAM.scala 148:48:@99963.4]
  assign _T_1165 = io_waddr == 6'h35; // @[SRAM.scala 148:37:@99971.4]
  assign _T_1166 = io_wen & _T_1165; // @[SRAM.scala 148:25:@99972.4]
  assign _GEN_53 = _T_1166 ? 1'h1 : regs_53; // @[SRAM.scala 148:48:@99974.4]
  assign _T_1174 = io_waddr == 6'h36; // @[SRAM.scala 148:37:@99982.4]
  assign _T_1175 = io_wen & _T_1174; // @[SRAM.scala 148:25:@99983.4]
  assign _GEN_54 = _T_1175 ? 1'h1 : regs_54; // @[SRAM.scala 148:48:@99985.4]
  assign _T_1183 = io_waddr == 6'h37; // @[SRAM.scala 148:37:@99993.4]
  assign _T_1184 = io_wen & _T_1183; // @[SRAM.scala 148:25:@99994.4]
  assign _GEN_55 = _T_1184 ? 1'h1 : regs_55; // @[SRAM.scala 148:48:@99996.4]
  assign _T_1192 = io_waddr == 6'h38; // @[SRAM.scala 148:37:@100004.4]
  assign _T_1193 = io_wen & _T_1192; // @[SRAM.scala 148:25:@100005.4]
  assign _GEN_56 = _T_1193 ? 1'h1 : regs_56; // @[SRAM.scala 148:48:@100007.4]
  assign _T_1201 = io_waddr == 6'h39; // @[SRAM.scala 148:37:@100015.4]
  assign _T_1202 = io_wen & _T_1201; // @[SRAM.scala 148:25:@100016.4]
  assign _GEN_57 = _T_1202 ? 1'h1 : regs_57; // @[SRAM.scala 148:48:@100018.4]
  assign _T_1210 = io_waddr == 6'h3a; // @[SRAM.scala 148:37:@100026.4]
  assign _T_1211 = io_wen & _T_1210; // @[SRAM.scala 148:25:@100027.4]
  assign _GEN_58 = _T_1211 ? 1'h1 : regs_58; // @[SRAM.scala 148:48:@100029.4]
  assign _T_1219 = io_waddr == 6'h3b; // @[SRAM.scala 148:37:@100037.4]
  assign _T_1220 = io_wen & _T_1219; // @[SRAM.scala 148:25:@100038.4]
  assign _GEN_59 = _T_1220 ? 1'h1 : regs_59; // @[SRAM.scala 148:48:@100040.4]
  assign _T_1228 = io_waddr == 6'h3c; // @[SRAM.scala 148:37:@100048.4]
  assign _T_1229 = io_wen & _T_1228; // @[SRAM.scala 148:25:@100049.4]
  assign _GEN_60 = _T_1229 ? 1'h1 : regs_60; // @[SRAM.scala 148:48:@100051.4]
  assign _T_1237 = io_waddr == 6'h3d; // @[SRAM.scala 148:37:@100059.4]
  assign _T_1238 = io_wen & _T_1237; // @[SRAM.scala 148:25:@100060.4]
  assign _GEN_61 = _T_1238 ? 1'h1 : regs_61; // @[SRAM.scala 148:48:@100062.4]
  assign _T_1246 = io_waddr == 6'h3e; // @[SRAM.scala 148:37:@100070.4]
  assign _T_1247 = io_wen & _T_1246; // @[SRAM.scala 148:25:@100071.4]
  assign _GEN_62 = _T_1247 ? 1'h1 : regs_62; // @[SRAM.scala 148:48:@100073.4]
  assign _T_1255 = io_waddr == 6'h3f; // @[SRAM.scala 148:37:@100081.4]
  assign _T_1256 = io_wen & _T_1255; // @[SRAM.scala 148:25:@100082.4]
  assign _GEN_63 = _T_1256 ? 1'h1 : regs_63; // @[SRAM.scala 148:48:@100084.4]
  assign _GEN_65 = 6'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_66 = 6'h2 == io_raddr ? regs_2 : _GEN_65; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_67 = 6'h3 == io_raddr ? regs_3 : _GEN_66; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_68 = 6'h4 == io_raddr ? regs_4 : _GEN_67; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_69 = 6'h5 == io_raddr ? regs_5 : _GEN_68; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_70 = 6'h6 == io_raddr ? regs_6 : _GEN_69; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_71 = 6'h7 == io_raddr ? regs_7 : _GEN_70; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_72 = 6'h8 == io_raddr ? regs_8 : _GEN_71; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_73 = 6'h9 == io_raddr ? regs_9 : _GEN_72; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_74 = 6'ha == io_raddr ? regs_10 : _GEN_73; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_75 = 6'hb == io_raddr ? regs_11 : _GEN_74; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_76 = 6'hc == io_raddr ? regs_12 : _GEN_75; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_77 = 6'hd == io_raddr ? regs_13 : _GEN_76; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_78 = 6'he == io_raddr ? regs_14 : _GEN_77; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_79 = 6'hf == io_raddr ? regs_15 : _GEN_78; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_80 = 6'h10 == io_raddr ? regs_16 : _GEN_79; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_81 = 6'h11 == io_raddr ? regs_17 : _GEN_80; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_82 = 6'h12 == io_raddr ? regs_18 : _GEN_81; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_83 = 6'h13 == io_raddr ? regs_19 : _GEN_82; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_84 = 6'h14 == io_raddr ? regs_20 : _GEN_83; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_85 = 6'h15 == io_raddr ? regs_21 : _GEN_84; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_86 = 6'h16 == io_raddr ? regs_22 : _GEN_85; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_87 = 6'h17 == io_raddr ? regs_23 : _GEN_86; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_88 = 6'h18 == io_raddr ? regs_24 : _GEN_87; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_89 = 6'h19 == io_raddr ? regs_25 : _GEN_88; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_90 = 6'h1a == io_raddr ? regs_26 : _GEN_89; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_91 = 6'h1b == io_raddr ? regs_27 : _GEN_90; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_92 = 6'h1c == io_raddr ? regs_28 : _GEN_91; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_93 = 6'h1d == io_raddr ? regs_29 : _GEN_92; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_94 = 6'h1e == io_raddr ? regs_30 : _GEN_93; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_95 = 6'h1f == io_raddr ? regs_31 : _GEN_94; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_96 = 6'h20 == io_raddr ? regs_32 : _GEN_95; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_97 = 6'h21 == io_raddr ? regs_33 : _GEN_96; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_98 = 6'h22 == io_raddr ? regs_34 : _GEN_97; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_99 = 6'h23 == io_raddr ? regs_35 : _GEN_98; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_100 = 6'h24 == io_raddr ? regs_36 : _GEN_99; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_101 = 6'h25 == io_raddr ? regs_37 : _GEN_100; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_102 = 6'h26 == io_raddr ? regs_38 : _GEN_101; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_103 = 6'h27 == io_raddr ? regs_39 : _GEN_102; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_104 = 6'h28 == io_raddr ? regs_40 : _GEN_103; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_105 = 6'h29 == io_raddr ? regs_41 : _GEN_104; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_106 = 6'h2a == io_raddr ? regs_42 : _GEN_105; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_107 = 6'h2b == io_raddr ? regs_43 : _GEN_106; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_108 = 6'h2c == io_raddr ? regs_44 : _GEN_107; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_109 = 6'h2d == io_raddr ? regs_45 : _GEN_108; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_110 = 6'h2e == io_raddr ? regs_46 : _GEN_109; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_111 = 6'h2f == io_raddr ? regs_47 : _GEN_110; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_112 = 6'h30 == io_raddr ? regs_48 : _GEN_111; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_113 = 6'h31 == io_raddr ? regs_49 : _GEN_112; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_114 = 6'h32 == io_raddr ? regs_50 : _GEN_113; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_115 = 6'h33 == io_raddr ? regs_51 : _GEN_114; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_116 = 6'h34 == io_raddr ? regs_52 : _GEN_115; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_117 = 6'h35 == io_raddr ? regs_53 : _GEN_116; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_118 = 6'h36 == io_raddr ? regs_54 : _GEN_117; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_119 = 6'h37 == io_raddr ? regs_55 : _GEN_118; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_120 = 6'h38 == io_raddr ? regs_56 : _GEN_119; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_121 = 6'h39 == io_raddr ? regs_57 : _GEN_120; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_122 = 6'h3a == io_raddr ? regs_58 : _GEN_121; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_123 = 6'h3b == io_raddr ? regs_59 : _GEN_122; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_124 = 6'h3c == io_raddr ? regs_60 : _GEN_123; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_125 = 6'h3d == io_raddr ? regs_61 : _GEN_124; // @[SRAM.scala 155:12:@100154.4]
  assign _GEN_126 = 6'h3e == io_raddr ? regs_62 : _GEN_125; // @[SRAM.scala 155:12:@100154.4]
  assign io_rdata = 6'h3f == io_raddr ? regs_63 : _GEN_126; // @[SRAM.scala 155:12:@100154.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_689) begin
        regs_0 <= 1'h1;
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_698) begin
        regs_1 <= 1'h1;
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_707) begin
        regs_2 <= 1'h1;
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_716) begin
        regs_3 <= 1'h1;
      end
    end
    if (reset) begin
      regs_4 <= 1'h0;
    end else begin
      if (_T_725) begin
        regs_4 <= 1'h1;
      end
    end
    if (reset) begin
      regs_5 <= 1'h0;
    end else begin
      if (_T_734) begin
        regs_5 <= 1'h1;
      end
    end
    if (reset) begin
      regs_6 <= 1'h0;
    end else begin
      if (_T_743) begin
        regs_6 <= 1'h1;
      end
    end
    if (reset) begin
      regs_7 <= 1'h0;
    end else begin
      if (_T_752) begin
        regs_7 <= 1'h1;
      end
    end
    if (reset) begin
      regs_8 <= 1'h0;
    end else begin
      if (_T_761) begin
        regs_8 <= 1'h1;
      end
    end
    if (reset) begin
      regs_9 <= 1'h0;
    end else begin
      if (_T_770) begin
        regs_9 <= 1'h1;
      end
    end
    if (reset) begin
      regs_10 <= 1'h0;
    end else begin
      if (_T_779) begin
        regs_10 <= 1'h1;
      end
    end
    if (reset) begin
      regs_11 <= 1'h0;
    end else begin
      if (_T_788) begin
        regs_11 <= 1'h1;
      end
    end
    if (reset) begin
      regs_12 <= 1'h0;
    end else begin
      if (_T_797) begin
        regs_12 <= 1'h1;
      end
    end
    if (reset) begin
      regs_13 <= 1'h0;
    end else begin
      if (_T_806) begin
        regs_13 <= 1'h1;
      end
    end
    if (reset) begin
      regs_14 <= 1'h0;
    end else begin
      if (_T_815) begin
        regs_14 <= 1'h1;
      end
    end
    if (reset) begin
      regs_15 <= 1'h0;
    end else begin
      if (_T_824) begin
        regs_15 <= 1'h1;
      end
    end
    if (reset) begin
      regs_16 <= 1'h0;
    end else begin
      if (_T_833) begin
        regs_16 <= 1'h1;
      end
    end
    if (reset) begin
      regs_17 <= 1'h0;
    end else begin
      if (_T_842) begin
        regs_17 <= 1'h1;
      end
    end
    if (reset) begin
      regs_18 <= 1'h0;
    end else begin
      if (_T_851) begin
        regs_18 <= 1'h1;
      end
    end
    if (reset) begin
      regs_19 <= 1'h0;
    end else begin
      if (_T_860) begin
        regs_19 <= 1'h1;
      end
    end
    if (reset) begin
      regs_20 <= 1'h0;
    end else begin
      if (_T_869) begin
        regs_20 <= 1'h1;
      end
    end
    if (reset) begin
      regs_21 <= 1'h0;
    end else begin
      if (_T_878) begin
        regs_21 <= 1'h1;
      end
    end
    if (reset) begin
      regs_22 <= 1'h0;
    end else begin
      if (_T_887) begin
        regs_22 <= 1'h1;
      end
    end
    if (reset) begin
      regs_23 <= 1'h0;
    end else begin
      if (_T_896) begin
        regs_23 <= 1'h1;
      end
    end
    if (reset) begin
      regs_24 <= 1'h0;
    end else begin
      if (_T_905) begin
        regs_24 <= 1'h1;
      end
    end
    if (reset) begin
      regs_25 <= 1'h0;
    end else begin
      if (_T_914) begin
        regs_25 <= 1'h1;
      end
    end
    if (reset) begin
      regs_26 <= 1'h0;
    end else begin
      if (_T_923) begin
        regs_26 <= 1'h1;
      end
    end
    if (reset) begin
      regs_27 <= 1'h0;
    end else begin
      if (_T_932) begin
        regs_27 <= 1'h1;
      end
    end
    if (reset) begin
      regs_28 <= 1'h0;
    end else begin
      if (_T_941) begin
        regs_28 <= 1'h1;
      end
    end
    if (reset) begin
      regs_29 <= 1'h0;
    end else begin
      if (_T_950) begin
        regs_29 <= 1'h1;
      end
    end
    if (reset) begin
      regs_30 <= 1'h0;
    end else begin
      if (_T_959) begin
        regs_30 <= 1'h1;
      end
    end
    if (reset) begin
      regs_31 <= 1'h0;
    end else begin
      if (_T_968) begin
        regs_31 <= 1'h1;
      end
    end
    if (reset) begin
      regs_32 <= 1'h0;
    end else begin
      if (_T_977) begin
        regs_32 <= 1'h1;
      end
    end
    if (reset) begin
      regs_33 <= 1'h0;
    end else begin
      if (_T_986) begin
        regs_33 <= 1'h1;
      end
    end
    if (reset) begin
      regs_34 <= 1'h0;
    end else begin
      if (_T_995) begin
        regs_34 <= 1'h1;
      end
    end
    if (reset) begin
      regs_35 <= 1'h0;
    end else begin
      if (_T_1004) begin
        regs_35 <= 1'h1;
      end
    end
    if (reset) begin
      regs_36 <= 1'h0;
    end else begin
      if (_T_1013) begin
        regs_36 <= 1'h1;
      end
    end
    if (reset) begin
      regs_37 <= 1'h0;
    end else begin
      if (_T_1022) begin
        regs_37 <= 1'h1;
      end
    end
    if (reset) begin
      regs_38 <= 1'h0;
    end else begin
      if (_T_1031) begin
        regs_38 <= 1'h1;
      end
    end
    if (reset) begin
      regs_39 <= 1'h0;
    end else begin
      if (_T_1040) begin
        regs_39 <= 1'h1;
      end
    end
    if (reset) begin
      regs_40 <= 1'h0;
    end else begin
      if (_T_1049) begin
        regs_40 <= 1'h1;
      end
    end
    if (reset) begin
      regs_41 <= 1'h0;
    end else begin
      if (_T_1058) begin
        regs_41 <= 1'h1;
      end
    end
    if (reset) begin
      regs_42 <= 1'h0;
    end else begin
      if (_T_1067) begin
        regs_42 <= 1'h1;
      end
    end
    if (reset) begin
      regs_43 <= 1'h0;
    end else begin
      if (_T_1076) begin
        regs_43 <= 1'h1;
      end
    end
    if (reset) begin
      regs_44 <= 1'h0;
    end else begin
      if (_T_1085) begin
        regs_44 <= 1'h1;
      end
    end
    if (reset) begin
      regs_45 <= 1'h0;
    end else begin
      if (_T_1094) begin
        regs_45 <= 1'h1;
      end
    end
    if (reset) begin
      regs_46 <= 1'h0;
    end else begin
      if (_T_1103) begin
        regs_46 <= 1'h1;
      end
    end
    if (reset) begin
      regs_47 <= 1'h0;
    end else begin
      if (_T_1112) begin
        regs_47 <= 1'h1;
      end
    end
    if (reset) begin
      regs_48 <= 1'h0;
    end else begin
      if (_T_1121) begin
        regs_48 <= 1'h1;
      end
    end
    if (reset) begin
      regs_49 <= 1'h0;
    end else begin
      if (_T_1130) begin
        regs_49 <= 1'h1;
      end
    end
    if (reset) begin
      regs_50 <= 1'h0;
    end else begin
      if (_T_1139) begin
        regs_50 <= 1'h1;
      end
    end
    if (reset) begin
      regs_51 <= 1'h0;
    end else begin
      if (_T_1148) begin
        regs_51 <= 1'h1;
      end
    end
    if (reset) begin
      regs_52 <= 1'h0;
    end else begin
      if (_T_1157) begin
        regs_52 <= 1'h1;
      end
    end
    if (reset) begin
      regs_53 <= 1'h0;
    end else begin
      if (_T_1166) begin
        regs_53 <= 1'h1;
      end
    end
    if (reset) begin
      regs_54 <= 1'h0;
    end else begin
      if (_T_1175) begin
        regs_54 <= 1'h1;
      end
    end
    if (reset) begin
      regs_55 <= 1'h0;
    end else begin
      if (_T_1184) begin
        regs_55 <= 1'h1;
      end
    end
    if (reset) begin
      regs_56 <= 1'h0;
    end else begin
      if (_T_1193) begin
        regs_56 <= 1'h1;
      end
    end
    if (reset) begin
      regs_57 <= 1'h0;
    end else begin
      if (_T_1202) begin
        regs_57 <= 1'h1;
      end
    end
    if (reset) begin
      regs_58 <= 1'h0;
    end else begin
      if (_T_1211) begin
        regs_58 <= 1'h1;
      end
    end
    if (reset) begin
      regs_59 <= 1'h0;
    end else begin
      if (_T_1220) begin
        regs_59 <= 1'h1;
      end
    end
    if (reset) begin
      regs_60 <= 1'h0;
    end else begin
      if (_T_1229) begin
        regs_60 <= 1'h1;
      end
    end
    if (reset) begin
      regs_61 <= 1'h0;
    end else begin
      if (_T_1238) begin
        regs_61 <= 1'h1;
      end
    end
    if (reset) begin
      regs_62 <= 1'h0;
    end else begin
      if (_T_1247) begin
        regs_62 <= 1'h1;
      end
    end
    if (reset) begin
      regs_63 <= 1'h0;
    end else begin
      if (_T_1256) begin
        regs_63 <= 1'h1;
      end
    end
  end
endmodule
module FIFO_51( // @[:@100156.2]
  input   clock, // @[:@100157.4]
  input   reset, // @[:@100158.4]
  output  io_in_ready, // @[:@100159.4]
  input   io_in_valid, // @[:@100159.4]
  input   io_out_ready, // @[:@100159.4]
  output  io_out_valid, // @[:@100159.4]
  output  io_out_bits // @[:@100159.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@100425.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@100425.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@100425.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@100425.4]
  wire [5:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@100425.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@100425.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@100425.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@100435.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@100435.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@100435.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@100435.4]
  wire [5:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@100435.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@100435.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@100435.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@100450.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@100450.4]
  wire [5:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@100450.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@100450.4]
  wire [5:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@100450.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@100450.4]
  wire  writeEn; // @[FIFO.scala 30:29:@100423.4]
  wire  readEn; // @[FIFO.scala 31:29:@100424.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@100445.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@100446.4]
  wire  _T_824; // @[FIFO.scala 45:27:@100447.4]
  wire  empty; // @[FIFO.scala 45:24:@100448.4]
  wire  full; // @[FIFO.scala 46:23:@100449.4]
  wire  _T_1657; // @[FIFO.scala 83:17:@101616.4]
  wire  _GEN_64; // @[FIFO.scala 83:29:@101617.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@100425.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@100435.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM_16 FFRAM ( // @[FIFO.scala 49:19:@100450.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_rdata(FFRAM_io_rdata)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@100423.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@100424.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@100446.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@100447.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@100448.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@100449.4]
  assign _T_1657 = writeEn != readEn; // @[FIFO.scala 83:17:@101616.4]
  assign _GEN_64 = _T_1657 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@101617.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@101623.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@101621.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@100655.4]
  assign enqCounter_clock = clock; // @[:@100426.4]
  assign enqCounter_reset = reset; // @[:@100427.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@100433.4]
  assign enqCounter_io_stride = 6'h1; // @[FIFO.scala 37:24:@100434.4]
  assign deqCounter_clock = clock; // @[:@100436.4]
  assign deqCounter_reset = reset; // @[:@100437.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@100443.4]
  assign deqCounter_io_stride = 6'h1; // @[FIFO.scala 41:24:@100444.4]
  assign FFRAM_clock = clock; // @[:@100451.4]
  assign FFRAM_reset = reset; // @[:@100452.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@100651.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@100652.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@100653.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_1657) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module StreamControllerStore( // @[:@101625.2]
  input         clock, // @[:@101626.4]
  input         reset, // @[:@101627.4]
  input         io_dram_cmd_ready, // @[:@101628.4]
  output        io_dram_cmd_valid, // @[:@101628.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@101628.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@101628.4]
  input         io_dram_wdata_ready, // @[:@101628.4]
  output        io_dram_wdata_valid, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_0, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_1, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_2, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_3, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_4, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_5, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_6, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_7, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_8, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_9, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_10, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_11, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_12, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_13, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_14, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_15, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_16, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_17, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_18, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_19, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_20, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_21, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_22, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_23, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_24, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_25, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_26, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_27, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_28, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_29, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_30, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_31, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_32, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_33, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_34, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_35, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_36, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_37, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_38, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_39, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_40, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_41, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_42, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_43, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_44, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_45, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_46, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_47, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_48, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_49, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_50, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_51, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_52, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_53, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_54, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_55, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_56, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_57, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_58, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_59, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_60, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_61, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_62, // @[:@101628.4]
  output [7:0]  io_dram_wdata_bits_wdata_63, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@101628.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@101628.4]
  output        io_dram_wresp_ready, // @[:@101628.4]
  input         io_dram_wresp_valid, // @[:@101628.4]
  output        io_store_cmd_ready, // @[:@101628.4]
  input         io_store_cmd_valid, // @[:@101628.4]
  input  [63:0] io_store_cmd_bits_addr, // @[:@101628.4]
  input  [31:0] io_store_cmd_bits_size, // @[:@101628.4]
  output        io_store_data_ready, // @[:@101628.4]
  input         io_store_data_valid, // @[:@101628.4]
  input  [31:0] io_store_data_bits_wdata_0, // @[:@101628.4]
  input         io_store_data_bits_wstrb, // @[:@101628.4]
  input         io_store_wresp_ready, // @[:@101628.4]
  output        io_store_wresp_valid, // @[:@101628.4]
  output        io_store_wresp_bits // @[:@101628.4]
);
  wire  cmd_clock; // @[StreamController.scala 75:19:@101849.4]
  wire  cmd_reset; // @[StreamController.scala 75:19:@101849.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 75:19:@101849.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 75:19:@101849.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 75:19:@101849.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 75:19:@101849.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 75:19:@101849.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 75:19:@101849.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 75:19:@101849.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 75:19:@101849.4]
  wire  wdata_clock; // @[StreamController.scala 88:21:@102255.4]
  wire  wdata_reset; // @[StreamController.scala 88:21:@102255.4]
  wire  wdata_io_in_ready; // @[StreamController.scala 88:21:@102255.4]
  wire  wdata_io_in_valid; // @[StreamController.scala 88:21:@102255.4]
  wire [31:0] wdata_io_in_bits_data_0; // @[StreamController.scala 88:21:@102255.4]
  wire  wdata_io_in_bits_strobe; // @[StreamController.scala 88:21:@102255.4]
  wire  wdata_io_out_ready; // @[StreamController.scala 88:21:@102255.4]
  wire  wdata_io_out_valid; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_0; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_1; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_2; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_3; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_4; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_5; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_6; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_7; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_8; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_9; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_10; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_11; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_12; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_13; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_14; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_15; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_16; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_17; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_18; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_19; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_20; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_21; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_22; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_23; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_24; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_25; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_26; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_27; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_28; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_29; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_30; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_31; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_32; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_33; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_34; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_35; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_36; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_37; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_38; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_39; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_40; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_41; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_42; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_43; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_44; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_45; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_46; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_47; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_48; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_49; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_50; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_51; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_52; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_53; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_54; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_55; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_56; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_57; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_58; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_59; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_60; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_61; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_62; // @[StreamController.scala 88:21:@102255.4]
  wire [7:0] wdata_io_out_bits_data_63; // @[StreamController.scala 88:21:@102255.4]
  wire [63:0] wdata_io_out_bits_strobe; // @[StreamController.scala 88:21:@102255.4]
  wire  wresp_clock; // @[StreamController.scala 100:21:@102592.4]
  wire  wresp_reset; // @[StreamController.scala 100:21:@102592.4]
  wire  wresp_io_in_ready; // @[StreamController.scala 100:21:@102592.4]
  wire  wresp_io_in_valid; // @[StreamController.scala 100:21:@102592.4]
  wire  wresp_io_out_ready; // @[StreamController.scala 100:21:@102592.4]
  wire  wresp_io_out_valid; // @[StreamController.scala 100:21:@102592.4]
  wire  wresp_io_out_bits; // @[StreamController.scala 100:21:@102592.4]
  wire [25:0] _T_111; // @[StreamController.scala 21:10:@102252.4]
  FIFO cmd ( // @[StreamController.scala 75:19:@101849.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert_1 wdata ( // @[StreamController.scala 88:21:@102255.4]
    .clock(wdata_clock),
    .reset(wdata_reset),
    .io_in_ready(wdata_io_in_ready),
    .io_in_valid(wdata_io_in_valid),
    .io_in_bits_data_0(wdata_io_in_bits_data_0),
    .io_in_bits_strobe(wdata_io_in_bits_strobe),
    .io_out_ready(wdata_io_out_ready),
    .io_out_valid(wdata_io_out_valid),
    .io_out_bits_data_0(wdata_io_out_bits_data_0),
    .io_out_bits_data_1(wdata_io_out_bits_data_1),
    .io_out_bits_data_2(wdata_io_out_bits_data_2),
    .io_out_bits_data_3(wdata_io_out_bits_data_3),
    .io_out_bits_data_4(wdata_io_out_bits_data_4),
    .io_out_bits_data_5(wdata_io_out_bits_data_5),
    .io_out_bits_data_6(wdata_io_out_bits_data_6),
    .io_out_bits_data_7(wdata_io_out_bits_data_7),
    .io_out_bits_data_8(wdata_io_out_bits_data_8),
    .io_out_bits_data_9(wdata_io_out_bits_data_9),
    .io_out_bits_data_10(wdata_io_out_bits_data_10),
    .io_out_bits_data_11(wdata_io_out_bits_data_11),
    .io_out_bits_data_12(wdata_io_out_bits_data_12),
    .io_out_bits_data_13(wdata_io_out_bits_data_13),
    .io_out_bits_data_14(wdata_io_out_bits_data_14),
    .io_out_bits_data_15(wdata_io_out_bits_data_15),
    .io_out_bits_data_16(wdata_io_out_bits_data_16),
    .io_out_bits_data_17(wdata_io_out_bits_data_17),
    .io_out_bits_data_18(wdata_io_out_bits_data_18),
    .io_out_bits_data_19(wdata_io_out_bits_data_19),
    .io_out_bits_data_20(wdata_io_out_bits_data_20),
    .io_out_bits_data_21(wdata_io_out_bits_data_21),
    .io_out_bits_data_22(wdata_io_out_bits_data_22),
    .io_out_bits_data_23(wdata_io_out_bits_data_23),
    .io_out_bits_data_24(wdata_io_out_bits_data_24),
    .io_out_bits_data_25(wdata_io_out_bits_data_25),
    .io_out_bits_data_26(wdata_io_out_bits_data_26),
    .io_out_bits_data_27(wdata_io_out_bits_data_27),
    .io_out_bits_data_28(wdata_io_out_bits_data_28),
    .io_out_bits_data_29(wdata_io_out_bits_data_29),
    .io_out_bits_data_30(wdata_io_out_bits_data_30),
    .io_out_bits_data_31(wdata_io_out_bits_data_31),
    .io_out_bits_data_32(wdata_io_out_bits_data_32),
    .io_out_bits_data_33(wdata_io_out_bits_data_33),
    .io_out_bits_data_34(wdata_io_out_bits_data_34),
    .io_out_bits_data_35(wdata_io_out_bits_data_35),
    .io_out_bits_data_36(wdata_io_out_bits_data_36),
    .io_out_bits_data_37(wdata_io_out_bits_data_37),
    .io_out_bits_data_38(wdata_io_out_bits_data_38),
    .io_out_bits_data_39(wdata_io_out_bits_data_39),
    .io_out_bits_data_40(wdata_io_out_bits_data_40),
    .io_out_bits_data_41(wdata_io_out_bits_data_41),
    .io_out_bits_data_42(wdata_io_out_bits_data_42),
    .io_out_bits_data_43(wdata_io_out_bits_data_43),
    .io_out_bits_data_44(wdata_io_out_bits_data_44),
    .io_out_bits_data_45(wdata_io_out_bits_data_45),
    .io_out_bits_data_46(wdata_io_out_bits_data_46),
    .io_out_bits_data_47(wdata_io_out_bits_data_47),
    .io_out_bits_data_48(wdata_io_out_bits_data_48),
    .io_out_bits_data_49(wdata_io_out_bits_data_49),
    .io_out_bits_data_50(wdata_io_out_bits_data_50),
    .io_out_bits_data_51(wdata_io_out_bits_data_51),
    .io_out_bits_data_52(wdata_io_out_bits_data_52),
    .io_out_bits_data_53(wdata_io_out_bits_data_53),
    .io_out_bits_data_54(wdata_io_out_bits_data_54),
    .io_out_bits_data_55(wdata_io_out_bits_data_55),
    .io_out_bits_data_56(wdata_io_out_bits_data_56),
    .io_out_bits_data_57(wdata_io_out_bits_data_57),
    .io_out_bits_data_58(wdata_io_out_bits_data_58),
    .io_out_bits_data_59(wdata_io_out_bits_data_59),
    .io_out_bits_data_60(wdata_io_out_bits_data_60),
    .io_out_bits_data_61(wdata_io_out_bits_data_61),
    .io_out_bits_data_62(wdata_io_out_bits_data_62),
    .io_out_bits_data_63(wdata_io_out_bits_data_63),
    .io_out_bits_strobe(wdata_io_out_bits_strobe)
  );
  FIFO_51 wresp ( // @[StreamController.scala 100:21:@102592.4]
    .clock(wresp_clock),
    .reset(wresp_reset),
    .io_in_ready(wresp_io_in_ready),
    .io_in_valid(wresp_io_in_valid),
    .io_out_ready(wresp_io_out_ready),
    .io_out_valid(wresp_io_out_valid),
    .io_out_bits(wresp_io_out_bits)
  );
  assign _T_111 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@102252.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 81:21:@102249.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 83:25:@102250.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_111}; // @[StreamController.scala 85:25:@102253.4]
  assign io_dram_wdata_valid = wdata_io_out_valid; // @[StreamController.scala 95:23:@102333.4]
  assign io_dram_wdata_bits_wdata_0 = wdata_io_out_bits_data_0; // @[StreamController.scala 96:28:@102334.4]
  assign io_dram_wdata_bits_wdata_1 = wdata_io_out_bits_data_1; // @[StreamController.scala 96:28:@102335.4]
  assign io_dram_wdata_bits_wdata_2 = wdata_io_out_bits_data_2; // @[StreamController.scala 96:28:@102336.4]
  assign io_dram_wdata_bits_wdata_3 = wdata_io_out_bits_data_3; // @[StreamController.scala 96:28:@102337.4]
  assign io_dram_wdata_bits_wdata_4 = wdata_io_out_bits_data_4; // @[StreamController.scala 96:28:@102338.4]
  assign io_dram_wdata_bits_wdata_5 = wdata_io_out_bits_data_5; // @[StreamController.scala 96:28:@102339.4]
  assign io_dram_wdata_bits_wdata_6 = wdata_io_out_bits_data_6; // @[StreamController.scala 96:28:@102340.4]
  assign io_dram_wdata_bits_wdata_7 = wdata_io_out_bits_data_7; // @[StreamController.scala 96:28:@102341.4]
  assign io_dram_wdata_bits_wdata_8 = wdata_io_out_bits_data_8; // @[StreamController.scala 96:28:@102342.4]
  assign io_dram_wdata_bits_wdata_9 = wdata_io_out_bits_data_9; // @[StreamController.scala 96:28:@102343.4]
  assign io_dram_wdata_bits_wdata_10 = wdata_io_out_bits_data_10; // @[StreamController.scala 96:28:@102344.4]
  assign io_dram_wdata_bits_wdata_11 = wdata_io_out_bits_data_11; // @[StreamController.scala 96:28:@102345.4]
  assign io_dram_wdata_bits_wdata_12 = wdata_io_out_bits_data_12; // @[StreamController.scala 96:28:@102346.4]
  assign io_dram_wdata_bits_wdata_13 = wdata_io_out_bits_data_13; // @[StreamController.scala 96:28:@102347.4]
  assign io_dram_wdata_bits_wdata_14 = wdata_io_out_bits_data_14; // @[StreamController.scala 96:28:@102348.4]
  assign io_dram_wdata_bits_wdata_15 = wdata_io_out_bits_data_15; // @[StreamController.scala 96:28:@102349.4]
  assign io_dram_wdata_bits_wdata_16 = wdata_io_out_bits_data_16; // @[StreamController.scala 96:28:@102350.4]
  assign io_dram_wdata_bits_wdata_17 = wdata_io_out_bits_data_17; // @[StreamController.scala 96:28:@102351.4]
  assign io_dram_wdata_bits_wdata_18 = wdata_io_out_bits_data_18; // @[StreamController.scala 96:28:@102352.4]
  assign io_dram_wdata_bits_wdata_19 = wdata_io_out_bits_data_19; // @[StreamController.scala 96:28:@102353.4]
  assign io_dram_wdata_bits_wdata_20 = wdata_io_out_bits_data_20; // @[StreamController.scala 96:28:@102354.4]
  assign io_dram_wdata_bits_wdata_21 = wdata_io_out_bits_data_21; // @[StreamController.scala 96:28:@102355.4]
  assign io_dram_wdata_bits_wdata_22 = wdata_io_out_bits_data_22; // @[StreamController.scala 96:28:@102356.4]
  assign io_dram_wdata_bits_wdata_23 = wdata_io_out_bits_data_23; // @[StreamController.scala 96:28:@102357.4]
  assign io_dram_wdata_bits_wdata_24 = wdata_io_out_bits_data_24; // @[StreamController.scala 96:28:@102358.4]
  assign io_dram_wdata_bits_wdata_25 = wdata_io_out_bits_data_25; // @[StreamController.scala 96:28:@102359.4]
  assign io_dram_wdata_bits_wdata_26 = wdata_io_out_bits_data_26; // @[StreamController.scala 96:28:@102360.4]
  assign io_dram_wdata_bits_wdata_27 = wdata_io_out_bits_data_27; // @[StreamController.scala 96:28:@102361.4]
  assign io_dram_wdata_bits_wdata_28 = wdata_io_out_bits_data_28; // @[StreamController.scala 96:28:@102362.4]
  assign io_dram_wdata_bits_wdata_29 = wdata_io_out_bits_data_29; // @[StreamController.scala 96:28:@102363.4]
  assign io_dram_wdata_bits_wdata_30 = wdata_io_out_bits_data_30; // @[StreamController.scala 96:28:@102364.4]
  assign io_dram_wdata_bits_wdata_31 = wdata_io_out_bits_data_31; // @[StreamController.scala 96:28:@102365.4]
  assign io_dram_wdata_bits_wdata_32 = wdata_io_out_bits_data_32; // @[StreamController.scala 96:28:@102366.4]
  assign io_dram_wdata_bits_wdata_33 = wdata_io_out_bits_data_33; // @[StreamController.scala 96:28:@102367.4]
  assign io_dram_wdata_bits_wdata_34 = wdata_io_out_bits_data_34; // @[StreamController.scala 96:28:@102368.4]
  assign io_dram_wdata_bits_wdata_35 = wdata_io_out_bits_data_35; // @[StreamController.scala 96:28:@102369.4]
  assign io_dram_wdata_bits_wdata_36 = wdata_io_out_bits_data_36; // @[StreamController.scala 96:28:@102370.4]
  assign io_dram_wdata_bits_wdata_37 = wdata_io_out_bits_data_37; // @[StreamController.scala 96:28:@102371.4]
  assign io_dram_wdata_bits_wdata_38 = wdata_io_out_bits_data_38; // @[StreamController.scala 96:28:@102372.4]
  assign io_dram_wdata_bits_wdata_39 = wdata_io_out_bits_data_39; // @[StreamController.scala 96:28:@102373.4]
  assign io_dram_wdata_bits_wdata_40 = wdata_io_out_bits_data_40; // @[StreamController.scala 96:28:@102374.4]
  assign io_dram_wdata_bits_wdata_41 = wdata_io_out_bits_data_41; // @[StreamController.scala 96:28:@102375.4]
  assign io_dram_wdata_bits_wdata_42 = wdata_io_out_bits_data_42; // @[StreamController.scala 96:28:@102376.4]
  assign io_dram_wdata_bits_wdata_43 = wdata_io_out_bits_data_43; // @[StreamController.scala 96:28:@102377.4]
  assign io_dram_wdata_bits_wdata_44 = wdata_io_out_bits_data_44; // @[StreamController.scala 96:28:@102378.4]
  assign io_dram_wdata_bits_wdata_45 = wdata_io_out_bits_data_45; // @[StreamController.scala 96:28:@102379.4]
  assign io_dram_wdata_bits_wdata_46 = wdata_io_out_bits_data_46; // @[StreamController.scala 96:28:@102380.4]
  assign io_dram_wdata_bits_wdata_47 = wdata_io_out_bits_data_47; // @[StreamController.scala 96:28:@102381.4]
  assign io_dram_wdata_bits_wdata_48 = wdata_io_out_bits_data_48; // @[StreamController.scala 96:28:@102382.4]
  assign io_dram_wdata_bits_wdata_49 = wdata_io_out_bits_data_49; // @[StreamController.scala 96:28:@102383.4]
  assign io_dram_wdata_bits_wdata_50 = wdata_io_out_bits_data_50; // @[StreamController.scala 96:28:@102384.4]
  assign io_dram_wdata_bits_wdata_51 = wdata_io_out_bits_data_51; // @[StreamController.scala 96:28:@102385.4]
  assign io_dram_wdata_bits_wdata_52 = wdata_io_out_bits_data_52; // @[StreamController.scala 96:28:@102386.4]
  assign io_dram_wdata_bits_wdata_53 = wdata_io_out_bits_data_53; // @[StreamController.scala 96:28:@102387.4]
  assign io_dram_wdata_bits_wdata_54 = wdata_io_out_bits_data_54; // @[StreamController.scala 96:28:@102388.4]
  assign io_dram_wdata_bits_wdata_55 = wdata_io_out_bits_data_55; // @[StreamController.scala 96:28:@102389.4]
  assign io_dram_wdata_bits_wdata_56 = wdata_io_out_bits_data_56; // @[StreamController.scala 96:28:@102390.4]
  assign io_dram_wdata_bits_wdata_57 = wdata_io_out_bits_data_57; // @[StreamController.scala 96:28:@102391.4]
  assign io_dram_wdata_bits_wdata_58 = wdata_io_out_bits_data_58; // @[StreamController.scala 96:28:@102392.4]
  assign io_dram_wdata_bits_wdata_59 = wdata_io_out_bits_data_59; // @[StreamController.scala 96:28:@102393.4]
  assign io_dram_wdata_bits_wdata_60 = wdata_io_out_bits_data_60; // @[StreamController.scala 96:28:@102394.4]
  assign io_dram_wdata_bits_wdata_61 = wdata_io_out_bits_data_61; // @[StreamController.scala 96:28:@102395.4]
  assign io_dram_wdata_bits_wdata_62 = wdata_io_out_bits_data_62; // @[StreamController.scala 96:28:@102396.4]
  assign io_dram_wdata_bits_wdata_63 = wdata_io_out_bits_data_63; // @[StreamController.scala 96:28:@102397.4]
  assign io_dram_wdata_bits_wstrb_0 = wdata_io_out_bits_strobe[63]; // @[StreamController.scala 97:28:@102527.4]
  assign io_dram_wdata_bits_wstrb_1 = wdata_io_out_bits_strobe[62]; // @[StreamController.scala 97:28:@102528.4]
  assign io_dram_wdata_bits_wstrb_2 = wdata_io_out_bits_strobe[61]; // @[StreamController.scala 97:28:@102529.4]
  assign io_dram_wdata_bits_wstrb_3 = wdata_io_out_bits_strobe[60]; // @[StreamController.scala 97:28:@102530.4]
  assign io_dram_wdata_bits_wstrb_4 = wdata_io_out_bits_strobe[59]; // @[StreamController.scala 97:28:@102531.4]
  assign io_dram_wdata_bits_wstrb_5 = wdata_io_out_bits_strobe[58]; // @[StreamController.scala 97:28:@102532.4]
  assign io_dram_wdata_bits_wstrb_6 = wdata_io_out_bits_strobe[57]; // @[StreamController.scala 97:28:@102533.4]
  assign io_dram_wdata_bits_wstrb_7 = wdata_io_out_bits_strobe[56]; // @[StreamController.scala 97:28:@102534.4]
  assign io_dram_wdata_bits_wstrb_8 = wdata_io_out_bits_strobe[55]; // @[StreamController.scala 97:28:@102535.4]
  assign io_dram_wdata_bits_wstrb_9 = wdata_io_out_bits_strobe[54]; // @[StreamController.scala 97:28:@102536.4]
  assign io_dram_wdata_bits_wstrb_10 = wdata_io_out_bits_strobe[53]; // @[StreamController.scala 97:28:@102537.4]
  assign io_dram_wdata_bits_wstrb_11 = wdata_io_out_bits_strobe[52]; // @[StreamController.scala 97:28:@102538.4]
  assign io_dram_wdata_bits_wstrb_12 = wdata_io_out_bits_strobe[51]; // @[StreamController.scala 97:28:@102539.4]
  assign io_dram_wdata_bits_wstrb_13 = wdata_io_out_bits_strobe[50]; // @[StreamController.scala 97:28:@102540.4]
  assign io_dram_wdata_bits_wstrb_14 = wdata_io_out_bits_strobe[49]; // @[StreamController.scala 97:28:@102541.4]
  assign io_dram_wdata_bits_wstrb_15 = wdata_io_out_bits_strobe[48]; // @[StreamController.scala 97:28:@102542.4]
  assign io_dram_wdata_bits_wstrb_16 = wdata_io_out_bits_strobe[47]; // @[StreamController.scala 97:28:@102543.4]
  assign io_dram_wdata_bits_wstrb_17 = wdata_io_out_bits_strobe[46]; // @[StreamController.scala 97:28:@102544.4]
  assign io_dram_wdata_bits_wstrb_18 = wdata_io_out_bits_strobe[45]; // @[StreamController.scala 97:28:@102545.4]
  assign io_dram_wdata_bits_wstrb_19 = wdata_io_out_bits_strobe[44]; // @[StreamController.scala 97:28:@102546.4]
  assign io_dram_wdata_bits_wstrb_20 = wdata_io_out_bits_strobe[43]; // @[StreamController.scala 97:28:@102547.4]
  assign io_dram_wdata_bits_wstrb_21 = wdata_io_out_bits_strobe[42]; // @[StreamController.scala 97:28:@102548.4]
  assign io_dram_wdata_bits_wstrb_22 = wdata_io_out_bits_strobe[41]; // @[StreamController.scala 97:28:@102549.4]
  assign io_dram_wdata_bits_wstrb_23 = wdata_io_out_bits_strobe[40]; // @[StreamController.scala 97:28:@102550.4]
  assign io_dram_wdata_bits_wstrb_24 = wdata_io_out_bits_strobe[39]; // @[StreamController.scala 97:28:@102551.4]
  assign io_dram_wdata_bits_wstrb_25 = wdata_io_out_bits_strobe[38]; // @[StreamController.scala 97:28:@102552.4]
  assign io_dram_wdata_bits_wstrb_26 = wdata_io_out_bits_strobe[37]; // @[StreamController.scala 97:28:@102553.4]
  assign io_dram_wdata_bits_wstrb_27 = wdata_io_out_bits_strobe[36]; // @[StreamController.scala 97:28:@102554.4]
  assign io_dram_wdata_bits_wstrb_28 = wdata_io_out_bits_strobe[35]; // @[StreamController.scala 97:28:@102555.4]
  assign io_dram_wdata_bits_wstrb_29 = wdata_io_out_bits_strobe[34]; // @[StreamController.scala 97:28:@102556.4]
  assign io_dram_wdata_bits_wstrb_30 = wdata_io_out_bits_strobe[33]; // @[StreamController.scala 97:28:@102557.4]
  assign io_dram_wdata_bits_wstrb_31 = wdata_io_out_bits_strobe[32]; // @[StreamController.scala 97:28:@102558.4]
  assign io_dram_wdata_bits_wstrb_32 = wdata_io_out_bits_strobe[31]; // @[StreamController.scala 97:28:@102559.4]
  assign io_dram_wdata_bits_wstrb_33 = wdata_io_out_bits_strobe[30]; // @[StreamController.scala 97:28:@102560.4]
  assign io_dram_wdata_bits_wstrb_34 = wdata_io_out_bits_strobe[29]; // @[StreamController.scala 97:28:@102561.4]
  assign io_dram_wdata_bits_wstrb_35 = wdata_io_out_bits_strobe[28]; // @[StreamController.scala 97:28:@102562.4]
  assign io_dram_wdata_bits_wstrb_36 = wdata_io_out_bits_strobe[27]; // @[StreamController.scala 97:28:@102563.4]
  assign io_dram_wdata_bits_wstrb_37 = wdata_io_out_bits_strobe[26]; // @[StreamController.scala 97:28:@102564.4]
  assign io_dram_wdata_bits_wstrb_38 = wdata_io_out_bits_strobe[25]; // @[StreamController.scala 97:28:@102565.4]
  assign io_dram_wdata_bits_wstrb_39 = wdata_io_out_bits_strobe[24]; // @[StreamController.scala 97:28:@102566.4]
  assign io_dram_wdata_bits_wstrb_40 = wdata_io_out_bits_strobe[23]; // @[StreamController.scala 97:28:@102567.4]
  assign io_dram_wdata_bits_wstrb_41 = wdata_io_out_bits_strobe[22]; // @[StreamController.scala 97:28:@102568.4]
  assign io_dram_wdata_bits_wstrb_42 = wdata_io_out_bits_strobe[21]; // @[StreamController.scala 97:28:@102569.4]
  assign io_dram_wdata_bits_wstrb_43 = wdata_io_out_bits_strobe[20]; // @[StreamController.scala 97:28:@102570.4]
  assign io_dram_wdata_bits_wstrb_44 = wdata_io_out_bits_strobe[19]; // @[StreamController.scala 97:28:@102571.4]
  assign io_dram_wdata_bits_wstrb_45 = wdata_io_out_bits_strobe[18]; // @[StreamController.scala 97:28:@102572.4]
  assign io_dram_wdata_bits_wstrb_46 = wdata_io_out_bits_strobe[17]; // @[StreamController.scala 97:28:@102573.4]
  assign io_dram_wdata_bits_wstrb_47 = wdata_io_out_bits_strobe[16]; // @[StreamController.scala 97:28:@102574.4]
  assign io_dram_wdata_bits_wstrb_48 = wdata_io_out_bits_strobe[15]; // @[StreamController.scala 97:28:@102575.4]
  assign io_dram_wdata_bits_wstrb_49 = wdata_io_out_bits_strobe[14]; // @[StreamController.scala 97:28:@102576.4]
  assign io_dram_wdata_bits_wstrb_50 = wdata_io_out_bits_strobe[13]; // @[StreamController.scala 97:28:@102577.4]
  assign io_dram_wdata_bits_wstrb_51 = wdata_io_out_bits_strobe[12]; // @[StreamController.scala 97:28:@102578.4]
  assign io_dram_wdata_bits_wstrb_52 = wdata_io_out_bits_strobe[11]; // @[StreamController.scala 97:28:@102579.4]
  assign io_dram_wdata_bits_wstrb_53 = wdata_io_out_bits_strobe[10]; // @[StreamController.scala 97:28:@102580.4]
  assign io_dram_wdata_bits_wstrb_54 = wdata_io_out_bits_strobe[9]; // @[StreamController.scala 97:28:@102581.4]
  assign io_dram_wdata_bits_wstrb_55 = wdata_io_out_bits_strobe[8]; // @[StreamController.scala 97:28:@102582.4]
  assign io_dram_wdata_bits_wstrb_56 = wdata_io_out_bits_strobe[7]; // @[StreamController.scala 97:28:@102583.4]
  assign io_dram_wdata_bits_wstrb_57 = wdata_io_out_bits_strobe[6]; // @[StreamController.scala 97:28:@102584.4]
  assign io_dram_wdata_bits_wstrb_58 = wdata_io_out_bits_strobe[5]; // @[StreamController.scala 97:28:@102585.4]
  assign io_dram_wdata_bits_wstrb_59 = wdata_io_out_bits_strobe[4]; // @[StreamController.scala 97:28:@102586.4]
  assign io_dram_wdata_bits_wstrb_60 = wdata_io_out_bits_strobe[3]; // @[StreamController.scala 97:28:@102587.4]
  assign io_dram_wdata_bits_wstrb_61 = wdata_io_out_bits_strobe[2]; // @[StreamController.scala 97:28:@102588.4]
  assign io_dram_wdata_bits_wstrb_62 = wdata_io_out_bits_strobe[1]; // @[StreamController.scala 97:28:@102589.4]
  assign io_dram_wdata_bits_wstrb_63 = wdata_io_out_bits_strobe[0]; // @[StreamController.scala 97:28:@102590.4]
  assign io_dram_wresp_ready = wresp_io_in_ready; // @[StreamController.scala 104:23:@102859.4]
  assign io_store_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 79:22:@102247.4]
  assign io_store_data_ready = wdata_io_in_ready; // @[StreamController.scala 93:23:@102332.4]
  assign io_store_wresp_valid = wresp_io_out_valid; // @[StreamController.scala 106:24:@102860.4]
  assign io_store_wresp_bits = wresp_io_out_bits; // @[StreamController.scala 107:23:@102861.4]
  assign cmd_clock = clock; // @[:@101850.4]
  assign cmd_reset = reset; // @[:@101851.4]
  assign cmd_io_in_valid = io_store_cmd_valid; // @[StreamController.scala 77:19:@102244.4]
  assign cmd_io_in_bits_addr = io_store_cmd_bits_addr; // @[StreamController.scala 78:18:@102246.4]
  assign cmd_io_in_bits_size = io_store_cmd_bits_size; // @[StreamController.scala 78:18:@102245.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 80:20:@102248.4]
  assign wdata_clock = clock; // @[:@102256.4]
  assign wdata_reset = reset; // @[:@102257.4]
  assign wdata_io_in_valid = io_store_data_valid; // @[StreamController.scala 90:21:@102329.4]
  assign wdata_io_in_bits_data_0 = io_store_data_bits_wdata_0; // @[StreamController.scala 91:25:@102330.4]
  assign wdata_io_in_bits_strobe = io_store_data_bits_wstrb; // @[StreamController.scala 92:27:@102331.4]
  assign wdata_io_out_ready = io_dram_wdata_ready; // @[StreamController.scala 98:22:@102591.4]
  assign wresp_clock = clock; // @[:@102593.4]
  assign wresp_reset = reset; // @[:@102594.4]
  assign wresp_io_in_valid = io_dram_wresp_valid; // @[StreamController.scala 102:21:@102857.4]
  assign wresp_io_out_ready = io_store_wresp_ready; // @[StreamController.scala 108:22:@102862.4]
endmodule
module MuxN( // @[:@102928.2]
  input  [63:0] io_ins_0_addr, // @[:@102931.4]
  input  [31:0] io_ins_0_size, // @[:@102931.4]
  input  [63:0] io_ins_1_addr, // @[:@102931.4]
  input  [31:0] io_ins_1_size, // @[:@102931.4]
  input         io_sel, // @[:@102931.4]
  output [63:0] io_out_addr, // @[:@102931.4]
  output [31:0] io_out_size, // @[:@102931.4]
  output        io_out_isWr, // @[:@102931.4]
  output [31:0] io_out_tag // @[:@102931.4]
);
  assign io_out_addr = io_sel ? io_ins_1_addr : io_ins_0_addr; // @[MuxN.scala 16:10:@102937.4]
  assign io_out_size = io_sel ? io_ins_1_size : io_ins_0_size; // @[MuxN.scala 16:10:@102936.4]
  assign io_out_isWr = io_sel; // @[MuxN.scala 16:10:@102934.4]
  assign io_out_tag = io_sel ? 32'h1 : 32'h0; // @[MuxN.scala 16:10:@102933.4]
endmodule
module MuxPipe( // @[:@102939.2]
  output        io_in_ready, // @[:@102942.4]
  input         io_in_valid, // @[:@102942.4]
  input  [63:0] io_in_bits_0_addr, // @[:@102942.4]
  input  [31:0] io_in_bits_0_size, // @[:@102942.4]
  input  [63:0] io_in_bits_1_addr, // @[:@102942.4]
  input  [31:0] io_in_bits_1_size, // @[:@102942.4]
  input         io_sel, // @[:@102942.4]
  input         io_out_ready, // @[:@102942.4]
  output        io_out_valid, // @[:@102942.4]
  output [63:0] io_out_bits_addr, // @[:@102942.4]
  output [31:0] io_out_bits_size, // @[:@102942.4]
  output        io_out_bits_isWr, // @[:@102942.4]
  output [31:0] io_out_bits_tag // @[:@102942.4]
);
  wire [63:0] MuxN_io_ins_0_addr; // @[MuxN.scala 40:23:@102957.4]
  wire [31:0] MuxN_io_ins_0_size; // @[MuxN.scala 40:23:@102957.4]
  wire [63:0] MuxN_io_ins_1_addr; // @[MuxN.scala 40:23:@102957.4]
  wire [31:0] MuxN_io_ins_1_size; // @[MuxN.scala 40:23:@102957.4]
  wire  MuxN_io_sel; // @[MuxN.scala 40:23:@102957.4]
  wire [63:0] MuxN_io_out_addr; // @[MuxN.scala 40:23:@102957.4]
  wire [31:0] MuxN_io_out_size; // @[MuxN.scala 40:23:@102957.4]
  wire  MuxN_io_out_isWr; // @[MuxN.scala 40:23:@102957.4]
  wire [31:0] MuxN_io_out_tag; // @[MuxN.scala 40:23:@102957.4]
  wire  _T_46; // @[MuxN.scala 28:31:@102944.4]
  MuxN MuxN ( // @[MuxN.scala 40:23:@102957.4]
    .io_ins_0_addr(MuxN_io_ins_0_addr),
    .io_ins_0_size(MuxN_io_ins_0_size),
    .io_ins_1_addr(MuxN_io_ins_1_addr),
    .io_ins_1_size(MuxN_io_ins_1_size),
    .io_sel(MuxN_io_sel),
    .io_out_addr(MuxN_io_out_addr),
    .io_out_size(MuxN_io_out_size),
    .io_out_isWr(MuxN_io_out_isWr),
    .io_out_tag(MuxN_io_out_tag)
  );
  assign _T_46 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@102944.4]
  assign io_in_ready = io_out_ready | _T_46; // @[MuxN.scala 71:15:@102973.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@102972.4]
  assign io_out_bits_addr = MuxN_io_out_addr; // @[MuxN.scala 72:15:@102978.4]
  assign io_out_bits_size = MuxN_io_out_size; // @[MuxN.scala 72:15:@102977.4]
  assign io_out_bits_isWr = MuxN_io_out_isWr; // @[MuxN.scala 72:15:@102975.4]
  assign io_out_bits_tag = MuxN_io_out_tag; // @[MuxN.scala 72:15:@102974.4]
  assign MuxN_io_ins_0_addr = io_in_bits_0_addr; // @[MuxN.scala 41:18:@102964.4]
  assign MuxN_io_ins_0_size = io_in_bits_0_size; // @[MuxN.scala 41:18:@102963.4]
  assign MuxN_io_ins_1_addr = io_in_bits_1_addr; // @[MuxN.scala 41:18:@102969.4]
  assign MuxN_io_ins_1_size = io_in_bits_1_size; // @[MuxN.scala 41:18:@102968.4]
  assign MuxN_io_sel = io_sel; // @[MuxN.scala 44:18:@102971.4]
endmodule
module MuxN_1( // @[:@102980.2]
  input  [7:0] io_ins_1_wdata_0, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_1, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_2, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_3, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_4, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_5, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_6, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_7, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_8, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_9, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_10, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_11, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_12, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_13, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_14, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_15, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_16, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_17, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_18, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_19, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_20, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_21, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_22, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_23, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_24, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_25, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_26, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_27, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_28, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_29, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_30, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_31, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_32, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_33, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_34, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_35, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_36, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_37, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_38, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_39, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_40, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_41, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_42, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_43, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_44, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_45, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_46, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_47, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_48, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_49, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_50, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_51, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_52, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_53, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_54, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_55, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_56, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_57, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_58, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_59, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_60, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_61, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_62, // @[:@102983.4]
  input  [7:0] io_ins_1_wdata_63, // @[:@102983.4]
  input        io_ins_1_wstrb_0, // @[:@102983.4]
  input        io_ins_1_wstrb_1, // @[:@102983.4]
  input        io_ins_1_wstrb_2, // @[:@102983.4]
  input        io_ins_1_wstrb_3, // @[:@102983.4]
  input        io_ins_1_wstrb_4, // @[:@102983.4]
  input        io_ins_1_wstrb_5, // @[:@102983.4]
  input        io_ins_1_wstrb_6, // @[:@102983.4]
  input        io_ins_1_wstrb_7, // @[:@102983.4]
  input        io_ins_1_wstrb_8, // @[:@102983.4]
  input        io_ins_1_wstrb_9, // @[:@102983.4]
  input        io_ins_1_wstrb_10, // @[:@102983.4]
  input        io_ins_1_wstrb_11, // @[:@102983.4]
  input        io_ins_1_wstrb_12, // @[:@102983.4]
  input        io_ins_1_wstrb_13, // @[:@102983.4]
  input        io_ins_1_wstrb_14, // @[:@102983.4]
  input        io_ins_1_wstrb_15, // @[:@102983.4]
  input        io_ins_1_wstrb_16, // @[:@102983.4]
  input        io_ins_1_wstrb_17, // @[:@102983.4]
  input        io_ins_1_wstrb_18, // @[:@102983.4]
  input        io_ins_1_wstrb_19, // @[:@102983.4]
  input        io_ins_1_wstrb_20, // @[:@102983.4]
  input        io_ins_1_wstrb_21, // @[:@102983.4]
  input        io_ins_1_wstrb_22, // @[:@102983.4]
  input        io_ins_1_wstrb_23, // @[:@102983.4]
  input        io_ins_1_wstrb_24, // @[:@102983.4]
  input        io_ins_1_wstrb_25, // @[:@102983.4]
  input        io_ins_1_wstrb_26, // @[:@102983.4]
  input        io_ins_1_wstrb_27, // @[:@102983.4]
  input        io_ins_1_wstrb_28, // @[:@102983.4]
  input        io_ins_1_wstrb_29, // @[:@102983.4]
  input        io_ins_1_wstrb_30, // @[:@102983.4]
  input        io_ins_1_wstrb_31, // @[:@102983.4]
  input        io_ins_1_wstrb_32, // @[:@102983.4]
  input        io_ins_1_wstrb_33, // @[:@102983.4]
  input        io_ins_1_wstrb_34, // @[:@102983.4]
  input        io_ins_1_wstrb_35, // @[:@102983.4]
  input        io_ins_1_wstrb_36, // @[:@102983.4]
  input        io_ins_1_wstrb_37, // @[:@102983.4]
  input        io_ins_1_wstrb_38, // @[:@102983.4]
  input        io_ins_1_wstrb_39, // @[:@102983.4]
  input        io_ins_1_wstrb_40, // @[:@102983.4]
  input        io_ins_1_wstrb_41, // @[:@102983.4]
  input        io_ins_1_wstrb_42, // @[:@102983.4]
  input        io_ins_1_wstrb_43, // @[:@102983.4]
  input        io_ins_1_wstrb_44, // @[:@102983.4]
  input        io_ins_1_wstrb_45, // @[:@102983.4]
  input        io_ins_1_wstrb_46, // @[:@102983.4]
  input        io_ins_1_wstrb_47, // @[:@102983.4]
  input        io_ins_1_wstrb_48, // @[:@102983.4]
  input        io_ins_1_wstrb_49, // @[:@102983.4]
  input        io_ins_1_wstrb_50, // @[:@102983.4]
  input        io_ins_1_wstrb_51, // @[:@102983.4]
  input        io_ins_1_wstrb_52, // @[:@102983.4]
  input        io_ins_1_wstrb_53, // @[:@102983.4]
  input        io_ins_1_wstrb_54, // @[:@102983.4]
  input        io_ins_1_wstrb_55, // @[:@102983.4]
  input        io_ins_1_wstrb_56, // @[:@102983.4]
  input        io_ins_1_wstrb_57, // @[:@102983.4]
  input        io_ins_1_wstrb_58, // @[:@102983.4]
  input        io_ins_1_wstrb_59, // @[:@102983.4]
  input        io_ins_1_wstrb_60, // @[:@102983.4]
  input        io_ins_1_wstrb_61, // @[:@102983.4]
  input        io_ins_1_wstrb_62, // @[:@102983.4]
  input        io_ins_1_wstrb_63, // @[:@102983.4]
  input        io_sel, // @[:@102983.4]
  output [7:0] io_out_wdata_0, // @[:@102983.4]
  output [7:0] io_out_wdata_1, // @[:@102983.4]
  output [7:0] io_out_wdata_2, // @[:@102983.4]
  output [7:0] io_out_wdata_3, // @[:@102983.4]
  output [7:0] io_out_wdata_4, // @[:@102983.4]
  output [7:0] io_out_wdata_5, // @[:@102983.4]
  output [7:0] io_out_wdata_6, // @[:@102983.4]
  output [7:0] io_out_wdata_7, // @[:@102983.4]
  output [7:0] io_out_wdata_8, // @[:@102983.4]
  output [7:0] io_out_wdata_9, // @[:@102983.4]
  output [7:0] io_out_wdata_10, // @[:@102983.4]
  output [7:0] io_out_wdata_11, // @[:@102983.4]
  output [7:0] io_out_wdata_12, // @[:@102983.4]
  output [7:0] io_out_wdata_13, // @[:@102983.4]
  output [7:0] io_out_wdata_14, // @[:@102983.4]
  output [7:0] io_out_wdata_15, // @[:@102983.4]
  output [7:0] io_out_wdata_16, // @[:@102983.4]
  output [7:0] io_out_wdata_17, // @[:@102983.4]
  output [7:0] io_out_wdata_18, // @[:@102983.4]
  output [7:0] io_out_wdata_19, // @[:@102983.4]
  output [7:0] io_out_wdata_20, // @[:@102983.4]
  output [7:0] io_out_wdata_21, // @[:@102983.4]
  output [7:0] io_out_wdata_22, // @[:@102983.4]
  output [7:0] io_out_wdata_23, // @[:@102983.4]
  output [7:0] io_out_wdata_24, // @[:@102983.4]
  output [7:0] io_out_wdata_25, // @[:@102983.4]
  output [7:0] io_out_wdata_26, // @[:@102983.4]
  output [7:0] io_out_wdata_27, // @[:@102983.4]
  output [7:0] io_out_wdata_28, // @[:@102983.4]
  output [7:0] io_out_wdata_29, // @[:@102983.4]
  output [7:0] io_out_wdata_30, // @[:@102983.4]
  output [7:0] io_out_wdata_31, // @[:@102983.4]
  output [7:0] io_out_wdata_32, // @[:@102983.4]
  output [7:0] io_out_wdata_33, // @[:@102983.4]
  output [7:0] io_out_wdata_34, // @[:@102983.4]
  output [7:0] io_out_wdata_35, // @[:@102983.4]
  output [7:0] io_out_wdata_36, // @[:@102983.4]
  output [7:0] io_out_wdata_37, // @[:@102983.4]
  output [7:0] io_out_wdata_38, // @[:@102983.4]
  output [7:0] io_out_wdata_39, // @[:@102983.4]
  output [7:0] io_out_wdata_40, // @[:@102983.4]
  output [7:0] io_out_wdata_41, // @[:@102983.4]
  output [7:0] io_out_wdata_42, // @[:@102983.4]
  output [7:0] io_out_wdata_43, // @[:@102983.4]
  output [7:0] io_out_wdata_44, // @[:@102983.4]
  output [7:0] io_out_wdata_45, // @[:@102983.4]
  output [7:0] io_out_wdata_46, // @[:@102983.4]
  output [7:0] io_out_wdata_47, // @[:@102983.4]
  output [7:0] io_out_wdata_48, // @[:@102983.4]
  output [7:0] io_out_wdata_49, // @[:@102983.4]
  output [7:0] io_out_wdata_50, // @[:@102983.4]
  output [7:0] io_out_wdata_51, // @[:@102983.4]
  output [7:0] io_out_wdata_52, // @[:@102983.4]
  output [7:0] io_out_wdata_53, // @[:@102983.4]
  output [7:0] io_out_wdata_54, // @[:@102983.4]
  output [7:0] io_out_wdata_55, // @[:@102983.4]
  output [7:0] io_out_wdata_56, // @[:@102983.4]
  output [7:0] io_out_wdata_57, // @[:@102983.4]
  output [7:0] io_out_wdata_58, // @[:@102983.4]
  output [7:0] io_out_wdata_59, // @[:@102983.4]
  output [7:0] io_out_wdata_60, // @[:@102983.4]
  output [7:0] io_out_wdata_61, // @[:@102983.4]
  output [7:0] io_out_wdata_62, // @[:@102983.4]
  output [7:0] io_out_wdata_63, // @[:@102983.4]
  output       io_out_wstrb_0, // @[:@102983.4]
  output       io_out_wstrb_1, // @[:@102983.4]
  output       io_out_wstrb_2, // @[:@102983.4]
  output       io_out_wstrb_3, // @[:@102983.4]
  output       io_out_wstrb_4, // @[:@102983.4]
  output       io_out_wstrb_5, // @[:@102983.4]
  output       io_out_wstrb_6, // @[:@102983.4]
  output       io_out_wstrb_7, // @[:@102983.4]
  output       io_out_wstrb_8, // @[:@102983.4]
  output       io_out_wstrb_9, // @[:@102983.4]
  output       io_out_wstrb_10, // @[:@102983.4]
  output       io_out_wstrb_11, // @[:@102983.4]
  output       io_out_wstrb_12, // @[:@102983.4]
  output       io_out_wstrb_13, // @[:@102983.4]
  output       io_out_wstrb_14, // @[:@102983.4]
  output       io_out_wstrb_15, // @[:@102983.4]
  output       io_out_wstrb_16, // @[:@102983.4]
  output       io_out_wstrb_17, // @[:@102983.4]
  output       io_out_wstrb_18, // @[:@102983.4]
  output       io_out_wstrb_19, // @[:@102983.4]
  output       io_out_wstrb_20, // @[:@102983.4]
  output       io_out_wstrb_21, // @[:@102983.4]
  output       io_out_wstrb_22, // @[:@102983.4]
  output       io_out_wstrb_23, // @[:@102983.4]
  output       io_out_wstrb_24, // @[:@102983.4]
  output       io_out_wstrb_25, // @[:@102983.4]
  output       io_out_wstrb_26, // @[:@102983.4]
  output       io_out_wstrb_27, // @[:@102983.4]
  output       io_out_wstrb_28, // @[:@102983.4]
  output       io_out_wstrb_29, // @[:@102983.4]
  output       io_out_wstrb_30, // @[:@102983.4]
  output       io_out_wstrb_31, // @[:@102983.4]
  output       io_out_wstrb_32, // @[:@102983.4]
  output       io_out_wstrb_33, // @[:@102983.4]
  output       io_out_wstrb_34, // @[:@102983.4]
  output       io_out_wstrb_35, // @[:@102983.4]
  output       io_out_wstrb_36, // @[:@102983.4]
  output       io_out_wstrb_37, // @[:@102983.4]
  output       io_out_wstrb_38, // @[:@102983.4]
  output       io_out_wstrb_39, // @[:@102983.4]
  output       io_out_wstrb_40, // @[:@102983.4]
  output       io_out_wstrb_41, // @[:@102983.4]
  output       io_out_wstrb_42, // @[:@102983.4]
  output       io_out_wstrb_43, // @[:@102983.4]
  output       io_out_wstrb_44, // @[:@102983.4]
  output       io_out_wstrb_45, // @[:@102983.4]
  output       io_out_wstrb_46, // @[:@102983.4]
  output       io_out_wstrb_47, // @[:@102983.4]
  output       io_out_wstrb_48, // @[:@102983.4]
  output       io_out_wstrb_49, // @[:@102983.4]
  output       io_out_wstrb_50, // @[:@102983.4]
  output       io_out_wstrb_51, // @[:@102983.4]
  output       io_out_wstrb_52, // @[:@102983.4]
  output       io_out_wstrb_53, // @[:@102983.4]
  output       io_out_wstrb_54, // @[:@102983.4]
  output       io_out_wstrb_55, // @[:@102983.4]
  output       io_out_wstrb_56, // @[:@102983.4]
  output       io_out_wstrb_57, // @[:@102983.4]
  output       io_out_wstrb_58, // @[:@102983.4]
  output       io_out_wstrb_59, // @[:@102983.4]
  output       io_out_wstrb_60, // @[:@102983.4]
  output       io_out_wstrb_61, // @[:@102983.4]
  output       io_out_wstrb_62, // @[:@102983.4]
  output       io_out_wstrb_63 // @[:@102983.4]
);
  assign io_out_wdata_0 = io_sel ? io_ins_1_wdata_0 : 8'h0; // @[MuxN.scala 16:10:@103050.4]
  assign io_out_wdata_1 = io_sel ? io_ins_1_wdata_1 : 8'h0; // @[MuxN.scala 16:10:@103051.4]
  assign io_out_wdata_2 = io_sel ? io_ins_1_wdata_2 : 8'h0; // @[MuxN.scala 16:10:@103052.4]
  assign io_out_wdata_3 = io_sel ? io_ins_1_wdata_3 : 8'h0; // @[MuxN.scala 16:10:@103053.4]
  assign io_out_wdata_4 = io_sel ? io_ins_1_wdata_4 : 8'h0; // @[MuxN.scala 16:10:@103054.4]
  assign io_out_wdata_5 = io_sel ? io_ins_1_wdata_5 : 8'h0; // @[MuxN.scala 16:10:@103055.4]
  assign io_out_wdata_6 = io_sel ? io_ins_1_wdata_6 : 8'h0; // @[MuxN.scala 16:10:@103056.4]
  assign io_out_wdata_7 = io_sel ? io_ins_1_wdata_7 : 8'h0; // @[MuxN.scala 16:10:@103057.4]
  assign io_out_wdata_8 = io_sel ? io_ins_1_wdata_8 : 8'h0; // @[MuxN.scala 16:10:@103058.4]
  assign io_out_wdata_9 = io_sel ? io_ins_1_wdata_9 : 8'h0; // @[MuxN.scala 16:10:@103059.4]
  assign io_out_wdata_10 = io_sel ? io_ins_1_wdata_10 : 8'h0; // @[MuxN.scala 16:10:@103060.4]
  assign io_out_wdata_11 = io_sel ? io_ins_1_wdata_11 : 8'h0; // @[MuxN.scala 16:10:@103061.4]
  assign io_out_wdata_12 = io_sel ? io_ins_1_wdata_12 : 8'h0; // @[MuxN.scala 16:10:@103062.4]
  assign io_out_wdata_13 = io_sel ? io_ins_1_wdata_13 : 8'h0; // @[MuxN.scala 16:10:@103063.4]
  assign io_out_wdata_14 = io_sel ? io_ins_1_wdata_14 : 8'h0; // @[MuxN.scala 16:10:@103064.4]
  assign io_out_wdata_15 = io_sel ? io_ins_1_wdata_15 : 8'h0; // @[MuxN.scala 16:10:@103065.4]
  assign io_out_wdata_16 = io_sel ? io_ins_1_wdata_16 : 8'h0; // @[MuxN.scala 16:10:@103066.4]
  assign io_out_wdata_17 = io_sel ? io_ins_1_wdata_17 : 8'h0; // @[MuxN.scala 16:10:@103067.4]
  assign io_out_wdata_18 = io_sel ? io_ins_1_wdata_18 : 8'h0; // @[MuxN.scala 16:10:@103068.4]
  assign io_out_wdata_19 = io_sel ? io_ins_1_wdata_19 : 8'h0; // @[MuxN.scala 16:10:@103069.4]
  assign io_out_wdata_20 = io_sel ? io_ins_1_wdata_20 : 8'h0; // @[MuxN.scala 16:10:@103070.4]
  assign io_out_wdata_21 = io_sel ? io_ins_1_wdata_21 : 8'h0; // @[MuxN.scala 16:10:@103071.4]
  assign io_out_wdata_22 = io_sel ? io_ins_1_wdata_22 : 8'h0; // @[MuxN.scala 16:10:@103072.4]
  assign io_out_wdata_23 = io_sel ? io_ins_1_wdata_23 : 8'h0; // @[MuxN.scala 16:10:@103073.4]
  assign io_out_wdata_24 = io_sel ? io_ins_1_wdata_24 : 8'h0; // @[MuxN.scala 16:10:@103074.4]
  assign io_out_wdata_25 = io_sel ? io_ins_1_wdata_25 : 8'h0; // @[MuxN.scala 16:10:@103075.4]
  assign io_out_wdata_26 = io_sel ? io_ins_1_wdata_26 : 8'h0; // @[MuxN.scala 16:10:@103076.4]
  assign io_out_wdata_27 = io_sel ? io_ins_1_wdata_27 : 8'h0; // @[MuxN.scala 16:10:@103077.4]
  assign io_out_wdata_28 = io_sel ? io_ins_1_wdata_28 : 8'h0; // @[MuxN.scala 16:10:@103078.4]
  assign io_out_wdata_29 = io_sel ? io_ins_1_wdata_29 : 8'h0; // @[MuxN.scala 16:10:@103079.4]
  assign io_out_wdata_30 = io_sel ? io_ins_1_wdata_30 : 8'h0; // @[MuxN.scala 16:10:@103080.4]
  assign io_out_wdata_31 = io_sel ? io_ins_1_wdata_31 : 8'h0; // @[MuxN.scala 16:10:@103081.4]
  assign io_out_wdata_32 = io_sel ? io_ins_1_wdata_32 : 8'h0; // @[MuxN.scala 16:10:@103082.4]
  assign io_out_wdata_33 = io_sel ? io_ins_1_wdata_33 : 8'h0; // @[MuxN.scala 16:10:@103083.4]
  assign io_out_wdata_34 = io_sel ? io_ins_1_wdata_34 : 8'h0; // @[MuxN.scala 16:10:@103084.4]
  assign io_out_wdata_35 = io_sel ? io_ins_1_wdata_35 : 8'h0; // @[MuxN.scala 16:10:@103085.4]
  assign io_out_wdata_36 = io_sel ? io_ins_1_wdata_36 : 8'h0; // @[MuxN.scala 16:10:@103086.4]
  assign io_out_wdata_37 = io_sel ? io_ins_1_wdata_37 : 8'h0; // @[MuxN.scala 16:10:@103087.4]
  assign io_out_wdata_38 = io_sel ? io_ins_1_wdata_38 : 8'h0; // @[MuxN.scala 16:10:@103088.4]
  assign io_out_wdata_39 = io_sel ? io_ins_1_wdata_39 : 8'h0; // @[MuxN.scala 16:10:@103089.4]
  assign io_out_wdata_40 = io_sel ? io_ins_1_wdata_40 : 8'h0; // @[MuxN.scala 16:10:@103090.4]
  assign io_out_wdata_41 = io_sel ? io_ins_1_wdata_41 : 8'h0; // @[MuxN.scala 16:10:@103091.4]
  assign io_out_wdata_42 = io_sel ? io_ins_1_wdata_42 : 8'h0; // @[MuxN.scala 16:10:@103092.4]
  assign io_out_wdata_43 = io_sel ? io_ins_1_wdata_43 : 8'h0; // @[MuxN.scala 16:10:@103093.4]
  assign io_out_wdata_44 = io_sel ? io_ins_1_wdata_44 : 8'h0; // @[MuxN.scala 16:10:@103094.4]
  assign io_out_wdata_45 = io_sel ? io_ins_1_wdata_45 : 8'h0; // @[MuxN.scala 16:10:@103095.4]
  assign io_out_wdata_46 = io_sel ? io_ins_1_wdata_46 : 8'h0; // @[MuxN.scala 16:10:@103096.4]
  assign io_out_wdata_47 = io_sel ? io_ins_1_wdata_47 : 8'h0; // @[MuxN.scala 16:10:@103097.4]
  assign io_out_wdata_48 = io_sel ? io_ins_1_wdata_48 : 8'h0; // @[MuxN.scala 16:10:@103098.4]
  assign io_out_wdata_49 = io_sel ? io_ins_1_wdata_49 : 8'h0; // @[MuxN.scala 16:10:@103099.4]
  assign io_out_wdata_50 = io_sel ? io_ins_1_wdata_50 : 8'h0; // @[MuxN.scala 16:10:@103100.4]
  assign io_out_wdata_51 = io_sel ? io_ins_1_wdata_51 : 8'h0; // @[MuxN.scala 16:10:@103101.4]
  assign io_out_wdata_52 = io_sel ? io_ins_1_wdata_52 : 8'h0; // @[MuxN.scala 16:10:@103102.4]
  assign io_out_wdata_53 = io_sel ? io_ins_1_wdata_53 : 8'h0; // @[MuxN.scala 16:10:@103103.4]
  assign io_out_wdata_54 = io_sel ? io_ins_1_wdata_54 : 8'h0; // @[MuxN.scala 16:10:@103104.4]
  assign io_out_wdata_55 = io_sel ? io_ins_1_wdata_55 : 8'h0; // @[MuxN.scala 16:10:@103105.4]
  assign io_out_wdata_56 = io_sel ? io_ins_1_wdata_56 : 8'h0; // @[MuxN.scala 16:10:@103106.4]
  assign io_out_wdata_57 = io_sel ? io_ins_1_wdata_57 : 8'h0; // @[MuxN.scala 16:10:@103107.4]
  assign io_out_wdata_58 = io_sel ? io_ins_1_wdata_58 : 8'h0; // @[MuxN.scala 16:10:@103108.4]
  assign io_out_wdata_59 = io_sel ? io_ins_1_wdata_59 : 8'h0; // @[MuxN.scala 16:10:@103109.4]
  assign io_out_wdata_60 = io_sel ? io_ins_1_wdata_60 : 8'h0; // @[MuxN.scala 16:10:@103110.4]
  assign io_out_wdata_61 = io_sel ? io_ins_1_wdata_61 : 8'h0; // @[MuxN.scala 16:10:@103111.4]
  assign io_out_wdata_62 = io_sel ? io_ins_1_wdata_62 : 8'h0; // @[MuxN.scala 16:10:@103112.4]
  assign io_out_wdata_63 = io_sel ? io_ins_1_wdata_63 : 8'h0; // @[MuxN.scala 16:10:@103113.4]
  assign io_out_wstrb_0 = io_sel ? io_ins_1_wstrb_0 : 1'h0; // @[MuxN.scala 16:10:@102986.4]
  assign io_out_wstrb_1 = io_sel ? io_ins_1_wstrb_1 : 1'h0; // @[MuxN.scala 16:10:@102987.4]
  assign io_out_wstrb_2 = io_sel ? io_ins_1_wstrb_2 : 1'h0; // @[MuxN.scala 16:10:@102988.4]
  assign io_out_wstrb_3 = io_sel ? io_ins_1_wstrb_3 : 1'h0; // @[MuxN.scala 16:10:@102989.4]
  assign io_out_wstrb_4 = io_sel ? io_ins_1_wstrb_4 : 1'h0; // @[MuxN.scala 16:10:@102990.4]
  assign io_out_wstrb_5 = io_sel ? io_ins_1_wstrb_5 : 1'h0; // @[MuxN.scala 16:10:@102991.4]
  assign io_out_wstrb_6 = io_sel ? io_ins_1_wstrb_6 : 1'h0; // @[MuxN.scala 16:10:@102992.4]
  assign io_out_wstrb_7 = io_sel ? io_ins_1_wstrb_7 : 1'h0; // @[MuxN.scala 16:10:@102993.4]
  assign io_out_wstrb_8 = io_sel ? io_ins_1_wstrb_8 : 1'h0; // @[MuxN.scala 16:10:@102994.4]
  assign io_out_wstrb_9 = io_sel ? io_ins_1_wstrb_9 : 1'h0; // @[MuxN.scala 16:10:@102995.4]
  assign io_out_wstrb_10 = io_sel ? io_ins_1_wstrb_10 : 1'h0; // @[MuxN.scala 16:10:@102996.4]
  assign io_out_wstrb_11 = io_sel ? io_ins_1_wstrb_11 : 1'h0; // @[MuxN.scala 16:10:@102997.4]
  assign io_out_wstrb_12 = io_sel ? io_ins_1_wstrb_12 : 1'h0; // @[MuxN.scala 16:10:@102998.4]
  assign io_out_wstrb_13 = io_sel ? io_ins_1_wstrb_13 : 1'h0; // @[MuxN.scala 16:10:@102999.4]
  assign io_out_wstrb_14 = io_sel ? io_ins_1_wstrb_14 : 1'h0; // @[MuxN.scala 16:10:@103000.4]
  assign io_out_wstrb_15 = io_sel ? io_ins_1_wstrb_15 : 1'h0; // @[MuxN.scala 16:10:@103001.4]
  assign io_out_wstrb_16 = io_sel ? io_ins_1_wstrb_16 : 1'h0; // @[MuxN.scala 16:10:@103002.4]
  assign io_out_wstrb_17 = io_sel ? io_ins_1_wstrb_17 : 1'h0; // @[MuxN.scala 16:10:@103003.4]
  assign io_out_wstrb_18 = io_sel ? io_ins_1_wstrb_18 : 1'h0; // @[MuxN.scala 16:10:@103004.4]
  assign io_out_wstrb_19 = io_sel ? io_ins_1_wstrb_19 : 1'h0; // @[MuxN.scala 16:10:@103005.4]
  assign io_out_wstrb_20 = io_sel ? io_ins_1_wstrb_20 : 1'h0; // @[MuxN.scala 16:10:@103006.4]
  assign io_out_wstrb_21 = io_sel ? io_ins_1_wstrb_21 : 1'h0; // @[MuxN.scala 16:10:@103007.4]
  assign io_out_wstrb_22 = io_sel ? io_ins_1_wstrb_22 : 1'h0; // @[MuxN.scala 16:10:@103008.4]
  assign io_out_wstrb_23 = io_sel ? io_ins_1_wstrb_23 : 1'h0; // @[MuxN.scala 16:10:@103009.4]
  assign io_out_wstrb_24 = io_sel ? io_ins_1_wstrb_24 : 1'h0; // @[MuxN.scala 16:10:@103010.4]
  assign io_out_wstrb_25 = io_sel ? io_ins_1_wstrb_25 : 1'h0; // @[MuxN.scala 16:10:@103011.4]
  assign io_out_wstrb_26 = io_sel ? io_ins_1_wstrb_26 : 1'h0; // @[MuxN.scala 16:10:@103012.4]
  assign io_out_wstrb_27 = io_sel ? io_ins_1_wstrb_27 : 1'h0; // @[MuxN.scala 16:10:@103013.4]
  assign io_out_wstrb_28 = io_sel ? io_ins_1_wstrb_28 : 1'h0; // @[MuxN.scala 16:10:@103014.4]
  assign io_out_wstrb_29 = io_sel ? io_ins_1_wstrb_29 : 1'h0; // @[MuxN.scala 16:10:@103015.4]
  assign io_out_wstrb_30 = io_sel ? io_ins_1_wstrb_30 : 1'h0; // @[MuxN.scala 16:10:@103016.4]
  assign io_out_wstrb_31 = io_sel ? io_ins_1_wstrb_31 : 1'h0; // @[MuxN.scala 16:10:@103017.4]
  assign io_out_wstrb_32 = io_sel ? io_ins_1_wstrb_32 : 1'h0; // @[MuxN.scala 16:10:@103018.4]
  assign io_out_wstrb_33 = io_sel ? io_ins_1_wstrb_33 : 1'h0; // @[MuxN.scala 16:10:@103019.4]
  assign io_out_wstrb_34 = io_sel ? io_ins_1_wstrb_34 : 1'h0; // @[MuxN.scala 16:10:@103020.4]
  assign io_out_wstrb_35 = io_sel ? io_ins_1_wstrb_35 : 1'h0; // @[MuxN.scala 16:10:@103021.4]
  assign io_out_wstrb_36 = io_sel ? io_ins_1_wstrb_36 : 1'h0; // @[MuxN.scala 16:10:@103022.4]
  assign io_out_wstrb_37 = io_sel ? io_ins_1_wstrb_37 : 1'h0; // @[MuxN.scala 16:10:@103023.4]
  assign io_out_wstrb_38 = io_sel ? io_ins_1_wstrb_38 : 1'h0; // @[MuxN.scala 16:10:@103024.4]
  assign io_out_wstrb_39 = io_sel ? io_ins_1_wstrb_39 : 1'h0; // @[MuxN.scala 16:10:@103025.4]
  assign io_out_wstrb_40 = io_sel ? io_ins_1_wstrb_40 : 1'h0; // @[MuxN.scala 16:10:@103026.4]
  assign io_out_wstrb_41 = io_sel ? io_ins_1_wstrb_41 : 1'h0; // @[MuxN.scala 16:10:@103027.4]
  assign io_out_wstrb_42 = io_sel ? io_ins_1_wstrb_42 : 1'h0; // @[MuxN.scala 16:10:@103028.4]
  assign io_out_wstrb_43 = io_sel ? io_ins_1_wstrb_43 : 1'h0; // @[MuxN.scala 16:10:@103029.4]
  assign io_out_wstrb_44 = io_sel ? io_ins_1_wstrb_44 : 1'h0; // @[MuxN.scala 16:10:@103030.4]
  assign io_out_wstrb_45 = io_sel ? io_ins_1_wstrb_45 : 1'h0; // @[MuxN.scala 16:10:@103031.4]
  assign io_out_wstrb_46 = io_sel ? io_ins_1_wstrb_46 : 1'h0; // @[MuxN.scala 16:10:@103032.4]
  assign io_out_wstrb_47 = io_sel ? io_ins_1_wstrb_47 : 1'h0; // @[MuxN.scala 16:10:@103033.4]
  assign io_out_wstrb_48 = io_sel ? io_ins_1_wstrb_48 : 1'h0; // @[MuxN.scala 16:10:@103034.4]
  assign io_out_wstrb_49 = io_sel ? io_ins_1_wstrb_49 : 1'h0; // @[MuxN.scala 16:10:@103035.4]
  assign io_out_wstrb_50 = io_sel ? io_ins_1_wstrb_50 : 1'h0; // @[MuxN.scala 16:10:@103036.4]
  assign io_out_wstrb_51 = io_sel ? io_ins_1_wstrb_51 : 1'h0; // @[MuxN.scala 16:10:@103037.4]
  assign io_out_wstrb_52 = io_sel ? io_ins_1_wstrb_52 : 1'h0; // @[MuxN.scala 16:10:@103038.4]
  assign io_out_wstrb_53 = io_sel ? io_ins_1_wstrb_53 : 1'h0; // @[MuxN.scala 16:10:@103039.4]
  assign io_out_wstrb_54 = io_sel ? io_ins_1_wstrb_54 : 1'h0; // @[MuxN.scala 16:10:@103040.4]
  assign io_out_wstrb_55 = io_sel ? io_ins_1_wstrb_55 : 1'h0; // @[MuxN.scala 16:10:@103041.4]
  assign io_out_wstrb_56 = io_sel ? io_ins_1_wstrb_56 : 1'h0; // @[MuxN.scala 16:10:@103042.4]
  assign io_out_wstrb_57 = io_sel ? io_ins_1_wstrb_57 : 1'h0; // @[MuxN.scala 16:10:@103043.4]
  assign io_out_wstrb_58 = io_sel ? io_ins_1_wstrb_58 : 1'h0; // @[MuxN.scala 16:10:@103044.4]
  assign io_out_wstrb_59 = io_sel ? io_ins_1_wstrb_59 : 1'h0; // @[MuxN.scala 16:10:@103045.4]
  assign io_out_wstrb_60 = io_sel ? io_ins_1_wstrb_60 : 1'h0; // @[MuxN.scala 16:10:@103046.4]
  assign io_out_wstrb_61 = io_sel ? io_ins_1_wstrb_61 : 1'h0; // @[MuxN.scala 16:10:@103047.4]
  assign io_out_wstrb_62 = io_sel ? io_ins_1_wstrb_62 : 1'h0; // @[MuxN.scala 16:10:@103048.4]
  assign io_out_wstrb_63 = io_sel ? io_ins_1_wstrb_63 : 1'h0; // @[MuxN.scala 16:10:@103049.4]
endmodule
module MuxPipe_1( // @[:@103115.2]
  output       io_in_ready, // @[:@103118.4]
  input        io_in_valid, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_0, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_1, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_2, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_3, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_4, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_5, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_6, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_7, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_8, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_9, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_10, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_11, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_12, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_13, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_14, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_15, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_16, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_17, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_18, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_19, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_20, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_21, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_22, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_23, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_24, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_25, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_26, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_27, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_28, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_29, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_30, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_31, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_32, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_33, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_34, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_35, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_36, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_37, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_38, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_39, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_40, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_41, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_42, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_43, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_44, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_45, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_46, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_47, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_48, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_49, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_50, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_51, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_52, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_53, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_54, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_55, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_56, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_57, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_58, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_59, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_60, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_61, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_62, // @[:@103118.4]
  input  [7:0] io_in_bits_1_wdata_63, // @[:@103118.4]
  input        io_in_bits_1_wstrb_0, // @[:@103118.4]
  input        io_in_bits_1_wstrb_1, // @[:@103118.4]
  input        io_in_bits_1_wstrb_2, // @[:@103118.4]
  input        io_in_bits_1_wstrb_3, // @[:@103118.4]
  input        io_in_bits_1_wstrb_4, // @[:@103118.4]
  input        io_in_bits_1_wstrb_5, // @[:@103118.4]
  input        io_in_bits_1_wstrb_6, // @[:@103118.4]
  input        io_in_bits_1_wstrb_7, // @[:@103118.4]
  input        io_in_bits_1_wstrb_8, // @[:@103118.4]
  input        io_in_bits_1_wstrb_9, // @[:@103118.4]
  input        io_in_bits_1_wstrb_10, // @[:@103118.4]
  input        io_in_bits_1_wstrb_11, // @[:@103118.4]
  input        io_in_bits_1_wstrb_12, // @[:@103118.4]
  input        io_in_bits_1_wstrb_13, // @[:@103118.4]
  input        io_in_bits_1_wstrb_14, // @[:@103118.4]
  input        io_in_bits_1_wstrb_15, // @[:@103118.4]
  input        io_in_bits_1_wstrb_16, // @[:@103118.4]
  input        io_in_bits_1_wstrb_17, // @[:@103118.4]
  input        io_in_bits_1_wstrb_18, // @[:@103118.4]
  input        io_in_bits_1_wstrb_19, // @[:@103118.4]
  input        io_in_bits_1_wstrb_20, // @[:@103118.4]
  input        io_in_bits_1_wstrb_21, // @[:@103118.4]
  input        io_in_bits_1_wstrb_22, // @[:@103118.4]
  input        io_in_bits_1_wstrb_23, // @[:@103118.4]
  input        io_in_bits_1_wstrb_24, // @[:@103118.4]
  input        io_in_bits_1_wstrb_25, // @[:@103118.4]
  input        io_in_bits_1_wstrb_26, // @[:@103118.4]
  input        io_in_bits_1_wstrb_27, // @[:@103118.4]
  input        io_in_bits_1_wstrb_28, // @[:@103118.4]
  input        io_in_bits_1_wstrb_29, // @[:@103118.4]
  input        io_in_bits_1_wstrb_30, // @[:@103118.4]
  input        io_in_bits_1_wstrb_31, // @[:@103118.4]
  input        io_in_bits_1_wstrb_32, // @[:@103118.4]
  input        io_in_bits_1_wstrb_33, // @[:@103118.4]
  input        io_in_bits_1_wstrb_34, // @[:@103118.4]
  input        io_in_bits_1_wstrb_35, // @[:@103118.4]
  input        io_in_bits_1_wstrb_36, // @[:@103118.4]
  input        io_in_bits_1_wstrb_37, // @[:@103118.4]
  input        io_in_bits_1_wstrb_38, // @[:@103118.4]
  input        io_in_bits_1_wstrb_39, // @[:@103118.4]
  input        io_in_bits_1_wstrb_40, // @[:@103118.4]
  input        io_in_bits_1_wstrb_41, // @[:@103118.4]
  input        io_in_bits_1_wstrb_42, // @[:@103118.4]
  input        io_in_bits_1_wstrb_43, // @[:@103118.4]
  input        io_in_bits_1_wstrb_44, // @[:@103118.4]
  input        io_in_bits_1_wstrb_45, // @[:@103118.4]
  input        io_in_bits_1_wstrb_46, // @[:@103118.4]
  input        io_in_bits_1_wstrb_47, // @[:@103118.4]
  input        io_in_bits_1_wstrb_48, // @[:@103118.4]
  input        io_in_bits_1_wstrb_49, // @[:@103118.4]
  input        io_in_bits_1_wstrb_50, // @[:@103118.4]
  input        io_in_bits_1_wstrb_51, // @[:@103118.4]
  input        io_in_bits_1_wstrb_52, // @[:@103118.4]
  input        io_in_bits_1_wstrb_53, // @[:@103118.4]
  input        io_in_bits_1_wstrb_54, // @[:@103118.4]
  input        io_in_bits_1_wstrb_55, // @[:@103118.4]
  input        io_in_bits_1_wstrb_56, // @[:@103118.4]
  input        io_in_bits_1_wstrb_57, // @[:@103118.4]
  input        io_in_bits_1_wstrb_58, // @[:@103118.4]
  input        io_in_bits_1_wstrb_59, // @[:@103118.4]
  input        io_in_bits_1_wstrb_60, // @[:@103118.4]
  input        io_in_bits_1_wstrb_61, // @[:@103118.4]
  input        io_in_bits_1_wstrb_62, // @[:@103118.4]
  input        io_in_bits_1_wstrb_63, // @[:@103118.4]
  input        io_sel, // @[:@103118.4]
  input        io_out_ready, // @[:@103118.4]
  output       io_out_valid, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_0, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_1, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_2, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_3, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_4, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_5, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_6, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_7, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_8, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_9, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_10, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_11, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_12, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_13, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_14, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_15, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_16, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_17, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_18, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_19, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_20, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_21, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_22, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_23, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_24, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_25, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_26, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_27, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_28, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_29, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_30, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_31, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_32, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_33, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_34, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_35, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_36, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_37, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_38, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_39, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_40, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_41, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_42, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_43, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_44, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_45, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_46, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_47, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_48, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_49, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_50, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_51, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_52, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_53, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_54, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_55, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_56, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_57, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_58, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_59, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_60, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_61, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_62, // @[:@103118.4]
  output [7:0] io_out_bits_wdata_63, // @[:@103118.4]
  output       io_out_bits_wstrb_0, // @[:@103118.4]
  output       io_out_bits_wstrb_1, // @[:@103118.4]
  output       io_out_bits_wstrb_2, // @[:@103118.4]
  output       io_out_bits_wstrb_3, // @[:@103118.4]
  output       io_out_bits_wstrb_4, // @[:@103118.4]
  output       io_out_bits_wstrb_5, // @[:@103118.4]
  output       io_out_bits_wstrb_6, // @[:@103118.4]
  output       io_out_bits_wstrb_7, // @[:@103118.4]
  output       io_out_bits_wstrb_8, // @[:@103118.4]
  output       io_out_bits_wstrb_9, // @[:@103118.4]
  output       io_out_bits_wstrb_10, // @[:@103118.4]
  output       io_out_bits_wstrb_11, // @[:@103118.4]
  output       io_out_bits_wstrb_12, // @[:@103118.4]
  output       io_out_bits_wstrb_13, // @[:@103118.4]
  output       io_out_bits_wstrb_14, // @[:@103118.4]
  output       io_out_bits_wstrb_15, // @[:@103118.4]
  output       io_out_bits_wstrb_16, // @[:@103118.4]
  output       io_out_bits_wstrb_17, // @[:@103118.4]
  output       io_out_bits_wstrb_18, // @[:@103118.4]
  output       io_out_bits_wstrb_19, // @[:@103118.4]
  output       io_out_bits_wstrb_20, // @[:@103118.4]
  output       io_out_bits_wstrb_21, // @[:@103118.4]
  output       io_out_bits_wstrb_22, // @[:@103118.4]
  output       io_out_bits_wstrb_23, // @[:@103118.4]
  output       io_out_bits_wstrb_24, // @[:@103118.4]
  output       io_out_bits_wstrb_25, // @[:@103118.4]
  output       io_out_bits_wstrb_26, // @[:@103118.4]
  output       io_out_bits_wstrb_27, // @[:@103118.4]
  output       io_out_bits_wstrb_28, // @[:@103118.4]
  output       io_out_bits_wstrb_29, // @[:@103118.4]
  output       io_out_bits_wstrb_30, // @[:@103118.4]
  output       io_out_bits_wstrb_31, // @[:@103118.4]
  output       io_out_bits_wstrb_32, // @[:@103118.4]
  output       io_out_bits_wstrb_33, // @[:@103118.4]
  output       io_out_bits_wstrb_34, // @[:@103118.4]
  output       io_out_bits_wstrb_35, // @[:@103118.4]
  output       io_out_bits_wstrb_36, // @[:@103118.4]
  output       io_out_bits_wstrb_37, // @[:@103118.4]
  output       io_out_bits_wstrb_38, // @[:@103118.4]
  output       io_out_bits_wstrb_39, // @[:@103118.4]
  output       io_out_bits_wstrb_40, // @[:@103118.4]
  output       io_out_bits_wstrb_41, // @[:@103118.4]
  output       io_out_bits_wstrb_42, // @[:@103118.4]
  output       io_out_bits_wstrb_43, // @[:@103118.4]
  output       io_out_bits_wstrb_44, // @[:@103118.4]
  output       io_out_bits_wstrb_45, // @[:@103118.4]
  output       io_out_bits_wstrb_46, // @[:@103118.4]
  output       io_out_bits_wstrb_47, // @[:@103118.4]
  output       io_out_bits_wstrb_48, // @[:@103118.4]
  output       io_out_bits_wstrb_49, // @[:@103118.4]
  output       io_out_bits_wstrb_50, // @[:@103118.4]
  output       io_out_bits_wstrb_51, // @[:@103118.4]
  output       io_out_bits_wstrb_52, // @[:@103118.4]
  output       io_out_bits_wstrb_53, // @[:@103118.4]
  output       io_out_bits_wstrb_54, // @[:@103118.4]
  output       io_out_bits_wstrb_55, // @[:@103118.4]
  output       io_out_bits_wstrb_56, // @[:@103118.4]
  output       io_out_bits_wstrb_57, // @[:@103118.4]
  output       io_out_bits_wstrb_58, // @[:@103118.4]
  output       io_out_bits_wstrb_59, // @[:@103118.4]
  output       io_out_bits_wstrb_60, // @[:@103118.4]
  output       io_out_bits_wstrb_61, // @[:@103118.4]
  output       io_out_bits_wstrb_62, // @[:@103118.4]
  output       io_out_bits_wstrb_63 // @[:@103118.4]
);
  wire [7:0] MuxN_io_ins_1_wdata_0; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_1; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_2; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_3; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_4; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_5; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_6; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_7; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_8; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_9; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_10; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_11; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_12; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_13; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_14; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_15; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_16; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_17; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_18; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_19; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_20; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_21; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_22; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_23; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_24; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_25; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_26; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_27; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_28; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_29; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_30; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_31; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_32; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_33; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_34; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_35; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_36; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_37; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_38; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_39; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_40; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_41; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_42; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_43; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_44; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_45; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_46; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_47; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_48; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_49; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_50; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_51; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_52; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_53; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_54; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_55; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_56; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_57; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_58; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_59; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_60; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_61; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_62; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_ins_1_wdata_63; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_0; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_1; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_2; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_3; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_4; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_5; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_6; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_7; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_8; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_9; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_10; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_11; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_12; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_13; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_14; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_15; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_16; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_17; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_18; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_19; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_20; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_21; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_22; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_23; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_24; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_25; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_26; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_27; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_28; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_29; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_30; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_31; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_32; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_33; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_34; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_35; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_36; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_37; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_38; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_39; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_40; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_41; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_42; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_43; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_44; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_45; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_46; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_47; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_48; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_49; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_50; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_51; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_52; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_53; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_54; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_55; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_56; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_57; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_58; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_59; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_60; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_61; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_62; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_ins_1_wstrb_63; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_sel; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_0; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_1; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_2; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_3; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_4; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_5; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_6; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_7; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_8; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_9; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_10; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_11; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_12; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_13; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_14; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_15; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_16; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_17; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_18; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_19; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_20; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_21; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_22; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_23; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_24; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_25; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_26; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_27; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_28; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_29; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_30; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_31; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_32; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_33; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_34; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_35; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_36; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_37; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_38; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_39; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_40; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_41; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_42; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_43; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_44; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_45; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_46; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_47; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_48; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_49; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_50; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_51; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_52; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_53; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_54; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_55; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_56; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_57; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_58; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_59; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_60; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_61; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_62; // @[MuxN.scala 40:23:@103381.4]
  wire [7:0] MuxN_io_out_wdata_63; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_0; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_1; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_2; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_3; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_4; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_5; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_6; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_7; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_8; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_9; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_10; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_11; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_12; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_13; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_14; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_15; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_16; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_17; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_18; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_19; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_20; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_21; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_22; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_23; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_24; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_25; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_26; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_27; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_28; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_29; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_30; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_31; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_32; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_33; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_34; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_35; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_36; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_37; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_38; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_39; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_40; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_41; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_42; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_43; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_44; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_45; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_46; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_47; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_48; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_49; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_50; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_51; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_52; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_53; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_54; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_55; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_56; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_57; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_58; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_59; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_60; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_61; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_62; // @[MuxN.scala 40:23:@103381.4]
  wire  MuxN_io_out_wstrb_63; // @[MuxN.scala 40:23:@103381.4]
  wire  _T_190; // @[MuxN.scala 28:31:@103120.4]
  MuxN_1 MuxN ( // @[MuxN.scala 40:23:@103381.4]
    .io_ins_1_wdata_0(MuxN_io_ins_1_wdata_0),
    .io_ins_1_wdata_1(MuxN_io_ins_1_wdata_1),
    .io_ins_1_wdata_2(MuxN_io_ins_1_wdata_2),
    .io_ins_1_wdata_3(MuxN_io_ins_1_wdata_3),
    .io_ins_1_wdata_4(MuxN_io_ins_1_wdata_4),
    .io_ins_1_wdata_5(MuxN_io_ins_1_wdata_5),
    .io_ins_1_wdata_6(MuxN_io_ins_1_wdata_6),
    .io_ins_1_wdata_7(MuxN_io_ins_1_wdata_7),
    .io_ins_1_wdata_8(MuxN_io_ins_1_wdata_8),
    .io_ins_1_wdata_9(MuxN_io_ins_1_wdata_9),
    .io_ins_1_wdata_10(MuxN_io_ins_1_wdata_10),
    .io_ins_1_wdata_11(MuxN_io_ins_1_wdata_11),
    .io_ins_1_wdata_12(MuxN_io_ins_1_wdata_12),
    .io_ins_1_wdata_13(MuxN_io_ins_1_wdata_13),
    .io_ins_1_wdata_14(MuxN_io_ins_1_wdata_14),
    .io_ins_1_wdata_15(MuxN_io_ins_1_wdata_15),
    .io_ins_1_wdata_16(MuxN_io_ins_1_wdata_16),
    .io_ins_1_wdata_17(MuxN_io_ins_1_wdata_17),
    .io_ins_1_wdata_18(MuxN_io_ins_1_wdata_18),
    .io_ins_1_wdata_19(MuxN_io_ins_1_wdata_19),
    .io_ins_1_wdata_20(MuxN_io_ins_1_wdata_20),
    .io_ins_1_wdata_21(MuxN_io_ins_1_wdata_21),
    .io_ins_1_wdata_22(MuxN_io_ins_1_wdata_22),
    .io_ins_1_wdata_23(MuxN_io_ins_1_wdata_23),
    .io_ins_1_wdata_24(MuxN_io_ins_1_wdata_24),
    .io_ins_1_wdata_25(MuxN_io_ins_1_wdata_25),
    .io_ins_1_wdata_26(MuxN_io_ins_1_wdata_26),
    .io_ins_1_wdata_27(MuxN_io_ins_1_wdata_27),
    .io_ins_1_wdata_28(MuxN_io_ins_1_wdata_28),
    .io_ins_1_wdata_29(MuxN_io_ins_1_wdata_29),
    .io_ins_1_wdata_30(MuxN_io_ins_1_wdata_30),
    .io_ins_1_wdata_31(MuxN_io_ins_1_wdata_31),
    .io_ins_1_wdata_32(MuxN_io_ins_1_wdata_32),
    .io_ins_1_wdata_33(MuxN_io_ins_1_wdata_33),
    .io_ins_1_wdata_34(MuxN_io_ins_1_wdata_34),
    .io_ins_1_wdata_35(MuxN_io_ins_1_wdata_35),
    .io_ins_1_wdata_36(MuxN_io_ins_1_wdata_36),
    .io_ins_1_wdata_37(MuxN_io_ins_1_wdata_37),
    .io_ins_1_wdata_38(MuxN_io_ins_1_wdata_38),
    .io_ins_1_wdata_39(MuxN_io_ins_1_wdata_39),
    .io_ins_1_wdata_40(MuxN_io_ins_1_wdata_40),
    .io_ins_1_wdata_41(MuxN_io_ins_1_wdata_41),
    .io_ins_1_wdata_42(MuxN_io_ins_1_wdata_42),
    .io_ins_1_wdata_43(MuxN_io_ins_1_wdata_43),
    .io_ins_1_wdata_44(MuxN_io_ins_1_wdata_44),
    .io_ins_1_wdata_45(MuxN_io_ins_1_wdata_45),
    .io_ins_1_wdata_46(MuxN_io_ins_1_wdata_46),
    .io_ins_1_wdata_47(MuxN_io_ins_1_wdata_47),
    .io_ins_1_wdata_48(MuxN_io_ins_1_wdata_48),
    .io_ins_1_wdata_49(MuxN_io_ins_1_wdata_49),
    .io_ins_1_wdata_50(MuxN_io_ins_1_wdata_50),
    .io_ins_1_wdata_51(MuxN_io_ins_1_wdata_51),
    .io_ins_1_wdata_52(MuxN_io_ins_1_wdata_52),
    .io_ins_1_wdata_53(MuxN_io_ins_1_wdata_53),
    .io_ins_1_wdata_54(MuxN_io_ins_1_wdata_54),
    .io_ins_1_wdata_55(MuxN_io_ins_1_wdata_55),
    .io_ins_1_wdata_56(MuxN_io_ins_1_wdata_56),
    .io_ins_1_wdata_57(MuxN_io_ins_1_wdata_57),
    .io_ins_1_wdata_58(MuxN_io_ins_1_wdata_58),
    .io_ins_1_wdata_59(MuxN_io_ins_1_wdata_59),
    .io_ins_1_wdata_60(MuxN_io_ins_1_wdata_60),
    .io_ins_1_wdata_61(MuxN_io_ins_1_wdata_61),
    .io_ins_1_wdata_62(MuxN_io_ins_1_wdata_62),
    .io_ins_1_wdata_63(MuxN_io_ins_1_wdata_63),
    .io_ins_1_wstrb_0(MuxN_io_ins_1_wstrb_0),
    .io_ins_1_wstrb_1(MuxN_io_ins_1_wstrb_1),
    .io_ins_1_wstrb_2(MuxN_io_ins_1_wstrb_2),
    .io_ins_1_wstrb_3(MuxN_io_ins_1_wstrb_3),
    .io_ins_1_wstrb_4(MuxN_io_ins_1_wstrb_4),
    .io_ins_1_wstrb_5(MuxN_io_ins_1_wstrb_5),
    .io_ins_1_wstrb_6(MuxN_io_ins_1_wstrb_6),
    .io_ins_1_wstrb_7(MuxN_io_ins_1_wstrb_7),
    .io_ins_1_wstrb_8(MuxN_io_ins_1_wstrb_8),
    .io_ins_1_wstrb_9(MuxN_io_ins_1_wstrb_9),
    .io_ins_1_wstrb_10(MuxN_io_ins_1_wstrb_10),
    .io_ins_1_wstrb_11(MuxN_io_ins_1_wstrb_11),
    .io_ins_1_wstrb_12(MuxN_io_ins_1_wstrb_12),
    .io_ins_1_wstrb_13(MuxN_io_ins_1_wstrb_13),
    .io_ins_1_wstrb_14(MuxN_io_ins_1_wstrb_14),
    .io_ins_1_wstrb_15(MuxN_io_ins_1_wstrb_15),
    .io_ins_1_wstrb_16(MuxN_io_ins_1_wstrb_16),
    .io_ins_1_wstrb_17(MuxN_io_ins_1_wstrb_17),
    .io_ins_1_wstrb_18(MuxN_io_ins_1_wstrb_18),
    .io_ins_1_wstrb_19(MuxN_io_ins_1_wstrb_19),
    .io_ins_1_wstrb_20(MuxN_io_ins_1_wstrb_20),
    .io_ins_1_wstrb_21(MuxN_io_ins_1_wstrb_21),
    .io_ins_1_wstrb_22(MuxN_io_ins_1_wstrb_22),
    .io_ins_1_wstrb_23(MuxN_io_ins_1_wstrb_23),
    .io_ins_1_wstrb_24(MuxN_io_ins_1_wstrb_24),
    .io_ins_1_wstrb_25(MuxN_io_ins_1_wstrb_25),
    .io_ins_1_wstrb_26(MuxN_io_ins_1_wstrb_26),
    .io_ins_1_wstrb_27(MuxN_io_ins_1_wstrb_27),
    .io_ins_1_wstrb_28(MuxN_io_ins_1_wstrb_28),
    .io_ins_1_wstrb_29(MuxN_io_ins_1_wstrb_29),
    .io_ins_1_wstrb_30(MuxN_io_ins_1_wstrb_30),
    .io_ins_1_wstrb_31(MuxN_io_ins_1_wstrb_31),
    .io_ins_1_wstrb_32(MuxN_io_ins_1_wstrb_32),
    .io_ins_1_wstrb_33(MuxN_io_ins_1_wstrb_33),
    .io_ins_1_wstrb_34(MuxN_io_ins_1_wstrb_34),
    .io_ins_1_wstrb_35(MuxN_io_ins_1_wstrb_35),
    .io_ins_1_wstrb_36(MuxN_io_ins_1_wstrb_36),
    .io_ins_1_wstrb_37(MuxN_io_ins_1_wstrb_37),
    .io_ins_1_wstrb_38(MuxN_io_ins_1_wstrb_38),
    .io_ins_1_wstrb_39(MuxN_io_ins_1_wstrb_39),
    .io_ins_1_wstrb_40(MuxN_io_ins_1_wstrb_40),
    .io_ins_1_wstrb_41(MuxN_io_ins_1_wstrb_41),
    .io_ins_1_wstrb_42(MuxN_io_ins_1_wstrb_42),
    .io_ins_1_wstrb_43(MuxN_io_ins_1_wstrb_43),
    .io_ins_1_wstrb_44(MuxN_io_ins_1_wstrb_44),
    .io_ins_1_wstrb_45(MuxN_io_ins_1_wstrb_45),
    .io_ins_1_wstrb_46(MuxN_io_ins_1_wstrb_46),
    .io_ins_1_wstrb_47(MuxN_io_ins_1_wstrb_47),
    .io_ins_1_wstrb_48(MuxN_io_ins_1_wstrb_48),
    .io_ins_1_wstrb_49(MuxN_io_ins_1_wstrb_49),
    .io_ins_1_wstrb_50(MuxN_io_ins_1_wstrb_50),
    .io_ins_1_wstrb_51(MuxN_io_ins_1_wstrb_51),
    .io_ins_1_wstrb_52(MuxN_io_ins_1_wstrb_52),
    .io_ins_1_wstrb_53(MuxN_io_ins_1_wstrb_53),
    .io_ins_1_wstrb_54(MuxN_io_ins_1_wstrb_54),
    .io_ins_1_wstrb_55(MuxN_io_ins_1_wstrb_55),
    .io_ins_1_wstrb_56(MuxN_io_ins_1_wstrb_56),
    .io_ins_1_wstrb_57(MuxN_io_ins_1_wstrb_57),
    .io_ins_1_wstrb_58(MuxN_io_ins_1_wstrb_58),
    .io_ins_1_wstrb_59(MuxN_io_ins_1_wstrb_59),
    .io_ins_1_wstrb_60(MuxN_io_ins_1_wstrb_60),
    .io_ins_1_wstrb_61(MuxN_io_ins_1_wstrb_61),
    .io_ins_1_wstrb_62(MuxN_io_ins_1_wstrb_62),
    .io_ins_1_wstrb_63(MuxN_io_ins_1_wstrb_63),
    .io_sel(MuxN_io_sel),
    .io_out_wdata_0(MuxN_io_out_wdata_0),
    .io_out_wdata_1(MuxN_io_out_wdata_1),
    .io_out_wdata_2(MuxN_io_out_wdata_2),
    .io_out_wdata_3(MuxN_io_out_wdata_3),
    .io_out_wdata_4(MuxN_io_out_wdata_4),
    .io_out_wdata_5(MuxN_io_out_wdata_5),
    .io_out_wdata_6(MuxN_io_out_wdata_6),
    .io_out_wdata_7(MuxN_io_out_wdata_7),
    .io_out_wdata_8(MuxN_io_out_wdata_8),
    .io_out_wdata_9(MuxN_io_out_wdata_9),
    .io_out_wdata_10(MuxN_io_out_wdata_10),
    .io_out_wdata_11(MuxN_io_out_wdata_11),
    .io_out_wdata_12(MuxN_io_out_wdata_12),
    .io_out_wdata_13(MuxN_io_out_wdata_13),
    .io_out_wdata_14(MuxN_io_out_wdata_14),
    .io_out_wdata_15(MuxN_io_out_wdata_15),
    .io_out_wdata_16(MuxN_io_out_wdata_16),
    .io_out_wdata_17(MuxN_io_out_wdata_17),
    .io_out_wdata_18(MuxN_io_out_wdata_18),
    .io_out_wdata_19(MuxN_io_out_wdata_19),
    .io_out_wdata_20(MuxN_io_out_wdata_20),
    .io_out_wdata_21(MuxN_io_out_wdata_21),
    .io_out_wdata_22(MuxN_io_out_wdata_22),
    .io_out_wdata_23(MuxN_io_out_wdata_23),
    .io_out_wdata_24(MuxN_io_out_wdata_24),
    .io_out_wdata_25(MuxN_io_out_wdata_25),
    .io_out_wdata_26(MuxN_io_out_wdata_26),
    .io_out_wdata_27(MuxN_io_out_wdata_27),
    .io_out_wdata_28(MuxN_io_out_wdata_28),
    .io_out_wdata_29(MuxN_io_out_wdata_29),
    .io_out_wdata_30(MuxN_io_out_wdata_30),
    .io_out_wdata_31(MuxN_io_out_wdata_31),
    .io_out_wdata_32(MuxN_io_out_wdata_32),
    .io_out_wdata_33(MuxN_io_out_wdata_33),
    .io_out_wdata_34(MuxN_io_out_wdata_34),
    .io_out_wdata_35(MuxN_io_out_wdata_35),
    .io_out_wdata_36(MuxN_io_out_wdata_36),
    .io_out_wdata_37(MuxN_io_out_wdata_37),
    .io_out_wdata_38(MuxN_io_out_wdata_38),
    .io_out_wdata_39(MuxN_io_out_wdata_39),
    .io_out_wdata_40(MuxN_io_out_wdata_40),
    .io_out_wdata_41(MuxN_io_out_wdata_41),
    .io_out_wdata_42(MuxN_io_out_wdata_42),
    .io_out_wdata_43(MuxN_io_out_wdata_43),
    .io_out_wdata_44(MuxN_io_out_wdata_44),
    .io_out_wdata_45(MuxN_io_out_wdata_45),
    .io_out_wdata_46(MuxN_io_out_wdata_46),
    .io_out_wdata_47(MuxN_io_out_wdata_47),
    .io_out_wdata_48(MuxN_io_out_wdata_48),
    .io_out_wdata_49(MuxN_io_out_wdata_49),
    .io_out_wdata_50(MuxN_io_out_wdata_50),
    .io_out_wdata_51(MuxN_io_out_wdata_51),
    .io_out_wdata_52(MuxN_io_out_wdata_52),
    .io_out_wdata_53(MuxN_io_out_wdata_53),
    .io_out_wdata_54(MuxN_io_out_wdata_54),
    .io_out_wdata_55(MuxN_io_out_wdata_55),
    .io_out_wdata_56(MuxN_io_out_wdata_56),
    .io_out_wdata_57(MuxN_io_out_wdata_57),
    .io_out_wdata_58(MuxN_io_out_wdata_58),
    .io_out_wdata_59(MuxN_io_out_wdata_59),
    .io_out_wdata_60(MuxN_io_out_wdata_60),
    .io_out_wdata_61(MuxN_io_out_wdata_61),
    .io_out_wdata_62(MuxN_io_out_wdata_62),
    .io_out_wdata_63(MuxN_io_out_wdata_63),
    .io_out_wstrb_0(MuxN_io_out_wstrb_0),
    .io_out_wstrb_1(MuxN_io_out_wstrb_1),
    .io_out_wstrb_2(MuxN_io_out_wstrb_2),
    .io_out_wstrb_3(MuxN_io_out_wstrb_3),
    .io_out_wstrb_4(MuxN_io_out_wstrb_4),
    .io_out_wstrb_5(MuxN_io_out_wstrb_5),
    .io_out_wstrb_6(MuxN_io_out_wstrb_6),
    .io_out_wstrb_7(MuxN_io_out_wstrb_7),
    .io_out_wstrb_8(MuxN_io_out_wstrb_8),
    .io_out_wstrb_9(MuxN_io_out_wstrb_9),
    .io_out_wstrb_10(MuxN_io_out_wstrb_10),
    .io_out_wstrb_11(MuxN_io_out_wstrb_11),
    .io_out_wstrb_12(MuxN_io_out_wstrb_12),
    .io_out_wstrb_13(MuxN_io_out_wstrb_13),
    .io_out_wstrb_14(MuxN_io_out_wstrb_14),
    .io_out_wstrb_15(MuxN_io_out_wstrb_15),
    .io_out_wstrb_16(MuxN_io_out_wstrb_16),
    .io_out_wstrb_17(MuxN_io_out_wstrb_17),
    .io_out_wstrb_18(MuxN_io_out_wstrb_18),
    .io_out_wstrb_19(MuxN_io_out_wstrb_19),
    .io_out_wstrb_20(MuxN_io_out_wstrb_20),
    .io_out_wstrb_21(MuxN_io_out_wstrb_21),
    .io_out_wstrb_22(MuxN_io_out_wstrb_22),
    .io_out_wstrb_23(MuxN_io_out_wstrb_23),
    .io_out_wstrb_24(MuxN_io_out_wstrb_24),
    .io_out_wstrb_25(MuxN_io_out_wstrb_25),
    .io_out_wstrb_26(MuxN_io_out_wstrb_26),
    .io_out_wstrb_27(MuxN_io_out_wstrb_27),
    .io_out_wstrb_28(MuxN_io_out_wstrb_28),
    .io_out_wstrb_29(MuxN_io_out_wstrb_29),
    .io_out_wstrb_30(MuxN_io_out_wstrb_30),
    .io_out_wstrb_31(MuxN_io_out_wstrb_31),
    .io_out_wstrb_32(MuxN_io_out_wstrb_32),
    .io_out_wstrb_33(MuxN_io_out_wstrb_33),
    .io_out_wstrb_34(MuxN_io_out_wstrb_34),
    .io_out_wstrb_35(MuxN_io_out_wstrb_35),
    .io_out_wstrb_36(MuxN_io_out_wstrb_36),
    .io_out_wstrb_37(MuxN_io_out_wstrb_37),
    .io_out_wstrb_38(MuxN_io_out_wstrb_38),
    .io_out_wstrb_39(MuxN_io_out_wstrb_39),
    .io_out_wstrb_40(MuxN_io_out_wstrb_40),
    .io_out_wstrb_41(MuxN_io_out_wstrb_41),
    .io_out_wstrb_42(MuxN_io_out_wstrb_42),
    .io_out_wstrb_43(MuxN_io_out_wstrb_43),
    .io_out_wstrb_44(MuxN_io_out_wstrb_44),
    .io_out_wstrb_45(MuxN_io_out_wstrb_45),
    .io_out_wstrb_46(MuxN_io_out_wstrb_46),
    .io_out_wstrb_47(MuxN_io_out_wstrb_47),
    .io_out_wstrb_48(MuxN_io_out_wstrb_48),
    .io_out_wstrb_49(MuxN_io_out_wstrb_49),
    .io_out_wstrb_50(MuxN_io_out_wstrb_50),
    .io_out_wstrb_51(MuxN_io_out_wstrb_51),
    .io_out_wstrb_52(MuxN_io_out_wstrb_52),
    .io_out_wstrb_53(MuxN_io_out_wstrb_53),
    .io_out_wstrb_54(MuxN_io_out_wstrb_54),
    .io_out_wstrb_55(MuxN_io_out_wstrb_55),
    .io_out_wstrb_56(MuxN_io_out_wstrb_56),
    .io_out_wstrb_57(MuxN_io_out_wstrb_57),
    .io_out_wstrb_58(MuxN_io_out_wstrb_58),
    .io_out_wstrb_59(MuxN_io_out_wstrb_59),
    .io_out_wstrb_60(MuxN_io_out_wstrb_60),
    .io_out_wstrb_61(MuxN_io_out_wstrb_61),
    .io_out_wstrb_62(MuxN_io_out_wstrb_62),
    .io_out_wstrb_63(MuxN_io_out_wstrb_63)
  );
  assign _T_190 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@103120.4]
  assign io_in_ready = io_out_ready | _T_190; // @[MuxN.scala 71:15:@103645.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@103644.4]
  assign io_out_bits_wdata_0 = MuxN_io_out_wdata_0; // @[MuxN.scala 72:15:@103711.4]
  assign io_out_bits_wdata_1 = MuxN_io_out_wdata_1; // @[MuxN.scala 72:15:@103712.4]
  assign io_out_bits_wdata_2 = MuxN_io_out_wdata_2; // @[MuxN.scala 72:15:@103713.4]
  assign io_out_bits_wdata_3 = MuxN_io_out_wdata_3; // @[MuxN.scala 72:15:@103714.4]
  assign io_out_bits_wdata_4 = MuxN_io_out_wdata_4; // @[MuxN.scala 72:15:@103715.4]
  assign io_out_bits_wdata_5 = MuxN_io_out_wdata_5; // @[MuxN.scala 72:15:@103716.4]
  assign io_out_bits_wdata_6 = MuxN_io_out_wdata_6; // @[MuxN.scala 72:15:@103717.4]
  assign io_out_bits_wdata_7 = MuxN_io_out_wdata_7; // @[MuxN.scala 72:15:@103718.4]
  assign io_out_bits_wdata_8 = MuxN_io_out_wdata_8; // @[MuxN.scala 72:15:@103719.4]
  assign io_out_bits_wdata_9 = MuxN_io_out_wdata_9; // @[MuxN.scala 72:15:@103720.4]
  assign io_out_bits_wdata_10 = MuxN_io_out_wdata_10; // @[MuxN.scala 72:15:@103721.4]
  assign io_out_bits_wdata_11 = MuxN_io_out_wdata_11; // @[MuxN.scala 72:15:@103722.4]
  assign io_out_bits_wdata_12 = MuxN_io_out_wdata_12; // @[MuxN.scala 72:15:@103723.4]
  assign io_out_bits_wdata_13 = MuxN_io_out_wdata_13; // @[MuxN.scala 72:15:@103724.4]
  assign io_out_bits_wdata_14 = MuxN_io_out_wdata_14; // @[MuxN.scala 72:15:@103725.4]
  assign io_out_bits_wdata_15 = MuxN_io_out_wdata_15; // @[MuxN.scala 72:15:@103726.4]
  assign io_out_bits_wdata_16 = MuxN_io_out_wdata_16; // @[MuxN.scala 72:15:@103727.4]
  assign io_out_bits_wdata_17 = MuxN_io_out_wdata_17; // @[MuxN.scala 72:15:@103728.4]
  assign io_out_bits_wdata_18 = MuxN_io_out_wdata_18; // @[MuxN.scala 72:15:@103729.4]
  assign io_out_bits_wdata_19 = MuxN_io_out_wdata_19; // @[MuxN.scala 72:15:@103730.4]
  assign io_out_bits_wdata_20 = MuxN_io_out_wdata_20; // @[MuxN.scala 72:15:@103731.4]
  assign io_out_bits_wdata_21 = MuxN_io_out_wdata_21; // @[MuxN.scala 72:15:@103732.4]
  assign io_out_bits_wdata_22 = MuxN_io_out_wdata_22; // @[MuxN.scala 72:15:@103733.4]
  assign io_out_bits_wdata_23 = MuxN_io_out_wdata_23; // @[MuxN.scala 72:15:@103734.4]
  assign io_out_bits_wdata_24 = MuxN_io_out_wdata_24; // @[MuxN.scala 72:15:@103735.4]
  assign io_out_bits_wdata_25 = MuxN_io_out_wdata_25; // @[MuxN.scala 72:15:@103736.4]
  assign io_out_bits_wdata_26 = MuxN_io_out_wdata_26; // @[MuxN.scala 72:15:@103737.4]
  assign io_out_bits_wdata_27 = MuxN_io_out_wdata_27; // @[MuxN.scala 72:15:@103738.4]
  assign io_out_bits_wdata_28 = MuxN_io_out_wdata_28; // @[MuxN.scala 72:15:@103739.4]
  assign io_out_bits_wdata_29 = MuxN_io_out_wdata_29; // @[MuxN.scala 72:15:@103740.4]
  assign io_out_bits_wdata_30 = MuxN_io_out_wdata_30; // @[MuxN.scala 72:15:@103741.4]
  assign io_out_bits_wdata_31 = MuxN_io_out_wdata_31; // @[MuxN.scala 72:15:@103742.4]
  assign io_out_bits_wdata_32 = MuxN_io_out_wdata_32; // @[MuxN.scala 72:15:@103743.4]
  assign io_out_bits_wdata_33 = MuxN_io_out_wdata_33; // @[MuxN.scala 72:15:@103744.4]
  assign io_out_bits_wdata_34 = MuxN_io_out_wdata_34; // @[MuxN.scala 72:15:@103745.4]
  assign io_out_bits_wdata_35 = MuxN_io_out_wdata_35; // @[MuxN.scala 72:15:@103746.4]
  assign io_out_bits_wdata_36 = MuxN_io_out_wdata_36; // @[MuxN.scala 72:15:@103747.4]
  assign io_out_bits_wdata_37 = MuxN_io_out_wdata_37; // @[MuxN.scala 72:15:@103748.4]
  assign io_out_bits_wdata_38 = MuxN_io_out_wdata_38; // @[MuxN.scala 72:15:@103749.4]
  assign io_out_bits_wdata_39 = MuxN_io_out_wdata_39; // @[MuxN.scala 72:15:@103750.4]
  assign io_out_bits_wdata_40 = MuxN_io_out_wdata_40; // @[MuxN.scala 72:15:@103751.4]
  assign io_out_bits_wdata_41 = MuxN_io_out_wdata_41; // @[MuxN.scala 72:15:@103752.4]
  assign io_out_bits_wdata_42 = MuxN_io_out_wdata_42; // @[MuxN.scala 72:15:@103753.4]
  assign io_out_bits_wdata_43 = MuxN_io_out_wdata_43; // @[MuxN.scala 72:15:@103754.4]
  assign io_out_bits_wdata_44 = MuxN_io_out_wdata_44; // @[MuxN.scala 72:15:@103755.4]
  assign io_out_bits_wdata_45 = MuxN_io_out_wdata_45; // @[MuxN.scala 72:15:@103756.4]
  assign io_out_bits_wdata_46 = MuxN_io_out_wdata_46; // @[MuxN.scala 72:15:@103757.4]
  assign io_out_bits_wdata_47 = MuxN_io_out_wdata_47; // @[MuxN.scala 72:15:@103758.4]
  assign io_out_bits_wdata_48 = MuxN_io_out_wdata_48; // @[MuxN.scala 72:15:@103759.4]
  assign io_out_bits_wdata_49 = MuxN_io_out_wdata_49; // @[MuxN.scala 72:15:@103760.4]
  assign io_out_bits_wdata_50 = MuxN_io_out_wdata_50; // @[MuxN.scala 72:15:@103761.4]
  assign io_out_bits_wdata_51 = MuxN_io_out_wdata_51; // @[MuxN.scala 72:15:@103762.4]
  assign io_out_bits_wdata_52 = MuxN_io_out_wdata_52; // @[MuxN.scala 72:15:@103763.4]
  assign io_out_bits_wdata_53 = MuxN_io_out_wdata_53; // @[MuxN.scala 72:15:@103764.4]
  assign io_out_bits_wdata_54 = MuxN_io_out_wdata_54; // @[MuxN.scala 72:15:@103765.4]
  assign io_out_bits_wdata_55 = MuxN_io_out_wdata_55; // @[MuxN.scala 72:15:@103766.4]
  assign io_out_bits_wdata_56 = MuxN_io_out_wdata_56; // @[MuxN.scala 72:15:@103767.4]
  assign io_out_bits_wdata_57 = MuxN_io_out_wdata_57; // @[MuxN.scala 72:15:@103768.4]
  assign io_out_bits_wdata_58 = MuxN_io_out_wdata_58; // @[MuxN.scala 72:15:@103769.4]
  assign io_out_bits_wdata_59 = MuxN_io_out_wdata_59; // @[MuxN.scala 72:15:@103770.4]
  assign io_out_bits_wdata_60 = MuxN_io_out_wdata_60; // @[MuxN.scala 72:15:@103771.4]
  assign io_out_bits_wdata_61 = MuxN_io_out_wdata_61; // @[MuxN.scala 72:15:@103772.4]
  assign io_out_bits_wdata_62 = MuxN_io_out_wdata_62; // @[MuxN.scala 72:15:@103773.4]
  assign io_out_bits_wdata_63 = MuxN_io_out_wdata_63; // @[MuxN.scala 72:15:@103774.4]
  assign io_out_bits_wstrb_0 = MuxN_io_out_wstrb_0; // @[MuxN.scala 72:15:@103647.4]
  assign io_out_bits_wstrb_1 = MuxN_io_out_wstrb_1; // @[MuxN.scala 72:15:@103648.4]
  assign io_out_bits_wstrb_2 = MuxN_io_out_wstrb_2; // @[MuxN.scala 72:15:@103649.4]
  assign io_out_bits_wstrb_3 = MuxN_io_out_wstrb_3; // @[MuxN.scala 72:15:@103650.4]
  assign io_out_bits_wstrb_4 = MuxN_io_out_wstrb_4; // @[MuxN.scala 72:15:@103651.4]
  assign io_out_bits_wstrb_5 = MuxN_io_out_wstrb_5; // @[MuxN.scala 72:15:@103652.4]
  assign io_out_bits_wstrb_6 = MuxN_io_out_wstrb_6; // @[MuxN.scala 72:15:@103653.4]
  assign io_out_bits_wstrb_7 = MuxN_io_out_wstrb_7; // @[MuxN.scala 72:15:@103654.4]
  assign io_out_bits_wstrb_8 = MuxN_io_out_wstrb_8; // @[MuxN.scala 72:15:@103655.4]
  assign io_out_bits_wstrb_9 = MuxN_io_out_wstrb_9; // @[MuxN.scala 72:15:@103656.4]
  assign io_out_bits_wstrb_10 = MuxN_io_out_wstrb_10; // @[MuxN.scala 72:15:@103657.4]
  assign io_out_bits_wstrb_11 = MuxN_io_out_wstrb_11; // @[MuxN.scala 72:15:@103658.4]
  assign io_out_bits_wstrb_12 = MuxN_io_out_wstrb_12; // @[MuxN.scala 72:15:@103659.4]
  assign io_out_bits_wstrb_13 = MuxN_io_out_wstrb_13; // @[MuxN.scala 72:15:@103660.4]
  assign io_out_bits_wstrb_14 = MuxN_io_out_wstrb_14; // @[MuxN.scala 72:15:@103661.4]
  assign io_out_bits_wstrb_15 = MuxN_io_out_wstrb_15; // @[MuxN.scala 72:15:@103662.4]
  assign io_out_bits_wstrb_16 = MuxN_io_out_wstrb_16; // @[MuxN.scala 72:15:@103663.4]
  assign io_out_bits_wstrb_17 = MuxN_io_out_wstrb_17; // @[MuxN.scala 72:15:@103664.4]
  assign io_out_bits_wstrb_18 = MuxN_io_out_wstrb_18; // @[MuxN.scala 72:15:@103665.4]
  assign io_out_bits_wstrb_19 = MuxN_io_out_wstrb_19; // @[MuxN.scala 72:15:@103666.4]
  assign io_out_bits_wstrb_20 = MuxN_io_out_wstrb_20; // @[MuxN.scala 72:15:@103667.4]
  assign io_out_bits_wstrb_21 = MuxN_io_out_wstrb_21; // @[MuxN.scala 72:15:@103668.4]
  assign io_out_bits_wstrb_22 = MuxN_io_out_wstrb_22; // @[MuxN.scala 72:15:@103669.4]
  assign io_out_bits_wstrb_23 = MuxN_io_out_wstrb_23; // @[MuxN.scala 72:15:@103670.4]
  assign io_out_bits_wstrb_24 = MuxN_io_out_wstrb_24; // @[MuxN.scala 72:15:@103671.4]
  assign io_out_bits_wstrb_25 = MuxN_io_out_wstrb_25; // @[MuxN.scala 72:15:@103672.4]
  assign io_out_bits_wstrb_26 = MuxN_io_out_wstrb_26; // @[MuxN.scala 72:15:@103673.4]
  assign io_out_bits_wstrb_27 = MuxN_io_out_wstrb_27; // @[MuxN.scala 72:15:@103674.4]
  assign io_out_bits_wstrb_28 = MuxN_io_out_wstrb_28; // @[MuxN.scala 72:15:@103675.4]
  assign io_out_bits_wstrb_29 = MuxN_io_out_wstrb_29; // @[MuxN.scala 72:15:@103676.4]
  assign io_out_bits_wstrb_30 = MuxN_io_out_wstrb_30; // @[MuxN.scala 72:15:@103677.4]
  assign io_out_bits_wstrb_31 = MuxN_io_out_wstrb_31; // @[MuxN.scala 72:15:@103678.4]
  assign io_out_bits_wstrb_32 = MuxN_io_out_wstrb_32; // @[MuxN.scala 72:15:@103679.4]
  assign io_out_bits_wstrb_33 = MuxN_io_out_wstrb_33; // @[MuxN.scala 72:15:@103680.4]
  assign io_out_bits_wstrb_34 = MuxN_io_out_wstrb_34; // @[MuxN.scala 72:15:@103681.4]
  assign io_out_bits_wstrb_35 = MuxN_io_out_wstrb_35; // @[MuxN.scala 72:15:@103682.4]
  assign io_out_bits_wstrb_36 = MuxN_io_out_wstrb_36; // @[MuxN.scala 72:15:@103683.4]
  assign io_out_bits_wstrb_37 = MuxN_io_out_wstrb_37; // @[MuxN.scala 72:15:@103684.4]
  assign io_out_bits_wstrb_38 = MuxN_io_out_wstrb_38; // @[MuxN.scala 72:15:@103685.4]
  assign io_out_bits_wstrb_39 = MuxN_io_out_wstrb_39; // @[MuxN.scala 72:15:@103686.4]
  assign io_out_bits_wstrb_40 = MuxN_io_out_wstrb_40; // @[MuxN.scala 72:15:@103687.4]
  assign io_out_bits_wstrb_41 = MuxN_io_out_wstrb_41; // @[MuxN.scala 72:15:@103688.4]
  assign io_out_bits_wstrb_42 = MuxN_io_out_wstrb_42; // @[MuxN.scala 72:15:@103689.4]
  assign io_out_bits_wstrb_43 = MuxN_io_out_wstrb_43; // @[MuxN.scala 72:15:@103690.4]
  assign io_out_bits_wstrb_44 = MuxN_io_out_wstrb_44; // @[MuxN.scala 72:15:@103691.4]
  assign io_out_bits_wstrb_45 = MuxN_io_out_wstrb_45; // @[MuxN.scala 72:15:@103692.4]
  assign io_out_bits_wstrb_46 = MuxN_io_out_wstrb_46; // @[MuxN.scala 72:15:@103693.4]
  assign io_out_bits_wstrb_47 = MuxN_io_out_wstrb_47; // @[MuxN.scala 72:15:@103694.4]
  assign io_out_bits_wstrb_48 = MuxN_io_out_wstrb_48; // @[MuxN.scala 72:15:@103695.4]
  assign io_out_bits_wstrb_49 = MuxN_io_out_wstrb_49; // @[MuxN.scala 72:15:@103696.4]
  assign io_out_bits_wstrb_50 = MuxN_io_out_wstrb_50; // @[MuxN.scala 72:15:@103697.4]
  assign io_out_bits_wstrb_51 = MuxN_io_out_wstrb_51; // @[MuxN.scala 72:15:@103698.4]
  assign io_out_bits_wstrb_52 = MuxN_io_out_wstrb_52; // @[MuxN.scala 72:15:@103699.4]
  assign io_out_bits_wstrb_53 = MuxN_io_out_wstrb_53; // @[MuxN.scala 72:15:@103700.4]
  assign io_out_bits_wstrb_54 = MuxN_io_out_wstrb_54; // @[MuxN.scala 72:15:@103701.4]
  assign io_out_bits_wstrb_55 = MuxN_io_out_wstrb_55; // @[MuxN.scala 72:15:@103702.4]
  assign io_out_bits_wstrb_56 = MuxN_io_out_wstrb_56; // @[MuxN.scala 72:15:@103703.4]
  assign io_out_bits_wstrb_57 = MuxN_io_out_wstrb_57; // @[MuxN.scala 72:15:@103704.4]
  assign io_out_bits_wstrb_58 = MuxN_io_out_wstrb_58; // @[MuxN.scala 72:15:@103705.4]
  assign io_out_bits_wstrb_59 = MuxN_io_out_wstrb_59; // @[MuxN.scala 72:15:@103706.4]
  assign io_out_bits_wstrb_60 = MuxN_io_out_wstrb_60; // @[MuxN.scala 72:15:@103707.4]
  assign io_out_bits_wstrb_61 = MuxN_io_out_wstrb_61; // @[MuxN.scala 72:15:@103708.4]
  assign io_out_bits_wstrb_62 = MuxN_io_out_wstrb_62; // @[MuxN.scala 72:15:@103709.4]
  assign io_out_bits_wstrb_63 = MuxN_io_out_wstrb_63; // @[MuxN.scala 72:15:@103710.4]
  assign MuxN_io_ins_1_wdata_0 = io_in_bits_1_wdata_0; // @[MuxN.scala 41:18:@103578.4]
  assign MuxN_io_ins_1_wdata_1 = io_in_bits_1_wdata_1; // @[MuxN.scala 41:18:@103579.4]
  assign MuxN_io_ins_1_wdata_2 = io_in_bits_1_wdata_2; // @[MuxN.scala 41:18:@103580.4]
  assign MuxN_io_ins_1_wdata_3 = io_in_bits_1_wdata_3; // @[MuxN.scala 41:18:@103581.4]
  assign MuxN_io_ins_1_wdata_4 = io_in_bits_1_wdata_4; // @[MuxN.scala 41:18:@103582.4]
  assign MuxN_io_ins_1_wdata_5 = io_in_bits_1_wdata_5; // @[MuxN.scala 41:18:@103583.4]
  assign MuxN_io_ins_1_wdata_6 = io_in_bits_1_wdata_6; // @[MuxN.scala 41:18:@103584.4]
  assign MuxN_io_ins_1_wdata_7 = io_in_bits_1_wdata_7; // @[MuxN.scala 41:18:@103585.4]
  assign MuxN_io_ins_1_wdata_8 = io_in_bits_1_wdata_8; // @[MuxN.scala 41:18:@103586.4]
  assign MuxN_io_ins_1_wdata_9 = io_in_bits_1_wdata_9; // @[MuxN.scala 41:18:@103587.4]
  assign MuxN_io_ins_1_wdata_10 = io_in_bits_1_wdata_10; // @[MuxN.scala 41:18:@103588.4]
  assign MuxN_io_ins_1_wdata_11 = io_in_bits_1_wdata_11; // @[MuxN.scala 41:18:@103589.4]
  assign MuxN_io_ins_1_wdata_12 = io_in_bits_1_wdata_12; // @[MuxN.scala 41:18:@103590.4]
  assign MuxN_io_ins_1_wdata_13 = io_in_bits_1_wdata_13; // @[MuxN.scala 41:18:@103591.4]
  assign MuxN_io_ins_1_wdata_14 = io_in_bits_1_wdata_14; // @[MuxN.scala 41:18:@103592.4]
  assign MuxN_io_ins_1_wdata_15 = io_in_bits_1_wdata_15; // @[MuxN.scala 41:18:@103593.4]
  assign MuxN_io_ins_1_wdata_16 = io_in_bits_1_wdata_16; // @[MuxN.scala 41:18:@103594.4]
  assign MuxN_io_ins_1_wdata_17 = io_in_bits_1_wdata_17; // @[MuxN.scala 41:18:@103595.4]
  assign MuxN_io_ins_1_wdata_18 = io_in_bits_1_wdata_18; // @[MuxN.scala 41:18:@103596.4]
  assign MuxN_io_ins_1_wdata_19 = io_in_bits_1_wdata_19; // @[MuxN.scala 41:18:@103597.4]
  assign MuxN_io_ins_1_wdata_20 = io_in_bits_1_wdata_20; // @[MuxN.scala 41:18:@103598.4]
  assign MuxN_io_ins_1_wdata_21 = io_in_bits_1_wdata_21; // @[MuxN.scala 41:18:@103599.4]
  assign MuxN_io_ins_1_wdata_22 = io_in_bits_1_wdata_22; // @[MuxN.scala 41:18:@103600.4]
  assign MuxN_io_ins_1_wdata_23 = io_in_bits_1_wdata_23; // @[MuxN.scala 41:18:@103601.4]
  assign MuxN_io_ins_1_wdata_24 = io_in_bits_1_wdata_24; // @[MuxN.scala 41:18:@103602.4]
  assign MuxN_io_ins_1_wdata_25 = io_in_bits_1_wdata_25; // @[MuxN.scala 41:18:@103603.4]
  assign MuxN_io_ins_1_wdata_26 = io_in_bits_1_wdata_26; // @[MuxN.scala 41:18:@103604.4]
  assign MuxN_io_ins_1_wdata_27 = io_in_bits_1_wdata_27; // @[MuxN.scala 41:18:@103605.4]
  assign MuxN_io_ins_1_wdata_28 = io_in_bits_1_wdata_28; // @[MuxN.scala 41:18:@103606.4]
  assign MuxN_io_ins_1_wdata_29 = io_in_bits_1_wdata_29; // @[MuxN.scala 41:18:@103607.4]
  assign MuxN_io_ins_1_wdata_30 = io_in_bits_1_wdata_30; // @[MuxN.scala 41:18:@103608.4]
  assign MuxN_io_ins_1_wdata_31 = io_in_bits_1_wdata_31; // @[MuxN.scala 41:18:@103609.4]
  assign MuxN_io_ins_1_wdata_32 = io_in_bits_1_wdata_32; // @[MuxN.scala 41:18:@103610.4]
  assign MuxN_io_ins_1_wdata_33 = io_in_bits_1_wdata_33; // @[MuxN.scala 41:18:@103611.4]
  assign MuxN_io_ins_1_wdata_34 = io_in_bits_1_wdata_34; // @[MuxN.scala 41:18:@103612.4]
  assign MuxN_io_ins_1_wdata_35 = io_in_bits_1_wdata_35; // @[MuxN.scala 41:18:@103613.4]
  assign MuxN_io_ins_1_wdata_36 = io_in_bits_1_wdata_36; // @[MuxN.scala 41:18:@103614.4]
  assign MuxN_io_ins_1_wdata_37 = io_in_bits_1_wdata_37; // @[MuxN.scala 41:18:@103615.4]
  assign MuxN_io_ins_1_wdata_38 = io_in_bits_1_wdata_38; // @[MuxN.scala 41:18:@103616.4]
  assign MuxN_io_ins_1_wdata_39 = io_in_bits_1_wdata_39; // @[MuxN.scala 41:18:@103617.4]
  assign MuxN_io_ins_1_wdata_40 = io_in_bits_1_wdata_40; // @[MuxN.scala 41:18:@103618.4]
  assign MuxN_io_ins_1_wdata_41 = io_in_bits_1_wdata_41; // @[MuxN.scala 41:18:@103619.4]
  assign MuxN_io_ins_1_wdata_42 = io_in_bits_1_wdata_42; // @[MuxN.scala 41:18:@103620.4]
  assign MuxN_io_ins_1_wdata_43 = io_in_bits_1_wdata_43; // @[MuxN.scala 41:18:@103621.4]
  assign MuxN_io_ins_1_wdata_44 = io_in_bits_1_wdata_44; // @[MuxN.scala 41:18:@103622.4]
  assign MuxN_io_ins_1_wdata_45 = io_in_bits_1_wdata_45; // @[MuxN.scala 41:18:@103623.4]
  assign MuxN_io_ins_1_wdata_46 = io_in_bits_1_wdata_46; // @[MuxN.scala 41:18:@103624.4]
  assign MuxN_io_ins_1_wdata_47 = io_in_bits_1_wdata_47; // @[MuxN.scala 41:18:@103625.4]
  assign MuxN_io_ins_1_wdata_48 = io_in_bits_1_wdata_48; // @[MuxN.scala 41:18:@103626.4]
  assign MuxN_io_ins_1_wdata_49 = io_in_bits_1_wdata_49; // @[MuxN.scala 41:18:@103627.4]
  assign MuxN_io_ins_1_wdata_50 = io_in_bits_1_wdata_50; // @[MuxN.scala 41:18:@103628.4]
  assign MuxN_io_ins_1_wdata_51 = io_in_bits_1_wdata_51; // @[MuxN.scala 41:18:@103629.4]
  assign MuxN_io_ins_1_wdata_52 = io_in_bits_1_wdata_52; // @[MuxN.scala 41:18:@103630.4]
  assign MuxN_io_ins_1_wdata_53 = io_in_bits_1_wdata_53; // @[MuxN.scala 41:18:@103631.4]
  assign MuxN_io_ins_1_wdata_54 = io_in_bits_1_wdata_54; // @[MuxN.scala 41:18:@103632.4]
  assign MuxN_io_ins_1_wdata_55 = io_in_bits_1_wdata_55; // @[MuxN.scala 41:18:@103633.4]
  assign MuxN_io_ins_1_wdata_56 = io_in_bits_1_wdata_56; // @[MuxN.scala 41:18:@103634.4]
  assign MuxN_io_ins_1_wdata_57 = io_in_bits_1_wdata_57; // @[MuxN.scala 41:18:@103635.4]
  assign MuxN_io_ins_1_wdata_58 = io_in_bits_1_wdata_58; // @[MuxN.scala 41:18:@103636.4]
  assign MuxN_io_ins_1_wdata_59 = io_in_bits_1_wdata_59; // @[MuxN.scala 41:18:@103637.4]
  assign MuxN_io_ins_1_wdata_60 = io_in_bits_1_wdata_60; // @[MuxN.scala 41:18:@103638.4]
  assign MuxN_io_ins_1_wdata_61 = io_in_bits_1_wdata_61; // @[MuxN.scala 41:18:@103639.4]
  assign MuxN_io_ins_1_wdata_62 = io_in_bits_1_wdata_62; // @[MuxN.scala 41:18:@103640.4]
  assign MuxN_io_ins_1_wdata_63 = io_in_bits_1_wdata_63; // @[MuxN.scala 41:18:@103641.4]
  assign MuxN_io_ins_1_wstrb_0 = io_in_bits_1_wstrb_0; // @[MuxN.scala 41:18:@103514.4]
  assign MuxN_io_ins_1_wstrb_1 = io_in_bits_1_wstrb_1; // @[MuxN.scala 41:18:@103515.4]
  assign MuxN_io_ins_1_wstrb_2 = io_in_bits_1_wstrb_2; // @[MuxN.scala 41:18:@103516.4]
  assign MuxN_io_ins_1_wstrb_3 = io_in_bits_1_wstrb_3; // @[MuxN.scala 41:18:@103517.4]
  assign MuxN_io_ins_1_wstrb_4 = io_in_bits_1_wstrb_4; // @[MuxN.scala 41:18:@103518.4]
  assign MuxN_io_ins_1_wstrb_5 = io_in_bits_1_wstrb_5; // @[MuxN.scala 41:18:@103519.4]
  assign MuxN_io_ins_1_wstrb_6 = io_in_bits_1_wstrb_6; // @[MuxN.scala 41:18:@103520.4]
  assign MuxN_io_ins_1_wstrb_7 = io_in_bits_1_wstrb_7; // @[MuxN.scala 41:18:@103521.4]
  assign MuxN_io_ins_1_wstrb_8 = io_in_bits_1_wstrb_8; // @[MuxN.scala 41:18:@103522.4]
  assign MuxN_io_ins_1_wstrb_9 = io_in_bits_1_wstrb_9; // @[MuxN.scala 41:18:@103523.4]
  assign MuxN_io_ins_1_wstrb_10 = io_in_bits_1_wstrb_10; // @[MuxN.scala 41:18:@103524.4]
  assign MuxN_io_ins_1_wstrb_11 = io_in_bits_1_wstrb_11; // @[MuxN.scala 41:18:@103525.4]
  assign MuxN_io_ins_1_wstrb_12 = io_in_bits_1_wstrb_12; // @[MuxN.scala 41:18:@103526.4]
  assign MuxN_io_ins_1_wstrb_13 = io_in_bits_1_wstrb_13; // @[MuxN.scala 41:18:@103527.4]
  assign MuxN_io_ins_1_wstrb_14 = io_in_bits_1_wstrb_14; // @[MuxN.scala 41:18:@103528.4]
  assign MuxN_io_ins_1_wstrb_15 = io_in_bits_1_wstrb_15; // @[MuxN.scala 41:18:@103529.4]
  assign MuxN_io_ins_1_wstrb_16 = io_in_bits_1_wstrb_16; // @[MuxN.scala 41:18:@103530.4]
  assign MuxN_io_ins_1_wstrb_17 = io_in_bits_1_wstrb_17; // @[MuxN.scala 41:18:@103531.4]
  assign MuxN_io_ins_1_wstrb_18 = io_in_bits_1_wstrb_18; // @[MuxN.scala 41:18:@103532.4]
  assign MuxN_io_ins_1_wstrb_19 = io_in_bits_1_wstrb_19; // @[MuxN.scala 41:18:@103533.4]
  assign MuxN_io_ins_1_wstrb_20 = io_in_bits_1_wstrb_20; // @[MuxN.scala 41:18:@103534.4]
  assign MuxN_io_ins_1_wstrb_21 = io_in_bits_1_wstrb_21; // @[MuxN.scala 41:18:@103535.4]
  assign MuxN_io_ins_1_wstrb_22 = io_in_bits_1_wstrb_22; // @[MuxN.scala 41:18:@103536.4]
  assign MuxN_io_ins_1_wstrb_23 = io_in_bits_1_wstrb_23; // @[MuxN.scala 41:18:@103537.4]
  assign MuxN_io_ins_1_wstrb_24 = io_in_bits_1_wstrb_24; // @[MuxN.scala 41:18:@103538.4]
  assign MuxN_io_ins_1_wstrb_25 = io_in_bits_1_wstrb_25; // @[MuxN.scala 41:18:@103539.4]
  assign MuxN_io_ins_1_wstrb_26 = io_in_bits_1_wstrb_26; // @[MuxN.scala 41:18:@103540.4]
  assign MuxN_io_ins_1_wstrb_27 = io_in_bits_1_wstrb_27; // @[MuxN.scala 41:18:@103541.4]
  assign MuxN_io_ins_1_wstrb_28 = io_in_bits_1_wstrb_28; // @[MuxN.scala 41:18:@103542.4]
  assign MuxN_io_ins_1_wstrb_29 = io_in_bits_1_wstrb_29; // @[MuxN.scala 41:18:@103543.4]
  assign MuxN_io_ins_1_wstrb_30 = io_in_bits_1_wstrb_30; // @[MuxN.scala 41:18:@103544.4]
  assign MuxN_io_ins_1_wstrb_31 = io_in_bits_1_wstrb_31; // @[MuxN.scala 41:18:@103545.4]
  assign MuxN_io_ins_1_wstrb_32 = io_in_bits_1_wstrb_32; // @[MuxN.scala 41:18:@103546.4]
  assign MuxN_io_ins_1_wstrb_33 = io_in_bits_1_wstrb_33; // @[MuxN.scala 41:18:@103547.4]
  assign MuxN_io_ins_1_wstrb_34 = io_in_bits_1_wstrb_34; // @[MuxN.scala 41:18:@103548.4]
  assign MuxN_io_ins_1_wstrb_35 = io_in_bits_1_wstrb_35; // @[MuxN.scala 41:18:@103549.4]
  assign MuxN_io_ins_1_wstrb_36 = io_in_bits_1_wstrb_36; // @[MuxN.scala 41:18:@103550.4]
  assign MuxN_io_ins_1_wstrb_37 = io_in_bits_1_wstrb_37; // @[MuxN.scala 41:18:@103551.4]
  assign MuxN_io_ins_1_wstrb_38 = io_in_bits_1_wstrb_38; // @[MuxN.scala 41:18:@103552.4]
  assign MuxN_io_ins_1_wstrb_39 = io_in_bits_1_wstrb_39; // @[MuxN.scala 41:18:@103553.4]
  assign MuxN_io_ins_1_wstrb_40 = io_in_bits_1_wstrb_40; // @[MuxN.scala 41:18:@103554.4]
  assign MuxN_io_ins_1_wstrb_41 = io_in_bits_1_wstrb_41; // @[MuxN.scala 41:18:@103555.4]
  assign MuxN_io_ins_1_wstrb_42 = io_in_bits_1_wstrb_42; // @[MuxN.scala 41:18:@103556.4]
  assign MuxN_io_ins_1_wstrb_43 = io_in_bits_1_wstrb_43; // @[MuxN.scala 41:18:@103557.4]
  assign MuxN_io_ins_1_wstrb_44 = io_in_bits_1_wstrb_44; // @[MuxN.scala 41:18:@103558.4]
  assign MuxN_io_ins_1_wstrb_45 = io_in_bits_1_wstrb_45; // @[MuxN.scala 41:18:@103559.4]
  assign MuxN_io_ins_1_wstrb_46 = io_in_bits_1_wstrb_46; // @[MuxN.scala 41:18:@103560.4]
  assign MuxN_io_ins_1_wstrb_47 = io_in_bits_1_wstrb_47; // @[MuxN.scala 41:18:@103561.4]
  assign MuxN_io_ins_1_wstrb_48 = io_in_bits_1_wstrb_48; // @[MuxN.scala 41:18:@103562.4]
  assign MuxN_io_ins_1_wstrb_49 = io_in_bits_1_wstrb_49; // @[MuxN.scala 41:18:@103563.4]
  assign MuxN_io_ins_1_wstrb_50 = io_in_bits_1_wstrb_50; // @[MuxN.scala 41:18:@103564.4]
  assign MuxN_io_ins_1_wstrb_51 = io_in_bits_1_wstrb_51; // @[MuxN.scala 41:18:@103565.4]
  assign MuxN_io_ins_1_wstrb_52 = io_in_bits_1_wstrb_52; // @[MuxN.scala 41:18:@103566.4]
  assign MuxN_io_ins_1_wstrb_53 = io_in_bits_1_wstrb_53; // @[MuxN.scala 41:18:@103567.4]
  assign MuxN_io_ins_1_wstrb_54 = io_in_bits_1_wstrb_54; // @[MuxN.scala 41:18:@103568.4]
  assign MuxN_io_ins_1_wstrb_55 = io_in_bits_1_wstrb_55; // @[MuxN.scala 41:18:@103569.4]
  assign MuxN_io_ins_1_wstrb_56 = io_in_bits_1_wstrb_56; // @[MuxN.scala 41:18:@103570.4]
  assign MuxN_io_ins_1_wstrb_57 = io_in_bits_1_wstrb_57; // @[MuxN.scala 41:18:@103571.4]
  assign MuxN_io_ins_1_wstrb_58 = io_in_bits_1_wstrb_58; // @[MuxN.scala 41:18:@103572.4]
  assign MuxN_io_ins_1_wstrb_59 = io_in_bits_1_wstrb_59; // @[MuxN.scala 41:18:@103573.4]
  assign MuxN_io_ins_1_wstrb_60 = io_in_bits_1_wstrb_60; // @[MuxN.scala 41:18:@103574.4]
  assign MuxN_io_ins_1_wstrb_61 = io_in_bits_1_wstrb_61; // @[MuxN.scala 41:18:@103575.4]
  assign MuxN_io_ins_1_wstrb_62 = io_in_bits_1_wstrb_62; // @[MuxN.scala 41:18:@103576.4]
  assign MuxN_io_ins_1_wstrb_63 = io_in_bits_1_wstrb_63; // @[MuxN.scala 41:18:@103577.4]
  assign MuxN_io_sel = io_sel; // @[MuxN.scala 44:18:@103643.4]
endmodule
module ElementCounter( // @[:@103776.2]
  input         clock, // @[:@103777.4]
  input         reset, // @[:@103778.4]
  input         io_reset, // @[:@103779.4]
  input         io_enable, // @[:@103779.4]
  output [31:0] io_out // @[:@103779.4]
);
  reg [31:0] count; // @[Counter.scala 37:22:@103781.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_14; // @[Counter.scala 39:24:@103782.4]
  wire [31:0] newCount; // @[Counter.scala 39:24:@103783.4]
  wire [31:0] _GEN_0; // @[Counter.scala 43:26:@103788.6]
  wire [31:0] _GEN_1; // @[Counter.scala 41:18:@103784.4]
  assign _T_14 = count + 32'h1; // @[Counter.scala 39:24:@103782.4]
  assign newCount = count + 32'h1; // @[Counter.scala 39:24:@103783.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 43:26:@103788.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 41:18:@103784.4]
  assign io_out = count; // @[Counter.scala 47:10:@103791.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module StreamArbiter( // @[:@103793.2]
  input         clock, // @[:@103794.4]
  input         reset, // @[:@103795.4]
  output        io_app_0_cmd_ready, // @[:@103796.4]
  input         io_app_0_cmd_valid, // @[:@103796.4]
  input  [63:0] io_app_0_cmd_bits_addr, // @[:@103796.4]
  input  [31:0] io_app_0_cmd_bits_size, // @[:@103796.4]
  input         io_app_0_rresp_ready, // @[:@103796.4]
  output        io_app_0_rresp_valid, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_0, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_1, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_2, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_3, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_4, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_5, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_6, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_7, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_8, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_9, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_10, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_11, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_12, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_13, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_14, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_15, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_16, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_17, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_18, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_19, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_20, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_21, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_22, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_23, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_24, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_25, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_26, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_27, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_28, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_29, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_30, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_31, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_32, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_33, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_34, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_35, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_36, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_37, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_38, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_39, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_40, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_41, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_42, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_43, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_44, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_45, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_46, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_47, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_48, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_49, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_50, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_51, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_52, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_53, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_54, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_55, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_56, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_57, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_58, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_59, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_60, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_61, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_62, // @[:@103796.4]
  output [7:0]  io_app_0_rresp_bits_rdata_63, // @[:@103796.4]
  output        io_app_1_cmd_ready, // @[:@103796.4]
  input         io_app_1_cmd_valid, // @[:@103796.4]
  input  [63:0] io_app_1_cmd_bits_addr, // @[:@103796.4]
  input  [31:0] io_app_1_cmd_bits_size, // @[:@103796.4]
  output        io_app_1_wdata_ready, // @[:@103796.4]
  input         io_app_1_wdata_valid, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_0, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_1, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_2, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_3, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_4, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_5, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_6, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_7, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_8, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_9, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_10, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_11, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_12, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_13, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_14, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_15, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_16, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_17, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_18, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_19, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_20, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_21, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_22, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_23, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_24, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_25, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_26, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_27, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_28, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_29, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_30, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_31, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_32, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_33, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_34, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_35, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_36, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_37, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_38, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_39, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_40, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_41, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_42, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_43, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_44, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_45, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_46, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_47, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_48, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_49, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_50, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_51, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_52, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_53, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_54, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_55, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_56, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_57, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_58, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_59, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_60, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_61, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_62, // @[:@103796.4]
  input  [7:0]  io_app_1_wdata_bits_wdata_63, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_0, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_1, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_2, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_3, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_4, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_5, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_6, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_7, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_8, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_9, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_10, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_11, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_12, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_13, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_14, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_15, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_16, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_17, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_18, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_19, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_20, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_21, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_22, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_23, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_24, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_25, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_26, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_27, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_28, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_29, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_30, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_31, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_32, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_33, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_34, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_35, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_36, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_37, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_38, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_39, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_40, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_41, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_42, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_43, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_44, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_45, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_46, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_47, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_48, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_49, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_50, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_51, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_52, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_53, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_54, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_55, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_56, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_57, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_58, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_59, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_60, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_61, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_62, // @[:@103796.4]
  input         io_app_1_wdata_bits_wstrb_63, // @[:@103796.4]
  input         io_app_1_wresp_ready, // @[:@103796.4]
  output        io_app_1_wresp_valid, // @[:@103796.4]
  input         io_dram_cmd_ready, // @[:@103796.4]
  output        io_dram_cmd_valid, // @[:@103796.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@103796.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@103796.4]
  output        io_dram_cmd_bits_isWr, // @[:@103796.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@103796.4]
  input         io_dram_wdata_ready, // @[:@103796.4]
  output        io_dram_wdata_valid, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_0, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_1, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_2, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_3, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_4, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_5, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_6, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_7, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_8, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_9, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_10, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_11, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_12, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_13, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_14, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_15, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_16, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_17, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_18, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_19, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_20, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_21, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_22, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_23, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_24, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_25, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_26, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_27, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_28, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_29, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_30, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_31, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_32, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_33, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_34, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_35, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_36, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_37, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_38, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_39, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_40, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_41, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_42, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_43, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_44, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_45, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_46, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_47, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_48, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_49, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_50, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_51, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_52, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_53, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_54, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_55, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_56, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_57, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_58, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_59, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_60, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_61, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_62, // @[:@103796.4]
  output [7:0]  io_dram_wdata_bits_wdata_63, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@103796.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@103796.4]
  output        io_dram_rresp_ready, // @[:@103796.4]
  input         io_dram_rresp_valid, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_0, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_1, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_2, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_3, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_4, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_5, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_6, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_7, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_8, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_9, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_10, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_11, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_12, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_13, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_14, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_15, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_16, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_17, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_18, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_19, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_20, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_21, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_22, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_23, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_24, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_25, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_26, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_27, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_28, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_29, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_30, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_31, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_32, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_33, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_34, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_35, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_36, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_37, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_38, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_39, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_40, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_41, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_42, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_43, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_44, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_45, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_46, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_47, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_48, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_49, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_50, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_51, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_52, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_53, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_54, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_55, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_56, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_57, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_58, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_59, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_60, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_61, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_62, // @[:@103796.4]
  input  [7:0]  io_dram_rresp_bits_rdata_63, // @[:@103796.4]
  input  [31:0] io_dram_rresp_bits_tag, // @[:@103796.4]
  output        io_dram_wresp_ready, // @[:@103796.4]
  input         io_dram_wresp_valid, // @[:@103796.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@103796.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@104427.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@104427.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@104427.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@104427.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@104427.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@104434.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@104434.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@104434.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@104434.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@104434.4]
  wire  cmdMux_io_in_ready; // @[StreamArbiter.scala 25:22:@104444.4]
  wire  cmdMux_io_in_valid; // @[StreamArbiter.scala 25:22:@104444.4]
  wire [63:0] cmdMux_io_in_bits_0_addr; // @[StreamArbiter.scala 25:22:@104444.4]
  wire [31:0] cmdMux_io_in_bits_0_size; // @[StreamArbiter.scala 25:22:@104444.4]
  wire [63:0] cmdMux_io_in_bits_1_addr; // @[StreamArbiter.scala 25:22:@104444.4]
  wire [31:0] cmdMux_io_in_bits_1_size; // @[StreamArbiter.scala 25:22:@104444.4]
  wire  cmdMux_io_sel; // @[StreamArbiter.scala 25:22:@104444.4]
  wire  cmdMux_io_out_ready; // @[StreamArbiter.scala 25:22:@104444.4]
  wire  cmdMux_io_out_valid; // @[StreamArbiter.scala 25:22:@104444.4]
  wire [63:0] cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 25:22:@104444.4]
  wire [31:0] cmdMux_io_out_bits_size; // @[StreamArbiter.scala 25:22:@104444.4]
  wire  cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 25:22:@104444.4]
  wire [31:0] cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 25:22:@104444.4]
  wire  wdataMux_io_in_ready; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_valid; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_0; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_1; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_2; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_3; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_4; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_5; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_6; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_7; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_8; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_9; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_10; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_11; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_12; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_13; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_14; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_15; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_16; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_17; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_18; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_19; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_20; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_21; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_22; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_23; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_24; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_25; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_26; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_27; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_28; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_29; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_30; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_31; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_32; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_33; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_34; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_35; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_36; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_37; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_38; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_39; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_40; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_41; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_42; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_43; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_44; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_45; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_46; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_47; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_48; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_49; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_50; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_51; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_52; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_53; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_54; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_55; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_56; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_57; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_58; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_59; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_60; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_61; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_62; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_in_bits_1_wdata_63; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_0; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_1; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_2; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_3; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_4; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_5; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_6; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_7; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_8; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_9; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_10; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_11; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_12; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_13; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_14; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_15; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_16; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_17; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_18; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_19; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_20; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_21; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_22; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_23; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_24; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_25; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_26; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_27; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_28; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_29; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_30; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_31; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_32; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_33; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_34; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_35; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_36; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_37; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_38; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_39; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_40; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_41; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_42; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_43; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_44; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_45; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_46; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_47; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_48; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_49; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_50; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_51; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_52; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_53; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_54; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_55; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_56; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_57; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_58; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_59; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_60; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_61; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_62; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_in_bits_1_wstrb_63; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_sel; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_ready; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_valid; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_16; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_17; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_18; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_19; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_20; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_21; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_22; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_23; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_24; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_25; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_26; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_27; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_28; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_29; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_30; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_31; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_32; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_33; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_34; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_35; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_36; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_37; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_38; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_39; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_40; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_41; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_42; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_43; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_44; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_45; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_46; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_47; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_48; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_49; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_50; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_51; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_52; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_53; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_54; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_55; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_56; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_57; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_58; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_59; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_60; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_61; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_62; // @[StreamArbiter.scala 35:24:@104486.4]
  wire [7:0] wdataMux_io_out_bits_wdata_63; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 35:24:@104486.4]
  wire  elementCtr_clock; // @[StreamArbiter.scala 36:26:@104489.4]
  wire  elementCtr_reset; // @[StreamArbiter.scala 36:26:@104489.4]
  wire  elementCtr_io_reset; // @[StreamArbiter.scala 36:26:@104489.4]
  wire  elementCtr_io_enable; // @[StreamArbiter.scala 36:26:@104489.4]
  wire [31:0] elementCtr_io_out; // @[StreamArbiter.scala 36:26:@104489.4]
  wire  priorityActive; // @[Mux.scala 31:69:@104422.4]
  wire  _T_408; // @[package.scala 96:25:@104432.4 package.scala 96:25:@104433.4]
  wire  _GEN_1; // @[StreamArbiter.scala 21:16:@104441.4]
  wire  _T_412; // @[package.scala 96:25:@104439.4 package.scala 96:25:@104440.4]
  wire  cmdIdx; // @[StreamArbiter.scala 21:16:@104441.4]
  wire [1:0] cmdInDecoder; // @[OneHot.scala 45:35:@104443.4]
  wire  _T_438; // @[StreamArbiter.scala 37:49:@104492.4]
  wire [31:0] _T_443; // @[:@104496.4 :@104497.4]
  wire [7:0] _T_444; // @[FringeBundles.scala 114:28:@104498.4]
  wire [255:0] cmdOutDecoder; // @[OneHot.scala 45:35:@104504.4]
  wire  _T_457; // @[:@104508.4]
  wire  _GEN_3; // @[StreamArbiter.scala 42:78:@104509.4]
  wire  _T_458; // @[StreamArbiter.scala 42:78:@104509.4]
  wire  _T_459; // @[StreamArbiter.scala 42:121:@104510.4]
  wire [7:0] _T_466; // @[FringeBundles.scala 132:28:@104913.4]
  wire [7:0] _T_474; // @[FringeBundles.scala 140:28:@104922.4]
  wire [255:0] rrespDecoder; // @[OneHot.scala 45:35:@104928.4]
  wire [255:0] wrespDecoder; // @[OneHot.scala 45:35:@104929.4]
  wire  _T_479; // @[StreamArbiter.scala 61:55:@104934.4]
  wire  _T_486; // @[StreamArbiter.scala 64:58:@104943.4]
  wire  _T_490; // @[StreamArbiter.scala 61:55:@105015.4]
  wire  _T_493; // @[StreamArbiter.scala 62:85:@105019.4]
  wire  _T_494; // @[StreamArbiter.scala 62:70:@105020.4]
  wire  _T_499; // @[StreamArbiter.scala 67:58:@105092.4]
  wire  _T_510; // @[:@105099.4]
  wire  _T_520; // @[:@105104.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@104427.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@104434.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  MuxPipe cmdMux ( // @[StreamArbiter.scala 25:22:@104444.4]
    .io_in_ready(cmdMux_io_in_ready),
    .io_in_valid(cmdMux_io_in_valid),
    .io_in_bits_0_addr(cmdMux_io_in_bits_0_addr),
    .io_in_bits_0_size(cmdMux_io_in_bits_0_size),
    .io_in_bits_1_addr(cmdMux_io_in_bits_1_addr),
    .io_in_bits_1_size(cmdMux_io_in_bits_1_size),
    .io_sel(cmdMux_io_sel),
    .io_out_ready(cmdMux_io_out_ready),
    .io_out_valid(cmdMux_io_out_valid),
    .io_out_bits_addr(cmdMux_io_out_bits_addr),
    .io_out_bits_size(cmdMux_io_out_bits_size),
    .io_out_bits_isWr(cmdMux_io_out_bits_isWr),
    .io_out_bits_tag(cmdMux_io_out_bits_tag)
  );
  MuxPipe_1 wdataMux ( // @[StreamArbiter.scala 35:24:@104486.4]
    .io_in_ready(wdataMux_io_in_ready),
    .io_in_valid(wdataMux_io_in_valid),
    .io_in_bits_1_wdata_0(wdataMux_io_in_bits_1_wdata_0),
    .io_in_bits_1_wdata_1(wdataMux_io_in_bits_1_wdata_1),
    .io_in_bits_1_wdata_2(wdataMux_io_in_bits_1_wdata_2),
    .io_in_bits_1_wdata_3(wdataMux_io_in_bits_1_wdata_3),
    .io_in_bits_1_wdata_4(wdataMux_io_in_bits_1_wdata_4),
    .io_in_bits_1_wdata_5(wdataMux_io_in_bits_1_wdata_5),
    .io_in_bits_1_wdata_6(wdataMux_io_in_bits_1_wdata_6),
    .io_in_bits_1_wdata_7(wdataMux_io_in_bits_1_wdata_7),
    .io_in_bits_1_wdata_8(wdataMux_io_in_bits_1_wdata_8),
    .io_in_bits_1_wdata_9(wdataMux_io_in_bits_1_wdata_9),
    .io_in_bits_1_wdata_10(wdataMux_io_in_bits_1_wdata_10),
    .io_in_bits_1_wdata_11(wdataMux_io_in_bits_1_wdata_11),
    .io_in_bits_1_wdata_12(wdataMux_io_in_bits_1_wdata_12),
    .io_in_bits_1_wdata_13(wdataMux_io_in_bits_1_wdata_13),
    .io_in_bits_1_wdata_14(wdataMux_io_in_bits_1_wdata_14),
    .io_in_bits_1_wdata_15(wdataMux_io_in_bits_1_wdata_15),
    .io_in_bits_1_wdata_16(wdataMux_io_in_bits_1_wdata_16),
    .io_in_bits_1_wdata_17(wdataMux_io_in_bits_1_wdata_17),
    .io_in_bits_1_wdata_18(wdataMux_io_in_bits_1_wdata_18),
    .io_in_bits_1_wdata_19(wdataMux_io_in_bits_1_wdata_19),
    .io_in_bits_1_wdata_20(wdataMux_io_in_bits_1_wdata_20),
    .io_in_bits_1_wdata_21(wdataMux_io_in_bits_1_wdata_21),
    .io_in_bits_1_wdata_22(wdataMux_io_in_bits_1_wdata_22),
    .io_in_bits_1_wdata_23(wdataMux_io_in_bits_1_wdata_23),
    .io_in_bits_1_wdata_24(wdataMux_io_in_bits_1_wdata_24),
    .io_in_bits_1_wdata_25(wdataMux_io_in_bits_1_wdata_25),
    .io_in_bits_1_wdata_26(wdataMux_io_in_bits_1_wdata_26),
    .io_in_bits_1_wdata_27(wdataMux_io_in_bits_1_wdata_27),
    .io_in_bits_1_wdata_28(wdataMux_io_in_bits_1_wdata_28),
    .io_in_bits_1_wdata_29(wdataMux_io_in_bits_1_wdata_29),
    .io_in_bits_1_wdata_30(wdataMux_io_in_bits_1_wdata_30),
    .io_in_bits_1_wdata_31(wdataMux_io_in_bits_1_wdata_31),
    .io_in_bits_1_wdata_32(wdataMux_io_in_bits_1_wdata_32),
    .io_in_bits_1_wdata_33(wdataMux_io_in_bits_1_wdata_33),
    .io_in_bits_1_wdata_34(wdataMux_io_in_bits_1_wdata_34),
    .io_in_bits_1_wdata_35(wdataMux_io_in_bits_1_wdata_35),
    .io_in_bits_1_wdata_36(wdataMux_io_in_bits_1_wdata_36),
    .io_in_bits_1_wdata_37(wdataMux_io_in_bits_1_wdata_37),
    .io_in_bits_1_wdata_38(wdataMux_io_in_bits_1_wdata_38),
    .io_in_bits_1_wdata_39(wdataMux_io_in_bits_1_wdata_39),
    .io_in_bits_1_wdata_40(wdataMux_io_in_bits_1_wdata_40),
    .io_in_bits_1_wdata_41(wdataMux_io_in_bits_1_wdata_41),
    .io_in_bits_1_wdata_42(wdataMux_io_in_bits_1_wdata_42),
    .io_in_bits_1_wdata_43(wdataMux_io_in_bits_1_wdata_43),
    .io_in_bits_1_wdata_44(wdataMux_io_in_bits_1_wdata_44),
    .io_in_bits_1_wdata_45(wdataMux_io_in_bits_1_wdata_45),
    .io_in_bits_1_wdata_46(wdataMux_io_in_bits_1_wdata_46),
    .io_in_bits_1_wdata_47(wdataMux_io_in_bits_1_wdata_47),
    .io_in_bits_1_wdata_48(wdataMux_io_in_bits_1_wdata_48),
    .io_in_bits_1_wdata_49(wdataMux_io_in_bits_1_wdata_49),
    .io_in_bits_1_wdata_50(wdataMux_io_in_bits_1_wdata_50),
    .io_in_bits_1_wdata_51(wdataMux_io_in_bits_1_wdata_51),
    .io_in_bits_1_wdata_52(wdataMux_io_in_bits_1_wdata_52),
    .io_in_bits_1_wdata_53(wdataMux_io_in_bits_1_wdata_53),
    .io_in_bits_1_wdata_54(wdataMux_io_in_bits_1_wdata_54),
    .io_in_bits_1_wdata_55(wdataMux_io_in_bits_1_wdata_55),
    .io_in_bits_1_wdata_56(wdataMux_io_in_bits_1_wdata_56),
    .io_in_bits_1_wdata_57(wdataMux_io_in_bits_1_wdata_57),
    .io_in_bits_1_wdata_58(wdataMux_io_in_bits_1_wdata_58),
    .io_in_bits_1_wdata_59(wdataMux_io_in_bits_1_wdata_59),
    .io_in_bits_1_wdata_60(wdataMux_io_in_bits_1_wdata_60),
    .io_in_bits_1_wdata_61(wdataMux_io_in_bits_1_wdata_61),
    .io_in_bits_1_wdata_62(wdataMux_io_in_bits_1_wdata_62),
    .io_in_bits_1_wdata_63(wdataMux_io_in_bits_1_wdata_63),
    .io_in_bits_1_wstrb_0(wdataMux_io_in_bits_1_wstrb_0),
    .io_in_bits_1_wstrb_1(wdataMux_io_in_bits_1_wstrb_1),
    .io_in_bits_1_wstrb_2(wdataMux_io_in_bits_1_wstrb_2),
    .io_in_bits_1_wstrb_3(wdataMux_io_in_bits_1_wstrb_3),
    .io_in_bits_1_wstrb_4(wdataMux_io_in_bits_1_wstrb_4),
    .io_in_bits_1_wstrb_5(wdataMux_io_in_bits_1_wstrb_5),
    .io_in_bits_1_wstrb_6(wdataMux_io_in_bits_1_wstrb_6),
    .io_in_bits_1_wstrb_7(wdataMux_io_in_bits_1_wstrb_7),
    .io_in_bits_1_wstrb_8(wdataMux_io_in_bits_1_wstrb_8),
    .io_in_bits_1_wstrb_9(wdataMux_io_in_bits_1_wstrb_9),
    .io_in_bits_1_wstrb_10(wdataMux_io_in_bits_1_wstrb_10),
    .io_in_bits_1_wstrb_11(wdataMux_io_in_bits_1_wstrb_11),
    .io_in_bits_1_wstrb_12(wdataMux_io_in_bits_1_wstrb_12),
    .io_in_bits_1_wstrb_13(wdataMux_io_in_bits_1_wstrb_13),
    .io_in_bits_1_wstrb_14(wdataMux_io_in_bits_1_wstrb_14),
    .io_in_bits_1_wstrb_15(wdataMux_io_in_bits_1_wstrb_15),
    .io_in_bits_1_wstrb_16(wdataMux_io_in_bits_1_wstrb_16),
    .io_in_bits_1_wstrb_17(wdataMux_io_in_bits_1_wstrb_17),
    .io_in_bits_1_wstrb_18(wdataMux_io_in_bits_1_wstrb_18),
    .io_in_bits_1_wstrb_19(wdataMux_io_in_bits_1_wstrb_19),
    .io_in_bits_1_wstrb_20(wdataMux_io_in_bits_1_wstrb_20),
    .io_in_bits_1_wstrb_21(wdataMux_io_in_bits_1_wstrb_21),
    .io_in_bits_1_wstrb_22(wdataMux_io_in_bits_1_wstrb_22),
    .io_in_bits_1_wstrb_23(wdataMux_io_in_bits_1_wstrb_23),
    .io_in_bits_1_wstrb_24(wdataMux_io_in_bits_1_wstrb_24),
    .io_in_bits_1_wstrb_25(wdataMux_io_in_bits_1_wstrb_25),
    .io_in_bits_1_wstrb_26(wdataMux_io_in_bits_1_wstrb_26),
    .io_in_bits_1_wstrb_27(wdataMux_io_in_bits_1_wstrb_27),
    .io_in_bits_1_wstrb_28(wdataMux_io_in_bits_1_wstrb_28),
    .io_in_bits_1_wstrb_29(wdataMux_io_in_bits_1_wstrb_29),
    .io_in_bits_1_wstrb_30(wdataMux_io_in_bits_1_wstrb_30),
    .io_in_bits_1_wstrb_31(wdataMux_io_in_bits_1_wstrb_31),
    .io_in_bits_1_wstrb_32(wdataMux_io_in_bits_1_wstrb_32),
    .io_in_bits_1_wstrb_33(wdataMux_io_in_bits_1_wstrb_33),
    .io_in_bits_1_wstrb_34(wdataMux_io_in_bits_1_wstrb_34),
    .io_in_bits_1_wstrb_35(wdataMux_io_in_bits_1_wstrb_35),
    .io_in_bits_1_wstrb_36(wdataMux_io_in_bits_1_wstrb_36),
    .io_in_bits_1_wstrb_37(wdataMux_io_in_bits_1_wstrb_37),
    .io_in_bits_1_wstrb_38(wdataMux_io_in_bits_1_wstrb_38),
    .io_in_bits_1_wstrb_39(wdataMux_io_in_bits_1_wstrb_39),
    .io_in_bits_1_wstrb_40(wdataMux_io_in_bits_1_wstrb_40),
    .io_in_bits_1_wstrb_41(wdataMux_io_in_bits_1_wstrb_41),
    .io_in_bits_1_wstrb_42(wdataMux_io_in_bits_1_wstrb_42),
    .io_in_bits_1_wstrb_43(wdataMux_io_in_bits_1_wstrb_43),
    .io_in_bits_1_wstrb_44(wdataMux_io_in_bits_1_wstrb_44),
    .io_in_bits_1_wstrb_45(wdataMux_io_in_bits_1_wstrb_45),
    .io_in_bits_1_wstrb_46(wdataMux_io_in_bits_1_wstrb_46),
    .io_in_bits_1_wstrb_47(wdataMux_io_in_bits_1_wstrb_47),
    .io_in_bits_1_wstrb_48(wdataMux_io_in_bits_1_wstrb_48),
    .io_in_bits_1_wstrb_49(wdataMux_io_in_bits_1_wstrb_49),
    .io_in_bits_1_wstrb_50(wdataMux_io_in_bits_1_wstrb_50),
    .io_in_bits_1_wstrb_51(wdataMux_io_in_bits_1_wstrb_51),
    .io_in_bits_1_wstrb_52(wdataMux_io_in_bits_1_wstrb_52),
    .io_in_bits_1_wstrb_53(wdataMux_io_in_bits_1_wstrb_53),
    .io_in_bits_1_wstrb_54(wdataMux_io_in_bits_1_wstrb_54),
    .io_in_bits_1_wstrb_55(wdataMux_io_in_bits_1_wstrb_55),
    .io_in_bits_1_wstrb_56(wdataMux_io_in_bits_1_wstrb_56),
    .io_in_bits_1_wstrb_57(wdataMux_io_in_bits_1_wstrb_57),
    .io_in_bits_1_wstrb_58(wdataMux_io_in_bits_1_wstrb_58),
    .io_in_bits_1_wstrb_59(wdataMux_io_in_bits_1_wstrb_59),
    .io_in_bits_1_wstrb_60(wdataMux_io_in_bits_1_wstrb_60),
    .io_in_bits_1_wstrb_61(wdataMux_io_in_bits_1_wstrb_61),
    .io_in_bits_1_wstrb_62(wdataMux_io_in_bits_1_wstrb_62),
    .io_in_bits_1_wstrb_63(wdataMux_io_in_bits_1_wstrb_63),
    .io_sel(wdataMux_io_sel),
    .io_out_ready(wdataMux_io_out_ready),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wdata_8(wdataMux_io_out_bits_wdata_8),
    .io_out_bits_wdata_9(wdataMux_io_out_bits_wdata_9),
    .io_out_bits_wdata_10(wdataMux_io_out_bits_wdata_10),
    .io_out_bits_wdata_11(wdataMux_io_out_bits_wdata_11),
    .io_out_bits_wdata_12(wdataMux_io_out_bits_wdata_12),
    .io_out_bits_wdata_13(wdataMux_io_out_bits_wdata_13),
    .io_out_bits_wdata_14(wdataMux_io_out_bits_wdata_14),
    .io_out_bits_wdata_15(wdataMux_io_out_bits_wdata_15),
    .io_out_bits_wdata_16(wdataMux_io_out_bits_wdata_16),
    .io_out_bits_wdata_17(wdataMux_io_out_bits_wdata_17),
    .io_out_bits_wdata_18(wdataMux_io_out_bits_wdata_18),
    .io_out_bits_wdata_19(wdataMux_io_out_bits_wdata_19),
    .io_out_bits_wdata_20(wdataMux_io_out_bits_wdata_20),
    .io_out_bits_wdata_21(wdataMux_io_out_bits_wdata_21),
    .io_out_bits_wdata_22(wdataMux_io_out_bits_wdata_22),
    .io_out_bits_wdata_23(wdataMux_io_out_bits_wdata_23),
    .io_out_bits_wdata_24(wdataMux_io_out_bits_wdata_24),
    .io_out_bits_wdata_25(wdataMux_io_out_bits_wdata_25),
    .io_out_bits_wdata_26(wdataMux_io_out_bits_wdata_26),
    .io_out_bits_wdata_27(wdataMux_io_out_bits_wdata_27),
    .io_out_bits_wdata_28(wdataMux_io_out_bits_wdata_28),
    .io_out_bits_wdata_29(wdataMux_io_out_bits_wdata_29),
    .io_out_bits_wdata_30(wdataMux_io_out_bits_wdata_30),
    .io_out_bits_wdata_31(wdataMux_io_out_bits_wdata_31),
    .io_out_bits_wdata_32(wdataMux_io_out_bits_wdata_32),
    .io_out_bits_wdata_33(wdataMux_io_out_bits_wdata_33),
    .io_out_bits_wdata_34(wdataMux_io_out_bits_wdata_34),
    .io_out_bits_wdata_35(wdataMux_io_out_bits_wdata_35),
    .io_out_bits_wdata_36(wdataMux_io_out_bits_wdata_36),
    .io_out_bits_wdata_37(wdataMux_io_out_bits_wdata_37),
    .io_out_bits_wdata_38(wdataMux_io_out_bits_wdata_38),
    .io_out_bits_wdata_39(wdataMux_io_out_bits_wdata_39),
    .io_out_bits_wdata_40(wdataMux_io_out_bits_wdata_40),
    .io_out_bits_wdata_41(wdataMux_io_out_bits_wdata_41),
    .io_out_bits_wdata_42(wdataMux_io_out_bits_wdata_42),
    .io_out_bits_wdata_43(wdataMux_io_out_bits_wdata_43),
    .io_out_bits_wdata_44(wdataMux_io_out_bits_wdata_44),
    .io_out_bits_wdata_45(wdataMux_io_out_bits_wdata_45),
    .io_out_bits_wdata_46(wdataMux_io_out_bits_wdata_46),
    .io_out_bits_wdata_47(wdataMux_io_out_bits_wdata_47),
    .io_out_bits_wdata_48(wdataMux_io_out_bits_wdata_48),
    .io_out_bits_wdata_49(wdataMux_io_out_bits_wdata_49),
    .io_out_bits_wdata_50(wdataMux_io_out_bits_wdata_50),
    .io_out_bits_wdata_51(wdataMux_io_out_bits_wdata_51),
    .io_out_bits_wdata_52(wdataMux_io_out_bits_wdata_52),
    .io_out_bits_wdata_53(wdataMux_io_out_bits_wdata_53),
    .io_out_bits_wdata_54(wdataMux_io_out_bits_wdata_54),
    .io_out_bits_wdata_55(wdataMux_io_out_bits_wdata_55),
    .io_out_bits_wdata_56(wdataMux_io_out_bits_wdata_56),
    .io_out_bits_wdata_57(wdataMux_io_out_bits_wdata_57),
    .io_out_bits_wdata_58(wdataMux_io_out_bits_wdata_58),
    .io_out_bits_wdata_59(wdataMux_io_out_bits_wdata_59),
    .io_out_bits_wdata_60(wdataMux_io_out_bits_wdata_60),
    .io_out_bits_wdata_61(wdataMux_io_out_bits_wdata_61),
    .io_out_bits_wdata_62(wdataMux_io_out_bits_wdata_62),
    .io_out_bits_wdata_63(wdataMux_io_out_bits_wdata_63),
    .io_out_bits_wstrb_0(wdataMux_io_out_bits_wstrb_0),
    .io_out_bits_wstrb_1(wdataMux_io_out_bits_wstrb_1),
    .io_out_bits_wstrb_2(wdataMux_io_out_bits_wstrb_2),
    .io_out_bits_wstrb_3(wdataMux_io_out_bits_wstrb_3),
    .io_out_bits_wstrb_4(wdataMux_io_out_bits_wstrb_4),
    .io_out_bits_wstrb_5(wdataMux_io_out_bits_wstrb_5),
    .io_out_bits_wstrb_6(wdataMux_io_out_bits_wstrb_6),
    .io_out_bits_wstrb_7(wdataMux_io_out_bits_wstrb_7),
    .io_out_bits_wstrb_8(wdataMux_io_out_bits_wstrb_8),
    .io_out_bits_wstrb_9(wdataMux_io_out_bits_wstrb_9),
    .io_out_bits_wstrb_10(wdataMux_io_out_bits_wstrb_10),
    .io_out_bits_wstrb_11(wdataMux_io_out_bits_wstrb_11),
    .io_out_bits_wstrb_12(wdataMux_io_out_bits_wstrb_12),
    .io_out_bits_wstrb_13(wdataMux_io_out_bits_wstrb_13),
    .io_out_bits_wstrb_14(wdataMux_io_out_bits_wstrb_14),
    .io_out_bits_wstrb_15(wdataMux_io_out_bits_wstrb_15),
    .io_out_bits_wstrb_16(wdataMux_io_out_bits_wstrb_16),
    .io_out_bits_wstrb_17(wdataMux_io_out_bits_wstrb_17),
    .io_out_bits_wstrb_18(wdataMux_io_out_bits_wstrb_18),
    .io_out_bits_wstrb_19(wdataMux_io_out_bits_wstrb_19),
    .io_out_bits_wstrb_20(wdataMux_io_out_bits_wstrb_20),
    .io_out_bits_wstrb_21(wdataMux_io_out_bits_wstrb_21),
    .io_out_bits_wstrb_22(wdataMux_io_out_bits_wstrb_22),
    .io_out_bits_wstrb_23(wdataMux_io_out_bits_wstrb_23),
    .io_out_bits_wstrb_24(wdataMux_io_out_bits_wstrb_24),
    .io_out_bits_wstrb_25(wdataMux_io_out_bits_wstrb_25),
    .io_out_bits_wstrb_26(wdataMux_io_out_bits_wstrb_26),
    .io_out_bits_wstrb_27(wdataMux_io_out_bits_wstrb_27),
    .io_out_bits_wstrb_28(wdataMux_io_out_bits_wstrb_28),
    .io_out_bits_wstrb_29(wdataMux_io_out_bits_wstrb_29),
    .io_out_bits_wstrb_30(wdataMux_io_out_bits_wstrb_30),
    .io_out_bits_wstrb_31(wdataMux_io_out_bits_wstrb_31),
    .io_out_bits_wstrb_32(wdataMux_io_out_bits_wstrb_32),
    .io_out_bits_wstrb_33(wdataMux_io_out_bits_wstrb_33),
    .io_out_bits_wstrb_34(wdataMux_io_out_bits_wstrb_34),
    .io_out_bits_wstrb_35(wdataMux_io_out_bits_wstrb_35),
    .io_out_bits_wstrb_36(wdataMux_io_out_bits_wstrb_36),
    .io_out_bits_wstrb_37(wdataMux_io_out_bits_wstrb_37),
    .io_out_bits_wstrb_38(wdataMux_io_out_bits_wstrb_38),
    .io_out_bits_wstrb_39(wdataMux_io_out_bits_wstrb_39),
    .io_out_bits_wstrb_40(wdataMux_io_out_bits_wstrb_40),
    .io_out_bits_wstrb_41(wdataMux_io_out_bits_wstrb_41),
    .io_out_bits_wstrb_42(wdataMux_io_out_bits_wstrb_42),
    .io_out_bits_wstrb_43(wdataMux_io_out_bits_wstrb_43),
    .io_out_bits_wstrb_44(wdataMux_io_out_bits_wstrb_44),
    .io_out_bits_wstrb_45(wdataMux_io_out_bits_wstrb_45),
    .io_out_bits_wstrb_46(wdataMux_io_out_bits_wstrb_46),
    .io_out_bits_wstrb_47(wdataMux_io_out_bits_wstrb_47),
    .io_out_bits_wstrb_48(wdataMux_io_out_bits_wstrb_48),
    .io_out_bits_wstrb_49(wdataMux_io_out_bits_wstrb_49),
    .io_out_bits_wstrb_50(wdataMux_io_out_bits_wstrb_50),
    .io_out_bits_wstrb_51(wdataMux_io_out_bits_wstrb_51),
    .io_out_bits_wstrb_52(wdataMux_io_out_bits_wstrb_52),
    .io_out_bits_wstrb_53(wdataMux_io_out_bits_wstrb_53),
    .io_out_bits_wstrb_54(wdataMux_io_out_bits_wstrb_54),
    .io_out_bits_wstrb_55(wdataMux_io_out_bits_wstrb_55),
    .io_out_bits_wstrb_56(wdataMux_io_out_bits_wstrb_56),
    .io_out_bits_wstrb_57(wdataMux_io_out_bits_wstrb_57),
    .io_out_bits_wstrb_58(wdataMux_io_out_bits_wstrb_58),
    .io_out_bits_wstrb_59(wdataMux_io_out_bits_wstrb_59),
    .io_out_bits_wstrb_60(wdataMux_io_out_bits_wstrb_60),
    .io_out_bits_wstrb_61(wdataMux_io_out_bits_wstrb_61),
    .io_out_bits_wstrb_62(wdataMux_io_out_bits_wstrb_62),
    .io_out_bits_wstrb_63(wdataMux_io_out_bits_wstrb_63)
  );
  ElementCounter elementCtr ( // @[StreamArbiter.scala 36:26:@104489.4]
    .clock(elementCtr_clock),
    .reset(elementCtr_reset),
    .io_reset(elementCtr_io_reset),
    .io_enable(elementCtr_io_enable),
    .io_out(elementCtr_io_out)
  );
  assign priorityActive = io_app_0_cmd_valid ? 1'h0 : 1'h1; // @[Mux.scala 31:69:@104422.4]
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@104432.4 package.scala 96:25:@104433.4]
  assign _GEN_1 = _T_408 ? io_app_1_cmd_valid : io_app_0_cmd_valid; // @[StreamArbiter.scala 21:16:@104441.4]
  assign _T_412 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@104439.4 package.scala 96:25:@104440.4]
  assign cmdIdx = _GEN_1 ? _T_412 : priorityActive; // @[StreamArbiter.scala 21:16:@104441.4]
  assign cmdInDecoder = 2'h1 << cmdIdx; // @[OneHot.scala 45:35:@104443.4]
  assign _T_438 = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:49:@104492.4]
  assign _T_443 = cmdMux_io_out_bits_tag; // @[:@104496.4 :@104497.4]
  assign _T_444 = _T_443[7:0]; // @[FringeBundles.scala 114:28:@104498.4]
  assign cmdOutDecoder = 256'h1 << _T_444; // @[OneHot.scala 45:35:@104504.4]
  assign _T_457 = _T_444[0]; // @[:@104508.4]
  assign _GEN_3 = _T_457 ? io_app_1_wdata_valid : 1'h0; // @[StreamArbiter.scala 42:78:@104509.4]
  assign _T_458 = _GEN_3 & cmdMux_io_out_valid; // @[StreamArbiter.scala 42:78:@104509.4]
  assign _T_459 = elementCtr_io_out < cmdMux_io_out_bits_size; // @[StreamArbiter.scala 42:121:@104510.4]
  assign _T_466 = io_dram_rresp_bits_tag[7:0]; // @[FringeBundles.scala 132:28:@104913.4]
  assign _T_474 = io_dram_wresp_bits_tag[7:0]; // @[FringeBundles.scala 140:28:@104922.4]
  assign rrespDecoder = 256'h1 << _T_466; // @[OneHot.scala 45:35:@104928.4]
  assign wrespDecoder = 256'h1 << _T_474; // @[OneHot.scala 45:35:@104929.4]
  assign _T_479 = cmdInDecoder[0]; // @[StreamArbiter.scala 61:55:@104934.4]
  assign _T_486 = rrespDecoder[0]; // @[StreamArbiter.scala 64:58:@104943.4]
  assign _T_490 = cmdInDecoder[1]; // @[StreamArbiter.scala 61:55:@105015.4]
  assign _T_493 = cmdOutDecoder[1]; // @[StreamArbiter.scala 62:85:@105019.4]
  assign _T_494 = _T_438 & _T_493; // @[StreamArbiter.scala 62:70:@105020.4]
  assign _T_499 = wrespDecoder[1]; // @[StreamArbiter.scala 67:58:@105092.4]
  assign _T_510 = _T_466[0]; // @[:@105099.4]
  assign _T_520 = _T_474[0]; // @[:@105104.4]
  assign io_app_0_cmd_ready = cmdMux_io_in_ready & _T_479; // @[StreamArbiter.scala 61:19:@104936.4]
  assign io_app_0_rresp_valid = io_dram_rresp_valid & _T_486; // @[StreamArbiter.scala 64:21:@104945.4]
  assign io_app_0_rresp_bits_rdata_0 = io_dram_rresp_bits_rdata_0; // @[StreamArbiter.scala 65:20:@104947.4]
  assign io_app_0_rresp_bits_rdata_1 = io_dram_rresp_bits_rdata_1; // @[StreamArbiter.scala 65:20:@104948.4]
  assign io_app_0_rresp_bits_rdata_2 = io_dram_rresp_bits_rdata_2; // @[StreamArbiter.scala 65:20:@104949.4]
  assign io_app_0_rresp_bits_rdata_3 = io_dram_rresp_bits_rdata_3; // @[StreamArbiter.scala 65:20:@104950.4]
  assign io_app_0_rresp_bits_rdata_4 = io_dram_rresp_bits_rdata_4; // @[StreamArbiter.scala 65:20:@104951.4]
  assign io_app_0_rresp_bits_rdata_5 = io_dram_rresp_bits_rdata_5; // @[StreamArbiter.scala 65:20:@104952.4]
  assign io_app_0_rresp_bits_rdata_6 = io_dram_rresp_bits_rdata_6; // @[StreamArbiter.scala 65:20:@104953.4]
  assign io_app_0_rresp_bits_rdata_7 = io_dram_rresp_bits_rdata_7; // @[StreamArbiter.scala 65:20:@104954.4]
  assign io_app_0_rresp_bits_rdata_8 = io_dram_rresp_bits_rdata_8; // @[StreamArbiter.scala 65:20:@104955.4]
  assign io_app_0_rresp_bits_rdata_9 = io_dram_rresp_bits_rdata_9; // @[StreamArbiter.scala 65:20:@104956.4]
  assign io_app_0_rresp_bits_rdata_10 = io_dram_rresp_bits_rdata_10; // @[StreamArbiter.scala 65:20:@104957.4]
  assign io_app_0_rresp_bits_rdata_11 = io_dram_rresp_bits_rdata_11; // @[StreamArbiter.scala 65:20:@104958.4]
  assign io_app_0_rresp_bits_rdata_12 = io_dram_rresp_bits_rdata_12; // @[StreamArbiter.scala 65:20:@104959.4]
  assign io_app_0_rresp_bits_rdata_13 = io_dram_rresp_bits_rdata_13; // @[StreamArbiter.scala 65:20:@104960.4]
  assign io_app_0_rresp_bits_rdata_14 = io_dram_rresp_bits_rdata_14; // @[StreamArbiter.scala 65:20:@104961.4]
  assign io_app_0_rresp_bits_rdata_15 = io_dram_rresp_bits_rdata_15; // @[StreamArbiter.scala 65:20:@104962.4]
  assign io_app_0_rresp_bits_rdata_16 = io_dram_rresp_bits_rdata_16; // @[StreamArbiter.scala 65:20:@104963.4]
  assign io_app_0_rresp_bits_rdata_17 = io_dram_rresp_bits_rdata_17; // @[StreamArbiter.scala 65:20:@104964.4]
  assign io_app_0_rresp_bits_rdata_18 = io_dram_rresp_bits_rdata_18; // @[StreamArbiter.scala 65:20:@104965.4]
  assign io_app_0_rresp_bits_rdata_19 = io_dram_rresp_bits_rdata_19; // @[StreamArbiter.scala 65:20:@104966.4]
  assign io_app_0_rresp_bits_rdata_20 = io_dram_rresp_bits_rdata_20; // @[StreamArbiter.scala 65:20:@104967.4]
  assign io_app_0_rresp_bits_rdata_21 = io_dram_rresp_bits_rdata_21; // @[StreamArbiter.scala 65:20:@104968.4]
  assign io_app_0_rresp_bits_rdata_22 = io_dram_rresp_bits_rdata_22; // @[StreamArbiter.scala 65:20:@104969.4]
  assign io_app_0_rresp_bits_rdata_23 = io_dram_rresp_bits_rdata_23; // @[StreamArbiter.scala 65:20:@104970.4]
  assign io_app_0_rresp_bits_rdata_24 = io_dram_rresp_bits_rdata_24; // @[StreamArbiter.scala 65:20:@104971.4]
  assign io_app_0_rresp_bits_rdata_25 = io_dram_rresp_bits_rdata_25; // @[StreamArbiter.scala 65:20:@104972.4]
  assign io_app_0_rresp_bits_rdata_26 = io_dram_rresp_bits_rdata_26; // @[StreamArbiter.scala 65:20:@104973.4]
  assign io_app_0_rresp_bits_rdata_27 = io_dram_rresp_bits_rdata_27; // @[StreamArbiter.scala 65:20:@104974.4]
  assign io_app_0_rresp_bits_rdata_28 = io_dram_rresp_bits_rdata_28; // @[StreamArbiter.scala 65:20:@104975.4]
  assign io_app_0_rresp_bits_rdata_29 = io_dram_rresp_bits_rdata_29; // @[StreamArbiter.scala 65:20:@104976.4]
  assign io_app_0_rresp_bits_rdata_30 = io_dram_rresp_bits_rdata_30; // @[StreamArbiter.scala 65:20:@104977.4]
  assign io_app_0_rresp_bits_rdata_31 = io_dram_rresp_bits_rdata_31; // @[StreamArbiter.scala 65:20:@104978.4]
  assign io_app_0_rresp_bits_rdata_32 = io_dram_rresp_bits_rdata_32; // @[StreamArbiter.scala 65:20:@104979.4]
  assign io_app_0_rresp_bits_rdata_33 = io_dram_rresp_bits_rdata_33; // @[StreamArbiter.scala 65:20:@104980.4]
  assign io_app_0_rresp_bits_rdata_34 = io_dram_rresp_bits_rdata_34; // @[StreamArbiter.scala 65:20:@104981.4]
  assign io_app_0_rresp_bits_rdata_35 = io_dram_rresp_bits_rdata_35; // @[StreamArbiter.scala 65:20:@104982.4]
  assign io_app_0_rresp_bits_rdata_36 = io_dram_rresp_bits_rdata_36; // @[StreamArbiter.scala 65:20:@104983.4]
  assign io_app_0_rresp_bits_rdata_37 = io_dram_rresp_bits_rdata_37; // @[StreamArbiter.scala 65:20:@104984.4]
  assign io_app_0_rresp_bits_rdata_38 = io_dram_rresp_bits_rdata_38; // @[StreamArbiter.scala 65:20:@104985.4]
  assign io_app_0_rresp_bits_rdata_39 = io_dram_rresp_bits_rdata_39; // @[StreamArbiter.scala 65:20:@104986.4]
  assign io_app_0_rresp_bits_rdata_40 = io_dram_rresp_bits_rdata_40; // @[StreamArbiter.scala 65:20:@104987.4]
  assign io_app_0_rresp_bits_rdata_41 = io_dram_rresp_bits_rdata_41; // @[StreamArbiter.scala 65:20:@104988.4]
  assign io_app_0_rresp_bits_rdata_42 = io_dram_rresp_bits_rdata_42; // @[StreamArbiter.scala 65:20:@104989.4]
  assign io_app_0_rresp_bits_rdata_43 = io_dram_rresp_bits_rdata_43; // @[StreamArbiter.scala 65:20:@104990.4]
  assign io_app_0_rresp_bits_rdata_44 = io_dram_rresp_bits_rdata_44; // @[StreamArbiter.scala 65:20:@104991.4]
  assign io_app_0_rresp_bits_rdata_45 = io_dram_rresp_bits_rdata_45; // @[StreamArbiter.scala 65:20:@104992.4]
  assign io_app_0_rresp_bits_rdata_46 = io_dram_rresp_bits_rdata_46; // @[StreamArbiter.scala 65:20:@104993.4]
  assign io_app_0_rresp_bits_rdata_47 = io_dram_rresp_bits_rdata_47; // @[StreamArbiter.scala 65:20:@104994.4]
  assign io_app_0_rresp_bits_rdata_48 = io_dram_rresp_bits_rdata_48; // @[StreamArbiter.scala 65:20:@104995.4]
  assign io_app_0_rresp_bits_rdata_49 = io_dram_rresp_bits_rdata_49; // @[StreamArbiter.scala 65:20:@104996.4]
  assign io_app_0_rresp_bits_rdata_50 = io_dram_rresp_bits_rdata_50; // @[StreamArbiter.scala 65:20:@104997.4]
  assign io_app_0_rresp_bits_rdata_51 = io_dram_rresp_bits_rdata_51; // @[StreamArbiter.scala 65:20:@104998.4]
  assign io_app_0_rresp_bits_rdata_52 = io_dram_rresp_bits_rdata_52; // @[StreamArbiter.scala 65:20:@104999.4]
  assign io_app_0_rresp_bits_rdata_53 = io_dram_rresp_bits_rdata_53; // @[StreamArbiter.scala 65:20:@105000.4]
  assign io_app_0_rresp_bits_rdata_54 = io_dram_rresp_bits_rdata_54; // @[StreamArbiter.scala 65:20:@105001.4]
  assign io_app_0_rresp_bits_rdata_55 = io_dram_rresp_bits_rdata_55; // @[StreamArbiter.scala 65:20:@105002.4]
  assign io_app_0_rresp_bits_rdata_56 = io_dram_rresp_bits_rdata_56; // @[StreamArbiter.scala 65:20:@105003.4]
  assign io_app_0_rresp_bits_rdata_57 = io_dram_rresp_bits_rdata_57; // @[StreamArbiter.scala 65:20:@105004.4]
  assign io_app_0_rresp_bits_rdata_58 = io_dram_rresp_bits_rdata_58; // @[StreamArbiter.scala 65:20:@105005.4]
  assign io_app_0_rresp_bits_rdata_59 = io_dram_rresp_bits_rdata_59; // @[StreamArbiter.scala 65:20:@105006.4]
  assign io_app_0_rresp_bits_rdata_60 = io_dram_rresp_bits_rdata_60; // @[StreamArbiter.scala 65:20:@105007.4]
  assign io_app_0_rresp_bits_rdata_61 = io_dram_rresp_bits_rdata_61; // @[StreamArbiter.scala 65:20:@105008.4]
  assign io_app_0_rresp_bits_rdata_62 = io_dram_rresp_bits_rdata_62; // @[StreamArbiter.scala 65:20:@105009.4]
  assign io_app_0_rresp_bits_rdata_63 = io_dram_rresp_bits_rdata_63; // @[StreamArbiter.scala 65:20:@105010.4]
  assign io_app_1_cmd_ready = cmdMux_io_in_ready & _T_490; // @[StreamArbiter.scala 61:19:@105017.4]
  assign io_app_1_wdata_ready = _T_494 & _T_459; // @[StreamArbiter.scala 62:21:@105023.4]
  assign io_app_1_wresp_valid = io_dram_wresp_valid & _T_499; // @[StreamArbiter.scala 67:21:@105094.4]
  assign io_dram_cmd_valid = cmdMux_io_out_valid; // @[StreamArbiter.scala 46:15:@104777.4]
  assign io_dram_cmd_bits_addr = cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 46:15:@104776.4]
  assign io_dram_cmd_bits_size = cmdMux_io_out_bits_size; // @[StreamArbiter.scala 46:15:@104775.4]
  assign io_dram_cmd_bits_isWr = cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 46:15:@104773.4]
  assign io_dram_cmd_bits_tag = cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 46:15:@104772.4]
  assign io_dram_wdata_valid = wdataMux_io_out_valid; // @[StreamArbiter.scala 47:17:@104908.4]
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 47:17:@104844.4]
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 47:17:@104845.4]
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 47:17:@104846.4]
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 47:17:@104847.4]
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 47:17:@104848.4]
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 47:17:@104849.4]
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 47:17:@104850.4]
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 47:17:@104851.4]
  assign io_dram_wdata_bits_wdata_8 = wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 47:17:@104852.4]
  assign io_dram_wdata_bits_wdata_9 = wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 47:17:@104853.4]
  assign io_dram_wdata_bits_wdata_10 = wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 47:17:@104854.4]
  assign io_dram_wdata_bits_wdata_11 = wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 47:17:@104855.4]
  assign io_dram_wdata_bits_wdata_12 = wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 47:17:@104856.4]
  assign io_dram_wdata_bits_wdata_13 = wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 47:17:@104857.4]
  assign io_dram_wdata_bits_wdata_14 = wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 47:17:@104858.4]
  assign io_dram_wdata_bits_wdata_15 = wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 47:17:@104859.4]
  assign io_dram_wdata_bits_wdata_16 = wdataMux_io_out_bits_wdata_16; // @[StreamArbiter.scala 47:17:@104860.4]
  assign io_dram_wdata_bits_wdata_17 = wdataMux_io_out_bits_wdata_17; // @[StreamArbiter.scala 47:17:@104861.4]
  assign io_dram_wdata_bits_wdata_18 = wdataMux_io_out_bits_wdata_18; // @[StreamArbiter.scala 47:17:@104862.4]
  assign io_dram_wdata_bits_wdata_19 = wdataMux_io_out_bits_wdata_19; // @[StreamArbiter.scala 47:17:@104863.4]
  assign io_dram_wdata_bits_wdata_20 = wdataMux_io_out_bits_wdata_20; // @[StreamArbiter.scala 47:17:@104864.4]
  assign io_dram_wdata_bits_wdata_21 = wdataMux_io_out_bits_wdata_21; // @[StreamArbiter.scala 47:17:@104865.4]
  assign io_dram_wdata_bits_wdata_22 = wdataMux_io_out_bits_wdata_22; // @[StreamArbiter.scala 47:17:@104866.4]
  assign io_dram_wdata_bits_wdata_23 = wdataMux_io_out_bits_wdata_23; // @[StreamArbiter.scala 47:17:@104867.4]
  assign io_dram_wdata_bits_wdata_24 = wdataMux_io_out_bits_wdata_24; // @[StreamArbiter.scala 47:17:@104868.4]
  assign io_dram_wdata_bits_wdata_25 = wdataMux_io_out_bits_wdata_25; // @[StreamArbiter.scala 47:17:@104869.4]
  assign io_dram_wdata_bits_wdata_26 = wdataMux_io_out_bits_wdata_26; // @[StreamArbiter.scala 47:17:@104870.4]
  assign io_dram_wdata_bits_wdata_27 = wdataMux_io_out_bits_wdata_27; // @[StreamArbiter.scala 47:17:@104871.4]
  assign io_dram_wdata_bits_wdata_28 = wdataMux_io_out_bits_wdata_28; // @[StreamArbiter.scala 47:17:@104872.4]
  assign io_dram_wdata_bits_wdata_29 = wdataMux_io_out_bits_wdata_29; // @[StreamArbiter.scala 47:17:@104873.4]
  assign io_dram_wdata_bits_wdata_30 = wdataMux_io_out_bits_wdata_30; // @[StreamArbiter.scala 47:17:@104874.4]
  assign io_dram_wdata_bits_wdata_31 = wdataMux_io_out_bits_wdata_31; // @[StreamArbiter.scala 47:17:@104875.4]
  assign io_dram_wdata_bits_wdata_32 = wdataMux_io_out_bits_wdata_32; // @[StreamArbiter.scala 47:17:@104876.4]
  assign io_dram_wdata_bits_wdata_33 = wdataMux_io_out_bits_wdata_33; // @[StreamArbiter.scala 47:17:@104877.4]
  assign io_dram_wdata_bits_wdata_34 = wdataMux_io_out_bits_wdata_34; // @[StreamArbiter.scala 47:17:@104878.4]
  assign io_dram_wdata_bits_wdata_35 = wdataMux_io_out_bits_wdata_35; // @[StreamArbiter.scala 47:17:@104879.4]
  assign io_dram_wdata_bits_wdata_36 = wdataMux_io_out_bits_wdata_36; // @[StreamArbiter.scala 47:17:@104880.4]
  assign io_dram_wdata_bits_wdata_37 = wdataMux_io_out_bits_wdata_37; // @[StreamArbiter.scala 47:17:@104881.4]
  assign io_dram_wdata_bits_wdata_38 = wdataMux_io_out_bits_wdata_38; // @[StreamArbiter.scala 47:17:@104882.4]
  assign io_dram_wdata_bits_wdata_39 = wdataMux_io_out_bits_wdata_39; // @[StreamArbiter.scala 47:17:@104883.4]
  assign io_dram_wdata_bits_wdata_40 = wdataMux_io_out_bits_wdata_40; // @[StreamArbiter.scala 47:17:@104884.4]
  assign io_dram_wdata_bits_wdata_41 = wdataMux_io_out_bits_wdata_41; // @[StreamArbiter.scala 47:17:@104885.4]
  assign io_dram_wdata_bits_wdata_42 = wdataMux_io_out_bits_wdata_42; // @[StreamArbiter.scala 47:17:@104886.4]
  assign io_dram_wdata_bits_wdata_43 = wdataMux_io_out_bits_wdata_43; // @[StreamArbiter.scala 47:17:@104887.4]
  assign io_dram_wdata_bits_wdata_44 = wdataMux_io_out_bits_wdata_44; // @[StreamArbiter.scala 47:17:@104888.4]
  assign io_dram_wdata_bits_wdata_45 = wdataMux_io_out_bits_wdata_45; // @[StreamArbiter.scala 47:17:@104889.4]
  assign io_dram_wdata_bits_wdata_46 = wdataMux_io_out_bits_wdata_46; // @[StreamArbiter.scala 47:17:@104890.4]
  assign io_dram_wdata_bits_wdata_47 = wdataMux_io_out_bits_wdata_47; // @[StreamArbiter.scala 47:17:@104891.4]
  assign io_dram_wdata_bits_wdata_48 = wdataMux_io_out_bits_wdata_48; // @[StreamArbiter.scala 47:17:@104892.4]
  assign io_dram_wdata_bits_wdata_49 = wdataMux_io_out_bits_wdata_49; // @[StreamArbiter.scala 47:17:@104893.4]
  assign io_dram_wdata_bits_wdata_50 = wdataMux_io_out_bits_wdata_50; // @[StreamArbiter.scala 47:17:@104894.4]
  assign io_dram_wdata_bits_wdata_51 = wdataMux_io_out_bits_wdata_51; // @[StreamArbiter.scala 47:17:@104895.4]
  assign io_dram_wdata_bits_wdata_52 = wdataMux_io_out_bits_wdata_52; // @[StreamArbiter.scala 47:17:@104896.4]
  assign io_dram_wdata_bits_wdata_53 = wdataMux_io_out_bits_wdata_53; // @[StreamArbiter.scala 47:17:@104897.4]
  assign io_dram_wdata_bits_wdata_54 = wdataMux_io_out_bits_wdata_54; // @[StreamArbiter.scala 47:17:@104898.4]
  assign io_dram_wdata_bits_wdata_55 = wdataMux_io_out_bits_wdata_55; // @[StreamArbiter.scala 47:17:@104899.4]
  assign io_dram_wdata_bits_wdata_56 = wdataMux_io_out_bits_wdata_56; // @[StreamArbiter.scala 47:17:@104900.4]
  assign io_dram_wdata_bits_wdata_57 = wdataMux_io_out_bits_wdata_57; // @[StreamArbiter.scala 47:17:@104901.4]
  assign io_dram_wdata_bits_wdata_58 = wdataMux_io_out_bits_wdata_58; // @[StreamArbiter.scala 47:17:@104902.4]
  assign io_dram_wdata_bits_wdata_59 = wdataMux_io_out_bits_wdata_59; // @[StreamArbiter.scala 47:17:@104903.4]
  assign io_dram_wdata_bits_wdata_60 = wdataMux_io_out_bits_wdata_60; // @[StreamArbiter.scala 47:17:@104904.4]
  assign io_dram_wdata_bits_wdata_61 = wdataMux_io_out_bits_wdata_61; // @[StreamArbiter.scala 47:17:@104905.4]
  assign io_dram_wdata_bits_wdata_62 = wdataMux_io_out_bits_wdata_62; // @[StreamArbiter.scala 47:17:@104906.4]
  assign io_dram_wdata_bits_wdata_63 = wdataMux_io_out_bits_wdata_63; // @[StreamArbiter.scala 47:17:@104907.4]
  assign io_dram_wdata_bits_wstrb_0 = wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 47:17:@104780.4]
  assign io_dram_wdata_bits_wstrb_1 = wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 47:17:@104781.4]
  assign io_dram_wdata_bits_wstrb_2 = wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 47:17:@104782.4]
  assign io_dram_wdata_bits_wstrb_3 = wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 47:17:@104783.4]
  assign io_dram_wdata_bits_wstrb_4 = wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 47:17:@104784.4]
  assign io_dram_wdata_bits_wstrb_5 = wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 47:17:@104785.4]
  assign io_dram_wdata_bits_wstrb_6 = wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 47:17:@104786.4]
  assign io_dram_wdata_bits_wstrb_7 = wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 47:17:@104787.4]
  assign io_dram_wdata_bits_wstrb_8 = wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 47:17:@104788.4]
  assign io_dram_wdata_bits_wstrb_9 = wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 47:17:@104789.4]
  assign io_dram_wdata_bits_wstrb_10 = wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 47:17:@104790.4]
  assign io_dram_wdata_bits_wstrb_11 = wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 47:17:@104791.4]
  assign io_dram_wdata_bits_wstrb_12 = wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 47:17:@104792.4]
  assign io_dram_wdata_bits_wstrb_13 = wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 47:17:@104793.4]
  assign io_dram_wdata_bits_wstrb_14 = wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 47:17:@104794.4]
  assign io_dram_wdata_bits_wstrb_15 = wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 47:17:@104795.4]
  assign io_dram_wdata_bits_wstrb_16 = wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 47:17:@104796.4]
  assign io_dram_wdata_bits_wstrb_17 = wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 47:17:@104797.4]
  assign io_dram_wdata_bits_wstrb_18 = wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 47:17:@104798.4]
  assign io_dram_wdata_bits_wstrb_19 = wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 47:17:@104799.4]
  assign io_dram_wdata_bits_wstrb_20 = wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 47:17:@104800.4]
  assign io_dram_wdata_bits_wstrb_21 = wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 47:17:@104801.4]
  assign io_dram_wdata_bits_wstrb_22 = wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 47:17:@104802.4]
  assign io_dram_wdata_bits_wstrb_23 = wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 47:17:@104803.4]
  assign io_dram_wdata_bits_wstrb_24 = wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 47:17:@104804.4]
  assign io_dram_wdata_bits_wstrb_25 = wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 47:17:@104805.4]
  assign io_dram_wdata_bits_wstrb_26 = wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 47:17:@104806.4]
  assign io_dram_wdata_bits_wstrb_27 = wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 47:17:@104807.4]
  assign io_dram_wdata_bits_wstrb_28 = wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 47:17:@104808.4]
  assign io_dram_wdata_bits_wstrb_29 = wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 47:17:@104809.4]
  assign io_dram_wdata_bits_wstrb_30 = wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 47:17:@104810.4]
  assign io_dram_wdata_bits_wstrb_31 = wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 47:17:@104811.4]
  assign io_dram_wdata_bits_wstrb_32 = wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 47:17:@104812.4]
  assign io_dram_wdata_bits_wstrb_33 = wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 47:17:@104813.4]
  assign io_dram_wdata_bits_wstrb_34 = wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 47:17:@104814.4]
  assign io_dram_wdata_bits_wstrb_35 = wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 47:17:@104815.4]
  assign io_dram_wdata_bits_wstrb_36 = wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 47:17:@104816.4]
  assign io_dram_wdata_bits_wstrb_37 = wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 47:17:@104817.4]
  assign io_dram_wdata_bits_wstrb_38 = wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 47:17:@104818.4]
  assign io_dram_wdata_bits_wstrb_39 = wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 47:17:@104819.4]
  assign io_dram_wdata_bits_wstrb_40 = wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 47:17:@104820.4]
  assign io_dram_wdata_bits_wstrb_41 = wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 47:17:@104821.4]
  assign io_dram_wdata_bits_wstrb_42 = wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 47:17:@104822.4]
  assign io_dram_wdata_bits_wstrb_43 = wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 47:17:@104823.4]
  assign io_dram_wdata_bits_wstrb_44 = wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 47:17:@104824.4]
  assign io_dram_wdata_bits_wstrb_45 = wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 47:17:@104825.4]
  assign io_dram_wdata_bits_wstrb_46 = wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 47:17:@104826.4]
  assign io_dram_wdata_bits_wstrb_47 = wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 47:17:@104827.4]
  assign io_dram_wdata_bits_wstrb_48 = wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 47:17:@104828.4]
  assign io_dram_wdata_bits_wstrb_49 = wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 47:17:@104829.4]
  assign io_dram_wdata_bits_wstrb_50 = wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 47:17:@104830.4]
  assign io_dram_wdata_bits_wstrb_51 = wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 47:17:@104831.4]
  assign io_dram_wdata_bits_wstrb_52 = wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 47:17:@104832.4]
  assign io_dram_wdata_bits_wstrb_53 = wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 47:17:@104833.4]
  assign io_dram_wdata_bits_wstrb_54 = wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 47:17:@104834.4]
  assign io_dram_wdata_bits_wstrb_55 = wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 47:17:@104835.4]
  assign io_dram_wdata_bits_wstrb_56 = wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 47:17:@104836.4]
  assign io_dram_wdata_bits_wstrb_57 = wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 47:17:@104837.4]
  assign io_dram_wdata_bits_wstrb_58 = wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 47:17:@104838.4]
  assign io_dram_wdata_bits_wstrb_59 = wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 47:17:@104839.4]
  assign io_dram_wdata_bits_wstrb_60 = wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 47:17:@104840.4]
  assign io_dram_wdata_bits_wstrb_61 = wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 47:17:@104841.4]
  assign io_dram_wdata_bits_wstrb_62 = wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 47:17:@104842.4]
  assign io_dram_wdata_bits_wstrb_63 = wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 47:17:@104843.4]
  assign io_dram_rresp_ready = _T_510 ? 1'h0 : io_app_0_rresp_ready; // @[StreamArbiter.scala 72:23:@105100.4]
  assign io_dram_wresp_ready = _T_520 ? io_app_1_wresp_ready : 1'h0; // @[StreamArbiter.scala 73:23:@105105.4]
  assign RetimeWrapper_clock = clock; // @[:@104428.4]
  assign RetimeWrapper_reset = reset; // @[:@104429.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@104431.4]
  assign RetimeWrapper_io_in = _GEN_1 ? _T_412 : priorityActive; // @[package.scala 94:16:@104430.4]
  assign RetimeWrapper_1_clock = clock; // @[:@104435.4]
  assign RetimeWrapper_1_reset = reset; // @[:@104436.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@104438.4]
  assign RetimeWrapper_1_io_in = _GEN_1 ? _T_412 : priorityActive; // @[package.scala 94:16:@104437.4]
  assign cmdMux_io_in_valid = io_app_0_cmd_valid | io_app_1_cmd_valid; // @[StreamArbiter.scala 26:22:@104448.4]
  assign cmdMux_io_in_bits_0_addr = io_app_0_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@104454.4]
  assign cmdMux_io_in_bits_0_size = io_app_0_cmd_bits_size; // @[StreamArbiter.scala 29:9:@104453.4]
  assign cmdMux_io_in_bits_1_addr = io_app_1_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@104472.4]
  assign cmdMux_io_in_bits_1_size = io_app_1_cmd_bits_size; // @[StreamArbiter.scala 29:9:@104471.4]
  assign cmdMux_io_sel = _GEN_1 ? _T_412 : priorityActive; // @[StreamArbiter.scala 27:17:@104449.4]
  assign cmdMux_io_out_ready = io_dram_cmd_valid & io_dram_cmd_ready; // @[StreamArbiter.scala 46:15:@104778.4 StreamArbiter.scala 57:23:@104932.4]
  assign wdataMux_io_in_valid = _T_458 & _T_459; // @[StreamArbiter.scala 42:24:@104512.4]
  assign wdataMux_io_in_bits_1_wdata_0 = io_app_1_wdata_bits_wdata_0; // @[StreamArbiter.scala 44:23:@104708.4]
  assign wdataMux_io_in_bits_1_wdata_1 = io_app_1_wdata_bits_wdata_1; // @[StreamArbiter.scala 44:23:@104709.4]
  assign wdataMux_io_in_bits_1_wdata_2 = io_app_1_wdata_bits_wdata_2; // @[StreamArbiter.scala 44:23:@104710.4]
  assign wdataMux_io_in_bits_1_wdata_3 = io_app_1_wdata_bits_wdata_3; // @[StreamArbiter.scala 44:23:@104711.4]
  assign wdataMux_io_in_bits_1_wdata_4 = io_app_1_wdata_bits_wdata_4; // @[StreamArbiter.scala 44:23:@104712.4]
  assign wdataMux_io_in_bits_1_wdata_5 = io_app_1_wdata_bits_wdata_5; // @[StreamArbiter.scala 44:23:@104713.4]
  assign wdataMux_io_in_bits_1_wdata_6 = io_app_1_wdata_bits_wdata_6; // @[StreamArbiter.scala 44:23:@104714.4]
  assign wdataMux_io_in_bits_1_wdata_7 = io_app_1_wdata_bits_wdata_7; // @[StreamArbiter.scala 44:23:@104715.4]
  assign wdataMux_io_in_bits_1_wdata_8 = io_app_1_wdata_bits_wdata_8; // @[StreamArbiter.scala 44:23:@104716.4]
  assign wdataMux_io_in_bits_1_wdata_9 = io_app_1_wdata_bits_wdata_9; // @[StreamArbiter.scala 44:23:@104717.4]
  assign wdataMux_io_in_bits_1_wdata_10 = io_app_1_wdata_bits_wdata_10; // @[StreamArbiter.scala 44:23:@104718.4]
  assign wdataMux_io_in_bits_1_wdata_11 = io_app_1_wdata_bits_wdata_11; // @[StreamArbiter.scala 44:23:@104719.4]
  assign wdataMux_io_in_bits_1_wdata_12 = io_app_1_wdata_bits_wdata_12; // @[StreamArbiter.scala 44:23:@104720.4]
  assign wdataMux_io_in_bits_1_wdata_13 = io_app_1_wdata_bits_wdata_13; // @[StreamArbiter.scala 44:23:@104721.4]
  assign wdataMux_io_in_bits_1_wdata_14 = io_app_1_wdata_bits_wdata_14; // @[StreamArbiter.scala 44:23:@104722.4]
  assign wdataMux_io_in_bits_1_wdata_15 = io_app_1_wdata_bits_wdata_15; // @[StreamArbiter.scala 44:23:@104723.4]
  assign wdataMux_io_in_bits_1_wdata_16 = io_app_1_wdata_bits_wdata_16; // @[StreamArbiter.scala 44:23:@104724.4]
  assign wdataMux_io_in_bits_1_wdata_17 = io_app_1_wdata_bits_wdata_17; // @[StreamArbiter.scala 44:23:@104725.4]
  assign wdataMux_io_in_bits_1_wdata_18 = io_app_1_wdata_bits_wdata_18; // @[StreamArbiter.scala 44:23:@104726.4]
  assign wdataMux_io_in_bits_1_wdata_19 = io_app_1_wdata_bits_wdata_19; // @[StreamArbiter.scala 44:23:@104727.4]
  assign wdataMux_io_in_bits_1_wdata_20 = io_app_1_wdata_bits_wdata_20; // @[StreamArbiter.scala 44:23:@104728.4]
  assign wdataMux_io_in_bits_1_wdata_21 = io_app_1_wdata_bits_wdata_21; // @[StreamArbiter.scala 44:23:@104729.4]
  assign wdataMux_io_in_bits_1_wdata_22 = io_app_1_wdata_bits_wdata_22; // @[StreamArbiter.scala 44:23:@104730.4]
  assign wdataMux_io_in_bits_1_wdata_23 = io_app_1_wdata_bits_wdata_23; // @[StreamArbiter.scala 44:23:@104731.4]
  assign wdataMux_io_in_bits_1_wdata_24 = io_app_1_wdata_bits_wdata_24; // @[StreamArbiter.scala 44:23:@104732.4]
  assign wdataMux_io_in_bits_1_wdata_25 = io_app_1_wdata_bits_wdata_25; // @[StreamArbiter.scala 44:23:@104733.4]
  assign wdataMux_io_in_bits_1_wdata_26 = io_app_1_wdata_bits_wdata_26; // @[StreamArbiter.scala 44:23:@104734.4]
  assign wdataMux_io_in_bits_1_wdata_27 = io_app_1_wdata_bits_wdata_27; // @[StreamArbiter.scala 44:23:@104735.4]
  assign wdataMux_io_in_bits_1_wdata_28 = io_app_1_wdata_bits_wdata_28; // @[StreamArbiter.scala 44:23:@104736.4]
  assign wdataMux_io_in_bits_1_wdata_29 = io_app_1_wdata_bits_wdata_29; // @[StreamArbiter.scala 44:23:@104737.4]
  assign wdataMux_io_in_bits_1_wdata_30 = io_app_1_wdata_bits_wdata_30; // @[StreamArbiter.scala 44:23:@104738.4]
  assign wdataMux_io_in_bits_1_wdata_31 = io_app_1_wdata_bits_wdata_31; // @[StreamArbiter.scala 44:23:@104739.4]
  assign wdataMux_io_in_bits_1_wdata_32 = io_app_1_wdata_bits_wdata_32; // @[StreamArbiter.scala 44:23:@104740.4]
  assign wdataMux_io_in_bits_1_wdata_33 = io_app_1_wdata_bits_wdata_33; // @[StreamArbiter.scala 44:23:@104741.4]
  assign wdataMux_io_in_bits_1_wdata_34 = io_app_1_wdata_bits_wdata_34; // @[StreamArbiter.scala 44:23:@104742.4]
  assign wdataMux_io_in_bits_1_wdata_35 = io_app_1_wdata_bits_wdata_35; // @[StreamArbiter.scala 44:23:@104743.4]
  assign wdataMux_io_in_bits_1_wdata_36 = io_app_1_wdata_bits_wdata_36; // @[StreamArbiter.scala 44:23:@104744.4]
  assign wdataMux_io_in_bits_1_wdata_37 = io_app_1_wdata_bits_wdata_37; // @[StreamArbiter.scala 44:23:@104745.4]
  assign wdataMux_io_in_bits_1_wdata_38 = io_app_1_wdata_bits_wdata_38; // @[StreamArbiter.scala 44:23:@104746.4]
  assign wdataMux_io_in_bits_1_wdata_39 = io_app_1_wdata_bits_wdata_39; // @[StreamArbiter.scala 44:23:@104747.4]
  assign wdataMux_io_in_bits_1_wdata_40 = io_app_1_wdata_bits_wdata_40; // @[StreamArbiter.scala 44:23:@104748.4]
  assign wdataMux_io_in_bits_1_wdata_41 = io_app_1_wdata_bits_wdata_41; // @[StreamArbiter.scala 44:23:@104749.4]
  assign wdataMux_io_in_bits_1_wdata_42 = io_app_1_wdata_bits_wdata_42; // @[StreamArbiter.scala 44:23:@104750.4]
  assign wdataMux_io_in_bits_1_wdata_43 = io_app_1_wdata_bits_wdata_43; // @[StreamArbiter.scala 44:23:@104751.4]
  assign wdataMux_io_in_bits_1_wdata_44 = io_app_1_wdata_bits_wdata_44; // @[StreamArbiter.scala 44:23:@104752.4]
  assign wdataMux_io_in_bits_1_wdata_45 = io_app_1_wdata_bits_wdata_45; // @[StreamArbiter.scala 44:23:@104753.4]
  assign wdataMux_io_in_bits_1_wdata_46 = io_app_1_wdata_bits_wdata_46; // @[StreamArbiter.scala 44:23:@104754.4]
  assign wdataMux_io_in_bits_1_wdata_47 = io_app_1_wdata_bits_wdata_47; // @[StreamArbiter.scala 44:23:@104755.4]
  assign wdataMux_io_in_bits_1_wdata_48 = io_app_1_wdata_bits_wdata_48; // @[StreamArbiter.scala 44:23:@104756.4]
  assign wdataMux_io_in_bits_1_wdata_49 = io_app_1_wdata_bits_wdata_49; // @[StreamArbiter.scala 44:23:@104757.4]
  assign wdataMux_io_in_bits_1_wdata_50 = io_app_1_wdata_bits_wdata_50; // @[StreamArbiter.scala 44:23:@104758.4]
  assign wdataMux_io_in_bits_1_wdata_51 = io_app_1_wdata_bits_wdata_51; // @[StreamArbiter.scala 44:23:@104759.4]
  assign wdataMux_io_in_bits_1_wdata_52 = io_app_1_wdata_bits_wdata_52; // @[StreamArbiter.scala 44:23:@104760.4]
  assign wdataMux_io_in_bits_1_wdata_53 = io_app_1_wdata_bits_wdata_53; // @[StreamArbiter.scala 44:23:@104761.4]
  assign wdataMux_io_in_bits_1_wdata_54 = io_app_1_wdata_bits_wdata_54; // @[StreamArbiter.scala 44:23:@104762.4]
  assign wdataMux_io_in_bits_1_wdata_55 = io_app_1_wdata_bits_wdata_55; // @[StreamArbiter.scala 44:23:@104763.4]
  assign wdataMux_io_in_bits_1_wdata_56 = io_app_1_wdata_bits_wdata_56; // @[StreamArbiter.scala 44:23:@104764.4]
  assign wdataMux_io_in_bits_1_wdata_57 = io_app_1_wdata_bits_wdata_57; // @[StreamArbiter.scala 44:23:@104765.4]
  assign wdataMux_io_in_bits_1_wdata_58 = io_app_1_wdata_bits_wdata_58; // @[StreamArbiter.scala 44:23:@104766.4]
  assign wdataMux_io_in_bits_1_wdata_59 = io_app_1_wdata_bits_wdata_59; // @[StreamArbiter.scala 44:23:@104767.4]
  assign wdataMux_io_in_bits_1_wdata_60 = io_app_1_wdata_bits_wdata_60; // @[StreamArbiter.scala 44:23:@104768.4]
  assign wdataMux_io_in_bits_1_wdata_61 = io_app_1_wdata_bits_wdata_61; // @[StreamArbiter.scala 44:23:@104769.4]
  assign wdataMux_io_in_bits_1_wdata_62 = io_app_1_wdata_bits_wdata_62; // @[StreamArbiter.scala 44:23:@104770.4]
  assign wdataMux_io_in_bits_1_wdata_63 = io_app_1_wdata_bits_wdata_63; // @[StreamArbiter.scala 44:23:@104771.4]
  assign wdataMux_io_in_bits_1_wstrb_0 = io_app_1_wdata_bits_wstrb_0; // @[StreamArbiter.scala 44:23:@104644.4]
  assign wdataMux_io_in_bits_1_wstrb_1 = io_app_1_wdata_bits_wstrb_1; // @[StreamArbiter.scala 44:23:@104645.4]
  assign wdataMux_io_in_bits_1_wstrb_2 = io_app_1_wdata_bits_wstrb_2; // @[StreamArbiter.scala 44:23:@104646.4]
  assign wdataMux_io_in_bits_1_wstrb_3 = io_app_1_wdata_bits_wstrb_3; // @[StreamArbiter.scala 44:23:@104647.4]
  assign wdataMux_io_in_bits_1_wstrb_4 = io_app_1_wdata_bits_wstrb_4; // @[StreamArbiter.scala 44:23:@104648.4]
  assign wdataMux_io_in_bits_1_wstrb_5 = io_app_1_wdata_bits_wstrb_5; // @[StreamArbiter.scala 44:23:@104649.4]
  assign wdataMux_io_in_bits_1_wstrb_6 = io_app_1_wdata_bits_wstrb_6; // @[StreamArbiter.scala 44:23:@104650.4]
  assign wdataMux_io_in_bits_1_wstrb_7 = io_app_1_wdata_bits_wstrb_7; // @[StreamArbiter.scala 44:23:@104651.4]
  assign wdataMux_io_in_bits_1_wstrb_8 = io_app_1_wdata_bits_wstrb_8; // @[StreamArbiter.scala 44:23:@104652.4]
  assign wdataMux_io_in_bits_1_wstrb_9 = io_app_1_wdata_bits_wstrb_9; // @[StreamArbiter.scala 44:23:@104653.4]
  assign wdataMux_io_in_bits_1_wstrb_10 = io_app_1_wdata_bits_wstrb_10; // @[StreamArbiter.scala 44:23:@104654.4]
  assign wdataMux_io_in_bits_1_wstrb_11 = io_app_1_wdata_bits_wstrb_11; // @[StreamArbiter.scala 44:23:@104655.4]
  assign wdataMux_io_in_bits_1_wstrb_12 = io_app_1_wdata_bits_wstrb_12; // @[StreamArbiter.scala 44:23:@104656.4]
  assign wdataMux_io_in_bits_1_wstrb_13 = io_app_1_wdata_bits_wstrb_13; // @[StreamArbiter.scala 44:23:@104657.4]
  assign wdataMux_io_in_bits_1_wstrb_14 = io_app_1_wdata_bits_wstrb_14; // @[StreamArbiter.scala 44:23:@104658.4]
  assign wdataMux_io_in_bits_1_wstrb_15 = io_app_1_wdata_bits_wstrb_15; // @[StreamArbiter.scala 44:23:@104659.4]
  assign wdataMux_io_in_bits_1_wstrb_16 = io_app_1_wdata_bits_wstrb_16; // @[StreamArbiter.scala 44:23:@104660.4]
  assign wdataMux_io_in_bits_1_wstrb_17 = io_app_1_wdata_bits_wstrb_17; // @[StreamArbiter.scala 44:23:@104661.4]
  assign wdataMux_io_in_bits_1_wstrb_18 = io_app_1_wdata_bits_wstrb_18; // @[StreamArbiter.scala 44:23:@104662.4]
  assign wdataMux_io_in_bits_1_wstrb_19 = io_app_1_wdata_bits_wstrb_19; // @[StreamArbiter.scala 44:23:@104663.4]
  assign wdataMux_io_in_bits_1_wstrb_20 = io_app_1_wdata_bits_wstrb_20; // @[StreamArbiter.scala 44:23:@104664.4]
  assign wdataMux_io_in_bits_1_wstrb_21 = io_app_1_wdata_bits_wstrb_21; // @[StreamArbiter.scala 44:23:@104665.4]
  assign wdataMux_io_in_bits_1_wstrb_22 = io_app_1_wdata_bits_wstrb_22; // @[StreamArbiter.scala 44:23:@104666.4]
  assign wdataMux_io_in_bits_1_wstrb_23 = io_app_1_wdata_bits_wstrb_23; // @[StreamArbiter.scala 44:23:@104667.4]
  assign wdataMux_io_in_bits_1_wstrb_24 = io_app_1_wdata_bits_wstrb_24; // @[StreamArbiter.scala 44:23:@104668.4]
  assign wdataMux_io_in_bits_1_wstrb_25 = io_app_1_wdata_bits_wstrb_25; // @[StreamArbiter.scala 44:23:@104669.4]
  assign wdataMux_io_in_bits_1_wstrb_26 = io_app_1_wdata_bits_wstrb_26; // @[StreamArbiter.scala 44:23:@104670.4]
  assign wdataMux_io_in_bits_1_wstrb_27 = io_app_1_wdata_bits_wstrb_27; // @[StreamArbiter.scala 44:23:@104671.4]
  assign wdataMux_io_in_bits_1_wstrb_28 = io_app_1_wdata_bits_wstrb_28; // @[StreamArbiter.scala 44:23:@104672.4]
  assign wdataMux_io_in_bits_1_wstrb_29 = io_app_1_wdata_bits_wstrb_29; // @[StreamArbiter.scala 44:23:@104673.4]
  assign wdataMux_io_in_bits_1_wstrb_30 = io_app_1_wdata_bits_wstrb_30; // @[StreamArbiter.scala 44:23:@104674.4]
  assign wdataMux_io_in_bits_1_wstrb_31 = io_app_1_wdata_bits_wstrb_31; // @[StreamArbiter.scala 44:23:@104675.4]
  assign wdataMux_io_in_bits_1_wstrb_32 = io_app_1_wdata_bits_wstrb_32; // @[StreamArbiter.scala 44:23:@104676.4]
  assign wdataMux_io_in_bits_1_wstrb_33 = io_app_1_wdata_bits_wstrb_33; // @[StreamArbiter.scala 44:23:@104677.4]
  assign wdataMux_io_in_bits_1_wstrb_34 = io_app_1_wdata_bits_wstrb_34; // @[StreamArbiter.scala 44:23:@104678.4]
  assign wdataMux_io_in_bits_1_wstrb_35 = io_app_1_wdata_bits_wstrb_35; // @[StreamArbiter.scala 44:23:@104679.4]
  assign wdataMux_io_in_bits_1_wstrb_36 = io_app_1_wdata_bits_wstrb_36; // @[StreamArbiter.scala 44:23:@104680.4]
  assign wdataMux_io_in_bits_1_wstrb_37 = io_app_1_wdata_bits_wstrb_37; // @[StreamArbiter.scala 44:23:@104681.4]
  assign wdataMux_io_in_bits_1_wstrb_38 = io_app_1_wdata_bits_wstrb_38; // @[StreamArbiter.scala 44:23:@104682.4]
  assign wdataMux_io_in_bits_1_wstrb_39 = io_app_1_wdata_bits_wstrb_39; // @[StreamArbiter.scala 44:23:@104683.4]
  assign wdataMux_io_in_bits_1_wstrb_40 = io_app_1_wdata_bits_wstrb_40; // @[StreamArbiter.scala 44:23:@104684.4]
  assign wdataMux_io_in_bits_1_wstrb_41 = io_app_1_wdata_bits_wstrb_41; // @[StreamArbiter.scala 44:23:@104685.4]
  assign wdataMux_io_in_bits_1_wstrb_42 = io_app_1_wdata_bits_wstrb_42; // @[StreamArbiter.scala 44:23:@104686.4]
  assign wdataMux_io_in_bits_1_wstrb_43 = io_app_1_wdata_bits_wstrb_43; // @[StreamArbiter.scala 44:23:@104687.4]
  assign wdataMux_io_in_bits_1_wstrb_44 = io_app_1_wdata_bits_wstrb_44; // @[StreamArbiter.scala 44:23:@104688.4]
  assign wdataMux_io_in_bits_1_wstrb_45 = io_app_1_wdata_bits_wstrb_45; // @[StreamArbiter.scala 44:23:@104689.4]
  assign wdataMux_io_in_bits_1_wstrb_46 = io_app_1_wdata_bits_wstrb_46; // @[StreamArbiter.scala 44:23:@104690.4]
  assign wdataMux_io_in_bits_1_wstrb_47 = io_app_1_wdata_bits_wstrb_47; // @[StreamArbiter.scala 44:23:@104691.4]
  assign wdataMux_io_in_bits_1_wstrb_48 = io_app_1_wdata_bits_wstrb_48; // @[StreamArbiter.scala 44:23:@104692.4]
  assign wdataMux_io_in_bits_1_wstrb_49 = io_app_1_wdata_bits_wstrb_49; // @[StreamArbiter.scala 44:23:@104693.4]
  assign wdataMux_io_in_bits_1_wstrb_50 = io_app_1_wdata_bits_wstrb_50; // @[StreamArbiter.scala 44:23:@104694.4]
  assign wdataMux_io_in_bits_1_wstrb_51 = io_app_1_wdata_bits_wstrb_51; // @[StreamArbiter.scala 44:23:@104695.4]
  assign wdataMux_io_in_bits_1_wstrb_52 = io_app_1_wdata_bits_wstrb_52; // @[StreamArbiter.scala 44:23:@104696.4]
  assign wdataMux_io_in_bits_1_wstrb_53 = io_app_1_wdata_bits_wstrb_53; // @[StreamArbiter.scala 44:23:@104697.4]
  assign wdataMux_io_in_bits_1_wstrb_54 = io_app_1_wdata_bits_wstrb_54; // @[StreamArbiter.scala 44:23:@104698.4]
  assign wdataMux_io_in_bits_1_wstrb_55 = io_app_1_wdata_bits_wstrb_55; // @[StreamArbiter.scala 44:23:@104699.4]
  assign wdataMux_io_in_bits_1_wstrb_56 = io_app_1_wdata_bits_wstrb_56; // @[StreamArbiter.scala 44:23:@104700.4]
  assign wdataMux_io_in_bits_1_wstrb_57 = io_app_1_wdata_bits_wstrb_57; // @[StreamArbiter.scala 44:23:@104701.4]
  assign wdataMux_io_in_bits_1_wstrb_58 = io_app_1_wdata_bits_wstrb_58; // @[StreamArbiter.scala 44:23:@104702.4]
  assign wdataMux_io_in_bits_1_wstrb_59 = io_app_1_wdata_bits_wstrb_59; // @[StreamArbiter.scala 44:23:@104703.4]
  assign wdataMux_io_in_bits_1_wstrb_60 = io_app_1_wdata_bits_wstrb_60; // @[StreamArbiter.scala 44:23:@104704.4]
  assign wdataMux_io_in_bits_1_wstrb_61 = io_app_1_wdata_bits_wstrb_61; // @[StreamArbiter.scala 44:23:@104705.4]
  assign wdataMux_io_in_bits_1_wstrb_62 = io_app_1_wdata_bits_wstrb_62; // @[StreamArbiter.scala 44:23:@104706.4]
  assign wdataMux_io_in_bits_1_wstrb_63 = io_app_1_wdata_bits_wstrb_63; // @[StreamArbiter.scala 44:23:@104707.4]
  assign wdataMux_io_sel = _T_444[0]; // @[StreamArbiter.scala 43:19:@104513.4]
  assign wdataMux_io_out_ready = io_dram_wdata_valid & io_dram_wdata_ready; // @[StreamArbiter.scala 47:17:@104909.4 StreamArbiter.scala 58:25:@104933.4]
  assign elementCtr_clock = clock; // @[:@104490.4]
  assign elementCtr_reset = reset; // @[:@104491.4]
  assign elementCtr_io_reset = cmdMux_io_out_ready; // @[StreamArbiter.scala 38:23:@104494.4]
  assign elementCtr_io_enable = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:24:@104493.4]
endmodule
module Counter_112( // @[:@105107.2]
  input         clock, // @[:@105108.4]
  input         reset, // @[:@105109.4]
  input         io_reset, // @[:@105110.4]
  input         io_enable, // @[:@105110.4]
  input  [31:0] io_stride, // @[:@105110.4]
  output [31:0] io_out, // @[:@105110.4]
  output [31:0] io_next // @[:@105110.4]
);
  reg [31:0] count; // @[Counter.scala 15:22:@105112.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_17; // @[Counter.scala 17:24:@105113.4]
  wire [31:0] newCount; // @[Counter.scala 17:24:@105114.4]
  wire [31:0] _GEN_0; // @[Counter.scala 21:26:@105119.6]
  wire [31:0] _GEN_1; // @[Counter.scala 19:18:@105115.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@105113.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@105114.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@105119.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 19:18:@105115.4]
  assign io_out = count; // @[Counter.scala 25:10:@105122.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@105123.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module AXICmdSplit( // @[:@105125.2]
  input         clock, // @[:@105126.4]
  input         reset, // @[:@105127.4]
  output        io_in_cmd_ready, // @[:@105128.4]
  input         io_in_cmd_valid, // @[:@105128.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@105128.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@105128.4]
  input         io_in_cmd_bits_isWr, // @[:@105128.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@105128.4]
  output        io_in_wdata_ready, // @[:@105128.4]
  input         io_in_wdata_valid, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_0, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_1, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_2, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_3, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_4, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_5, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_6, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_7, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_8, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_9, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_10, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_11, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_12, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_13, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_14, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_15, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_16, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_17, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_18, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_19, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_20, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_21, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_22, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_23, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_24, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_25, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_26, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_27, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_28, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_29, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_30, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_31, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_32, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_33, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_34, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_35, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_36, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_37, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_38, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_39, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_40, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_41, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_42, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_43, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_44, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_45, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_46, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_47, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_48, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_49, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_50, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_51, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_52, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_53, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_54, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_55, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_56, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_57, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_58, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_59, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_60, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_61, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_62, // @[:@105128.4]
  input  [7:0]  io_in_wdata_bits_wdata_63, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@105128.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@105128.4]
  input         io_in_rresp_ready, // @[:@105128.4]
  output        io_in_rresp_valid, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_0, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_1, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_2, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_3, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_4, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_5, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_6, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_7, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_8, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_9, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_10, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_11, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_12, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_13, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_14, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_15, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_16, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_17, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_18, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_19, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_20, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_21, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_22, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_23, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_24, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_25, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_26, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_27, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_28, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_29, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_30, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_31, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_32, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_33, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_34, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_35, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_36, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_37, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_38, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_39, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_40, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_41, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_42, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_43, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_44, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_45, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_46, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_47, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_48, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_49, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_50, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_51, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_52, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_53, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_54, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_55, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_56, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_57, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_58, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_59, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_60, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_61, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_62, // @[:@105128.4]
  output [7:0]  io_in_rresp_bits_rdata_63, // @[:@105128.4]
  output [31:0] io_in_rresp_bits_tag, // @[:@105128.4]
  input         io_in_wresp_ready, // @[:@105128.4]
  output        io_in_wresp_valid, // @[:@105128.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@105128.4]
  input         io_out_cmd_ready, // @[:@105128.4]
  output        io_out_cmd_valid, // @[:@105128.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@105128.4]
  output [31:0] io_out_cmd_bits_size, // @[:@105128.4]
  output [63:0] io_out_cmd_bits_rawAddr, // @[:@105128.4]
  output        io_out_cmd_bits_isWr, // @[:@105128.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@105128.4]
  input         io_out_wdata_ready, // @[:@105128.4]
  output        io_out_wdata_valid, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_0, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_1, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_2, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_3, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_4, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_5, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_6, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_7, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_8, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_9, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_10, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_11, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_12, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_13, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_14, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_15, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_16, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_17, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_18, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_19, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_20, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_21, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_22, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_23, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_24, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_25, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_26, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_27, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_28, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_29, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_30, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_31, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_32, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_33, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_34, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_35, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_36, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_37, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_38, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_39, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_40, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_41, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_42, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_43, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_44, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_45, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_46, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_47, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_48, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_49, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_50, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_51, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_52, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_53, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_54, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_55, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_56, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_57, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_58, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_59, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_60, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_61, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_62, // @[:@105128.4]
  output [7:0]  io_out_wdata_bits_wdata_63, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@105128.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@105128.4]
  output        io_out_rresp_ready, // @[:@105128.4]
  input         io_out_rresp_valid, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_0, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_1, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_2, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_3, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_4, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_5, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_6, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_7, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_8, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_9, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_10, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_11, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_12, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_13, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_14, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_15, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_16, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_17, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_18, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_19, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_20, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_21, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_22, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_23, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_24, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_25, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_26, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_27, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_28, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_29, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_30, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_31, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_32, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_33, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_34, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_35, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_36, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_37, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_38, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_39, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_40, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_41, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_42, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_43, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_44, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_45, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_46, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_47, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_48, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_49, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_50, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_51, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_52, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_53, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_54, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_55, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_56, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_57, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_58, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_59, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_60, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_61, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_62, // @[:@105128.4]
  input  [7:0]  io_out_rresp_bits_rdata_63, // @[:@105128.4]
  input  [31:0] io_out_rresp_bits_tag, // @[:@105128.4]
  output        io_out_wresp_ready, // @[:@105128.4]
  input         io_out_wresp_valid, // @[:@105128.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@105128.4]
);
  wire  cmdSizeCounter_clock; // @[AXIProtocol.scala 18:30:@105338.4]
  wire  cmdSizeCounter_reset; // @[AXIProtocol.scala 18:30:@105338.4]
  wire  cmdSizeCounter_io_reset; // @[AXIProtocol.scala 18:30:@105338.4]
  wire  cmdSizeCounter_io_enable; // @[AXIProtocol.scala 18:30:@105338.4]
  wire [31:0] cmdSizeCounter_io_stride; // @[AXIProtocol.scala 18:30:@105338.4]
  wire [31:0] cmdSizeCounter_io_out; // @[AXIProtocol.scala 18:30:@105338.4]
  wire [31:0] cmdSizeCounter_io_next; // @[AXIProtocol.scala 18:30:@105338.4]
  wire [32:0] _T_199; // @[AXIProtocol.scala 20:46:@105341.4]
  wire [32:0] _T_200; // @[AXIProtocol.scala 20:46:@105342.4]
  wire [31:0] cmdSizeRemaining; // @[AXIProtocol.scala 20:46:@105343.4]
  wire  lastCmd; // @[AXIProtocol.scala 23:35:@105344.4]
  wire [37:0] _GEN_0; // @[AXIProtocol.scala 27:47:@105347.4]
  wire [37:0] addrOffsetBytes; // @[AXIProtocol.scala 27:47:@105347.4]
  wire [63:0] _GEN_1; // @[AXIProtocol.scala 28:49:@105348.4]
  wire [64:0] _T_201; // @[AXIProtocol.scala 28:49:@105348.4]
  wire [63:0] cmdAddr_bits; // @[AXIProtocol.scala 28:49:@105349.4]
  wire [57:0] _T_204; // @[FringeBundles.scala 158:22:@105352.4]
  wire [7:0] cmdTag_streamID; // @[FringeBundles.scala 114:28:@105359.4]
  wire [22:0] cmdTag_uid; // @[FringeBundles.scala 114:28:@105363.4]
  wire [23:0] _T_214; // @[FringeBundles.scala 115:37:@105366.4]
  wire  cmdIssue; // @[AXIProtocol.scala 36:35:@105369.4]
  wire  _T_223; // @[FringeBundles.scala 140:28:@105380.4]
  Counter_112 cmdSizeCounter ( // @[AXIProtocol.scala 18:30:@105338.4]
    .clock(cmdSizeCounter_clock),
    .reset(cmdSizeCounter_reset),
    .io_reset(cmdSizeCounter_io_reset),
    .io_enable(cmdSizeCounter_io_enable),
    .io_stride(cmdSizeCounter_io_stride),
    .io_out(cmdSizeCounter_io_out),
    .io_next(cmdSizeCounter_io_next)
  );
  assign _T_199 = io_in_cmd_bits_size - cmdSizeCounter_io_out; // @[AXIProtocol.scala 20:46:@105341.4]
  assign _T_200 = $unsigned(_T_199); // @[AXIProtocol.scala 20:46:@105342.4]
  assign cmdSizeRemaining = _T_200[31:0]; // @[AXIProtocol.scala 20:46:@105343.4]
  assign lastCmd = cmdSizeRemaining <= 32'h100; // @[AXIProtocol.scala 23:35:@105344.4]
  assign _GEN_0 = {{6'd0}, cmdSizeCounter_io_out}; // @[AXIProtocol.scala 27:47:@105347.4]
  assign addrOffsetBytes = _GEN_0 << 6; // @[AXIProtocol.scala 27:47:@105347.4]
  assign _GEN_1 = {{26'd0}, addrOffsetBytes}; // @[AXIProtocol.scala 28:49:@105348.4]
  assign _T_201 = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@105348.4]
  assign cmdAddr_bits = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@105349.4]
  assign _T_204 = cmdAddr_bits[63:6]; // @[FringeBundles.scala 158:22:@105352.4]
  assign cmdTag_streamID = io_in_cmd_bits_tag[7:0]; // @[FringeBundles.scala 114:28:@105359.4]
  assign cmdTag_uid = io_in_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@105363.4]
  assign _T_214 = {cmdTag_uid,lastCmd}; // @[FringeBundles.scala 115:37:@105366.4]
  assign cmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 36:35:@105369.4]
  assign _T_223 = io_out_wresp_bits_tag[8]; // @[FringeBundles.scala 140:28:@105380.4]
  assign io_in_cmd_ready = lastCmd & cmdIssue; // @[AXIProtocol.scala 15:10:@105337.4 AXIProtocol.scala 38:19:@105371.4]
  assign io_in_wdata_ready = io_out_wdata_ready; // @[AXIProtocol.scala 15:10:@105330.4]
  assign io_in_rresp_valid = io_out_rresp_valid; // @[AXIProtocol.scala 15:10:@105198.4]
  assign io_in_rresp_bits_rdata_0 = io_out_rresp_bits_rdata_0; // @[AXIProtocol.scala 15:10:@105134.4]
  assign io_in_rresp_bits_rdata_1 = io_out_rresp_bits_rdata_1; // @[AXIProtocol.scala 15:10:@105135.4]
  assign io_in_rresp_bits_rdata_2 = io_out_rresp_bits_rdata_2; // @[AXIProtocol.scala 15:10:@105136.4]
  assign io_in_rresp_bits_rdata_3 = io_out_rresp_bits_rdata_3; // @[AXIProtocol.scala 15:10:@105137.4]
  assign io_in_rresp_bits_rdata_4 = io_out_rresp_bits_rdata_4; // @[AXIProtocol.scala 15:10:@105138.4]
  assign io_in_rresp_bits_rdata_5 = io_out_rresp_bits_rdata_5; // @[AXIProtocol.scala 15:10:@105139.4]
  assign io_in_rresp_bits_rdata_6 = io_out_rresp_bits_rdata_6; // @[AXIProtocol.scala 15:10:@105140.4]
  assign io_in_rresp_bits_rdata_7 = io_out_rresp_bits_rdata_7; // @[AXIProtocol.scala 15:10:@105141.4]
  assign io_in_rresp_bits_rdata_8 = io_out_rresp_bits_rdata_8; // @[AXIProtocol.scala 15:10:@105142.4]
  assign io_in_rresp_bits_rdata_9 = io_out_rresp_bits_rdata_9; // @[AXIProtocol.scala 15:10:@105143.4]
  assign io_in_rresp_bits_rdata_10 = io_out_rresp_bits_rdata_10; // @[AXIProtocol.scala 15:10:@105144.4]
  assign io_in_rresp_bits_rdata_11 = io_out_rresp_bits_rdata_11; // @[AXIProtocol.scala 15:10:@105145.4]
  assign io_in_rresp_bits_rdata_12 = io_out_rresp_bits_rdata_12; // @[AXIProtocol.scala 15:10:@105146.4]
  assign io_in_rresp_bits_rdata_13 = io_out_rresp_bits_rdata_13; // @[AXIProtocol.scala 15:10:@105147.4]
  assign io_in_rresp_bits_rdata_14 = io_out_rresp_bits_rdata_14; // @[AXIProtocol.scala 15:10:@105148.4]
  assign io_in_rresp_bits_rdata_15 = io_out_rresp_bits_rdata_15; // @[AXIProtocol.scala 15:10:@105149.4]
  assign io_in_rresp_bits_rdata_16 = io_out_rresp_bits_rdata_16; // @[AXIProtocol.scala 15:10:@105150.4]
  assign io_in_rresp_bits_rdata_17 = io_out_rresp_bits_rdata_17; // @[AXIProtocol.scala 15:10:@105151.4]
  assign io_in_rresp_bits_rdata_18 = io_out_rresp_bits_rdata_18; // @[AXIProtocol.scala 15:10:@105152.4]
  assign io_in_rresp_bits_rdata_19 = io_out_rresp_bits_rdata_19; // @[AXIProtocol.scala 15:10:@105153.4]
  assign io_in_rresp_bits_rdata_20 = io_out_rresp_bits_rdata_20; // @[AXIProtocol.scala 15:10:@105154.4]
  assign io_in_rresp_bits_rdata_21 = io_out_rresp_bits_rdata_21; // @[AXIProtocol.scala 15:10:@105155.4]
  assign io_in_rresp_bits_rdata_22 = io_out_rresp_bits_rdata_22; // @[AXIProtocol.scala 15:10:@105156.4]
  assign io_in_rresp_bits_rdata_23 = io_out_rresp_bits_rdata_23; // @[AXIProtocol.scala 15:10:@105157.4]
  assign io_in_rresp_bits_rdata_24 = io_out_rresp_bits_rdata_24; // @[AXIProtocol.scala 15:10:@105158.4]
  assign io_in_rresp_bits_rdata_25 = io_out_rresp_bits_rdata_25; // @[AXIProtocol.scala 15:10:@105159.4]
  assign io_in_rresp_bits_rdata_26 = io_out_rresp_bits_rdata_26; // @[AXIProtocol.scala 15:10:@105160.4]
  assign io_in_rresp_bits_rdata_27 = io_out_rresp_bits_rdata_27; // @[AXIProtocol.scala 15:10:@105161.4]
  assign io_in_rresp_bits_rdata_28 = io_out_rresp_bits_rdata_28; // @[AXIProtocol.scala 15:10:@105162.4]
  assign io_in_rresp_bits_rdata_29 = io_out_rresp_bits_rdata_29; // @[AXIProtocol.scala 15:10:@105163.4]
  assign io_in_rresp_bits_rdata_30 = io_out_rresp_bits_rdata_30; // @[AXIProtocol.scala 15:10:@105164.4]
  assign io_in_rresp_bits_rdata_31 = io_out_rresp_bits_rdata_31; // @[AXIProtocol.scala 15:10:@105165.4]
  assign io_in_rresp_bits_rdata_32 = io_out_rresp_bits_rdata_32; // @[AXIProtocol.scala 15:10:@105166.4]
  assign io_in_rresp_bits_rdata_33 = io_out_rresp_bits_rdata_33; // @[AXIProtocol.scala 15:10:@105167.4]
  assign io_in_rresp_bits_rdata_34 = io_out_rresp_bits_rdata_34; // @[AXIProtocol.scala 15:10:@105168.4]
  assign io_in_rresp_bits_rdata_35 = io_out_rresp_bits_rdata_35; // @[AXIProtocol.scala 15:10:@105169.4]
  assign io_in_rresp_bits_rdata_36 = io_out_rresp_bits_rdata_36; // @[AXIProtocol.scala 15:10:@105170.4]
  assign io_in_rresp_bits_rdata_37 = io_out_rresp_bits_rdata_37; // @[AXIProtocol.scala 15:10:@105171.4]
  assign io_in_rresp_bits_rdata_38 = io_out_rresp_bits_rdata_38; // @[AXIProtocol.scala 15:10:@105172.4]
  assign io_in_rresp_bits_rdata_39 = io_out_rresp_bits_rdata_39; // @[AXIProtocol.scala 15:10:@105173.4]
  assign io_in_rresp_bits_rdata_40 = io_out_rresp_bits_rdata_40; // @[AXIProtocol.scala 15:10:@105174.4]
  assign io_in_rresp_bits_rdata_41 = io_out_rresp_bits_rdata_41; // @[AXIProtocol.scala 15:10:@105175.4]
  assign io_in_rresp_bits_rdata_42 = io_out_rresp_bits_rdata_42; // @[AXIProtocol.scala 15:10:@105176.4]
  assign io_in_rresp_bits_rdata_43 = io_out_rresp_bits_rdata_43; // @[AXIProtocol.scala 15:10:@105177.4]
  assign io_in_rresp_bits_rdata_44 = io_out_rresp_bits_rdata_44; // @[AXIProtocol.scala 15:10:@105178.4]
  assign io_in_rresp_bits_rdata_45 = io_out_rresp_bits_rdata_45; // @[AXIProtocol.scala 15:10:@105179.4]
  assign io_in_rresp_bits_rdata_46 = io_out_rresp_bits_rdata_46; // @[AXIProtocol.scala 15:10:@105180.4]
  assign io_in_rresp_bits_rdata_47 = io_out_rresp_bits_rdata_47; // @[AXIProtocol.scala 15:10:@105181.4]
  assign io_in_rresp_bits_rdata_48 = io_out_rresp_bits_rdata_48; // @[AXIProtocol.scala 15:10:@105182.4]
  assign io_in_rresp_bits_rdata_49 = io_out_rresp_bits_rdata_49; // @[AXIProtocol.scala 15:10:@105183.4]
  assign io_in_rresp_bits_rdata_50 = io_out_rresp_bits_rdata_50; // @[AXIProtocol.scala 15:10:@105184.4]
  assign io_in_rresp_bits_rdata_51 = io_out_rresp_bits_rdata_51; // @[AXIProtocol.scala 15:10:@105185.4]
  assign io_in_rresp_bits_rdata_52 = io_out_rresp_bits_rdata_52; // @[AXIProtocol.scala 15:10:@105186.4]
  assign io_in_rresp_bits_rdata_53 = io_out_rresp_bits_rdata_53; // @[AXIProtocol.scala 15:10:@105187.4]
  assign io_in_rresp_bits_rdata_54 = io_out_rresp_bits_rdata_54; // @[AXIProtocol.scala 15:10:@105188.4]
  assign io_in_rresp_bits_rdata_55 = io_out_rresp_bits_rdata_55; // @[AXIProtocol.scala 15:10:@105189.4]
  assign io_in_rresp_bits_rdata_56 = io_out_rresp_bits_rdata_56; // @[AXIProtocol.scala 15:10:@105190.4]
  assign io_in_rresp_bits_rdata_57 = io_out_rresp_bits_rdata_57; // @[AXIProtocol.scala 15:10:@105191.4]
  assign io_in_rresp_bits_rdata_58 = io_out_rresp_bits_rdata_58; // @[AXIProtocol.scala 15:10:@105192.4]
  assign io_in_rresp_bits_rdata_59 = io_out_rresp_bits_rdata_59; // @[AXIProtocol.scala 15:10:@105193.4]
  assign io_in_rresp_bits_rdata_60 = io_out_rresp_bits_rdata_60; // @[AXIProtocol.scala 15:10:@105194.4]
  assign io_in_rresp_bits_rdata_61 = io_out_rresp_bits_rdata_61; // @[AXIProtocol.scala 15:10:@105195.4]
  assign io_in_rresp_bits_rdata_62 = io_out_rresp_bits_rdata_62; // @[AXIProtocol.scala 15:10:@105196.4]
  assign io_in_rresp_bits_rdata_63 = io_out_rresp_bits_rdata_63; // @[AXIProtocol.scala 15:10:@105197.4]
  assign io_in_rresp_bits_tag = io_out_rresp_bits_tag; // @[AXIProtocol.scala 15:10:@105133.4]
  assign io_in_wresp_valid = io_out_wresp_valid & _T_223; // @[AXIProtocol.scala 15:10:@105131.4 AXIProtocol.scala 46:21:@105385.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 15:10:@105130.4]
  assign io_out_cmd_valid = io_in_cmd_valid; // @[AXIProtocol.scala 15:10:@105336.4]
  assign io_out_cmd_bits_addr = {_T_204,6'h0}; // @[AXIProtocol.scala 15:10:@105335.4 AXIProtocol.scala 29:24:@105354.4]
  assign io_out_cmd_bits_size = lastCmd ? cmdSizeRemaining : 32'h100; // @[AXIProtocol.scala 15:10:@105334.4 AXIProtocol.scala 25:24:@105346.4]
  assign io_out_cmd_bits_rawAddr = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 15:10:@105333.4 AXIProtocol.scala 30:27:@105355.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 15:10:@105332.4]
  assign io_out_cmd_bits_tag = {_T_214,cmdTag_streamID}; // @[AXIProtocol.scala 15:10:@105331.4 FringeBundles.scala 115:32:@105368.4]
  assign io_out_wdata_valid = io_in_wdata_valid; // @[AXIProtocol.scala 15:10:@105329.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 15:10:@105265.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 15:10:@105266.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 15:10:@105267.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 15:10:@105268.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 15:10:@105269.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 15:10:@105270.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 15:10:@105271.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 15:10:@105272.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 15:10:@105273.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 15:10:@105274.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 15:10:@105275.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 15:10:@105276.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 15:10:@105277.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 15:10:@105278.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 15:10:@105279.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 15:10:@105280.4]
  assign io_out_wdata_bits_wdata_16 = io_in_wdata_bits_wdata_16; // @[AXIProtocol.scala 15:10:@105281.4]
  assign io_out_wdata_bits_wdata_17 = io_in_wdata_bits_wdata_17; // @[AXIProtocol.scala 15:10:@105282.4]
  assign io_out_wdata_bits_wdata_18 = io_in_wdata_bits_wdata_18; // @[AXIProtocol.scala 15:10:@105283.4]
  assign io_out_wdata_bits_wdata_19 = io_in_wdata_bits_wdata_19; // @[AXIProtocol.scala 15:10:@105284.4]
  assign io_out_wdata_bits_wdata_20 = io_in_wdata_bits_wdata_20; // @[AXIProtocol.scala 15:10:@105285.4]
  assign io_out_wdata_bits_wdata_21 = io_in_wdata_bits_wdata_21; // @[AXIProtocol.scala 15:10:@105286.4]
  assign io_out_wdata_bits_wdata_22 = io_in_wdata_bits_wdata_22; // @[AXIProtocol.scala 15:10:@105287.4]
  assign io_out_wdata_bits_wdata_23 = io_in_wdata_bits_wdata_23; // @[AXIProtocol.scala 15:10:@105288.4]
  assign io_out_wdata_bits_wdata_24 = io_in_wdata_bits_wdata_24; // @[AXIProtocol.scala 15:10:@105289.4]
  assign io_out_wdata_bits_wdata_25 = io_in_wdata_bits_wdata_25; // @[AXIProtocol.scala 15:10:@105290.4]
  assign io_out_wdata_bits_wdata_26 = io_in_wdata_bits_wdata_26; // @[AXIProtocol.scala 15:10:@105291.4]
  assign io_out_wdata_bits_wdata_27 = io_in_wdata_bits_wdata_27; // @[AXIProtocol.scala 15:10:@105292.4]
  assign io_out_wdata_bits_wdata_28 = io_in_wdata_bits_wdata_28; // @[AXIProtocol.scala 15:10:@105293.4]
  assign io_out_wdata_bits_wdata_29 = io_in_wdata_bits_wdata_29; // @[AXIProtocol.scala 15:10:@105294.4]
  assign io_out_wdata_bits_wdata_30 = io_in_wdata_bits_wdata_30; // @[AXIProtocol.scala 15:10:@105295.4]
  assign io_out_wdata_bits_wdata_31 = io_in_wdata_bits_wdata_31; // @[AXIProtocol.scala 15:10:@105296.4]
  assign io_out_wdata_bits_wdata_32 = io_in_wdata_bits_wdata_32; // @[AXIProtocol.scala 15:10:@105297.4]
  assign io_out_wdata_bits_wdata_33 = io_in_wdata_bits_wdata_33; // @[AXIProtocol.scala 15:10:@105298.4]
  assign io_out_wdata_bits_wdata_34 = io_in_wdata_bits_wdata_34; // @[AXIProtocol.scala 15:10:@105299.4]
  assign io_out_wdata_bits_wdata_35 = io_in_wdata_bits_wdata_35; // @[AXIProtocol.scala 15:10:@105300.4]
  assign io_out_wdata_bits_wdata_36 = io_in_wdata_bits_wdata_36; // @[AXIProtocol.scala 15:10:@105301.4]
  assign io_out_wdata_bits_wdata_37 = io_in_wdata_bits_wdata_37; // @[AXIProtocol.scala 15:10:@105302.4]
  assign io_out_wdata_bits_wdata_38 = io_in_wdata_bits_wdata_38; // @[AXIProtocol.scala 15:10:@105303.4]
  assign io_out_wdata_bits_wdata_39 = io_in_wdata_bits_wdata_39; // @[AXIProtocol.scala 15:10:@105304.4]
  assign io_out_wdata_bits_wdata_40 = io_in_wdata_bits_wdata_40; // @[AXIProtocol.scala 15:10:@105305.4]
  assign io_out_wdata_bits_wdata_41 = io_in_wdata_bits_wdata_41; // @[AXIProtocol.scala 15:10:@105306.4]
  assign io_out_wdata_bits_wdata_42 = io_in_wdata_bits_wdata_42; // @[AXIProtocol.scala 15:10:@105307.4]
  assign io_out_wdata_bits_wdata_43 = io_in_wdata_bits_wdata_43; // @[AXIProtocol.scala 15:10:@105308.4]
  assign io_out_wdata_bits_wdata_44 = io_in_wdata_bits_wdata_44; // @[AXIProtocol.scala 15:10:@105309.4]
  assign io_out_wdata_bits_wdata_45 = io_in_wdata_bits_wdata_45; // @[AXIProtocol.scala 15:10:@105310.4]
  assign io_out_wdata_bits_wdata_46 = io_in_wdata_bits_wdata_46; // @[AXIProtocol.scala 15:10:@105311.4]
  assign io_out_wdata_bits_wdata_47 = io_in_wdata_bits_wdata_47; // @[AXIProtocol.scala 15:10:@105312.4]
  assign io_out_wdata_bits_wdata_48 = io_in_wdata_bits_wdata_48; // @[AXIProtocol.scala 15:10:@105313.4]
  assign io_out_wdata_bits_wdata_49 = io_in_wdata_bits_wdata_49; // @[AXIProtocol.scala 15:10:@105314.4]
  assign io_out_wdata_bits_wdata_50 = io_in_wdata_bits_wdata_50; // @[AXIProtocol.scala 15:10:@105315.4]
  assign io_out_wdata_bits_wdata_51 = io_in_wdata_bits_wdata_51; // @[AXIProtocol.scala 15:10:@105316.4]
  assign io_out_wdata_bits_wdata_52 = io_in_wdata_bits_wdata_52; // @[AXIProtocol.scala 15:10:@105317.4]
  assign io_out_wdata_bits_wdata_53 = io_in_wdata_bits_wdata_53; // @[AXIProtocol.scala 15:10:@105318.4]
  assign io_out_wdata_bits_wdata_54 = io_in_wdata_bits_wdata_54; // @[AXIProtocol.scala 15:10:@105319.4]
  assign io_out_wdata_bits_wdata_55 = io_in_wdata_bits_wdata_55; // @[AXIProtocol.scala 15:10:@105320.4]
  assign io_out_wdata_bits_wdata_56 = io_in_wdata_bits_wdata_56; // @[AXIProtocol.scala 15:10:@105321.4]
  assign io_out_wdata_bits_wdata_57 = io_in_wdata_bits_wdata_57; // @[AXIProtocol.scala 15:10:@105322.4]
  assign io_out_wdata_bits_wdata_58 = io_in_wdata_bits_wdata_58; // @[AXIProtocol.scala 15:10:@105323.4]
  assign io_out_wdata_bits_wdata_59 = io_in_wdata_bits_wdata_59; // @[AXIProtocol.scala 15:10:@105324.4]
  assign io_out_wdata_bits_wdata_60 = io_in_wdata_bits_wdata_60; // @[AXIProtocol.scala 15:10:@105325.4]
  assign io_out_wdata_bits_wdata_61 = io_in_wdata_bits_wdata_61; // @[AXIProtocol.scala 15:10:@105326.4]
  assign io_out_wdata_bits_wdata_62 = io_in_wdata_bits_wdata_62; // @[AXIProtocol.scala 15:10:@105327.4]
  assign io_out_wdata_bits_wdata_63 = io_in_wdata_bits_wdata_63; // @[AXIProtocol.scala 15:10:@105328.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 15:10:@105201.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 15:10:@105202.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 15:10:@105203.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 15:10:@105204.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 15:10:@105205.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 15:10:@105206.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 15:10:@105207.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 15:10:@105208.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 15:10:@105209.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 15:10:@105210.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 15:10:@105211.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 15:10:@105212.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 15:10:@105213.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 15:10:@105214.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 15:10:@105215.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 15:10:@105216.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 15:10:@105217.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 15:10:@105218.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 15:10:@105219.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 15:10:@105220.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 15:10:@105221.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 15:10:@105222.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 15:10:@105223.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 15:10:@105224.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 15:10:@105225.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 15:10:@105226.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 15:10:@105227.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 15:10:@105228.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 15:10:@105229.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 15:10:@105230.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 15:10:@105231.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 15:10:@105232.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 15:10:@105233.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 15:10:@105234.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 15:10:@105235.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 15:10:@105236.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 15:10:@105237.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 15:10:@105238.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 15:10:@105239.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 15:10:@105240.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 15:10:@105241.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 15:10:@105242.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 15:10:@105243.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 15:10:@105244.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 15:10:@105245.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 15:10:@105246.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 15:10:@105247.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 15:10:@105248.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 15:10:@105249.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 15:10:@105250.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 15:10:@105251.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 15:10:@105252.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 15:10:@105253.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 15:10:@105254.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 15:10:@105255.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 15:10:@105256.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 15:10:@105257.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 15:10:@105258.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 15:10:@105259.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 15:10:@105260.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 15:10:@105261.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 15:10:@105262.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 15:10:@105263.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 15:10:@105264.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 15:10:@105199.4]
  assign io_out_wresp_ready = _T_223 ? io_in_wresp_ready : 1'h1; // @[AXIProtocol.scala 15:10:@105132.4 AXIProtocol.scala 47:22:@105387.4]
  assign cmdSizeCounter_clock = clock; // @[:@105339.4]
  assign cmdSizeCounter_reset = reset; // @[:@105340.4]
  assign cmdSizeCounter_io_reset = lastCmd & cmdIssue; // @[AXIProtocol.scala 40:27:@105372.4]
  assign cmdSizeCounter_io_enable = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 41:28:@105373.4]
  assign cmdSizeCounter_io_stride = 32'h100; // @[AXIProtocol.scala 42:28:@105374.4]
endmodule
module AXICmdIssue( // @[:@105407.2]
  input         clock, // @[:@105408.4]
  input         reset, // @[:@105409.4]
  output        io_in_cmd_ready, // @[:@105410.4]
  input         io_in_cmd_valid, // @[:@105410.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@105410.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@105410.4]
  input  [63:0] io_in_cmd_bits_rawAddr, // @[:@105410.4]
  input         io_in_cmd_bits_isWr, // @[:@105410.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@105410.4]
  output        io_in_wdata_ready, // @[:@105410.4]
  input         io_in_wdata_valid, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_0, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_1, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_2, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_3, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_4, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_5, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_6, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_7, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_8, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_9, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_10, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_11, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_12, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_13, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_14, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_15, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_16, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_17, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_18, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_19, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_20, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_21, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_22, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_23, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_24, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_25, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_26, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_27, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_28, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_29, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_30, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_31, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_32, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_33, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_34, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_35, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_36, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_37, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_38, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_39, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_40, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_41, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_42, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_43, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_44, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_45, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_46, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_47, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_48, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_49, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_50, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_51, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_52, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_53, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_54, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_55, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_56, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_57, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_58, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_59, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_60, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_61, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_62, // @[:@105410.4]
  input  [7:0]  io_in_wdata_bits_wdata_63, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@105410.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@105410.4]
  input         io_in_rresp_ready, // @[:@105410.4]
  output        io_in_rresp_valid, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_0, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_1, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_2, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_3, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_4, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_5, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_6, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_7, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_8, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_9, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_10, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_11, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_12, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_13, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_14, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_15, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_16, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_17, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_18, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_19, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_20, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_21, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_22, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_23, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_24, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_25, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_26, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_27, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_28, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_29, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_30, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_31, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_32, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_33, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_34, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_35, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_36, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_37, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_38, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_39, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_40, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_41, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_42, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_43, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_44, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_45, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_46, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_47, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_48, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_49, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_50, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_51, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_52, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_53, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_54, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_55, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_56, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_57, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_58, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_59, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_60, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_61, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_62, // @[:@105410.4]
  output [7:0]  io_in_rresp_bits_rdata_63, // @[:@105410.4]
  output [31:0] io_in_rresp_bits_tag, // @[:@105410.4]
  input         io_in_wresp_ready, // @[:@105410.4]
  output        io_in_wresp_valid, // @[:@105410.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@105410.4]
  input         io_out_cmd_ready, // @[:@105410.4]
  output        io_out_cmd_valid, // @[:@105410.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@105410.4]
  output [31:0] io_out_cmd_bits_size, // @[:@105410.4]
  output [63:0] io_out_cmd_bits_rawAddr, // @[:@105410.4]
  output        io_out_cmd_bits_isWr, // @[:@105410.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@105410.4]
  input         io_out_wdata_ready, // @[:@105410.4]
  output        io_out_wdata_valid, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_0, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_1, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_2, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_3, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_4, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_5, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_6, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_7, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_8, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_9, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_10, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_11, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_12, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_13, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_14, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_15, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_16, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_17, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_18, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_19, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_20, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_21, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_22, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_23, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_24, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_25, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_26, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_27, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_28, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_29, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_30, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_31, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_32, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_33, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_34, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_35, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_36, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_37, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_38, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_39, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_40, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_41, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_42, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_43, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_44, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_45, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_46, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_47, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_48, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_49, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_50, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_51, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_52, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_53, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_54, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_55, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_56, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_57, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_58, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_59, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_60, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_61, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_62, // @[:@105410.4]
  output [7:0]  io_out_wdata_bits_wdata_63, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@105410.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@105410.4]
  output        io_out_wdata_bits_wlast, // @[:@105410.4]
  output        io_out_rresp_ready, // @[:@105410.4]
  input         io_out_rresp_valid, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_0, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_1, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_2, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_3, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_4, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_5, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_6, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_7, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_8, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_9, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_10, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_11, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_12, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_13, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_14, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_15, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_16, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_17, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_18, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_19, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_20, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_21, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_22, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_23, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_24, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_25, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_26, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_27, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_28, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_29, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_30, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_31, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_32, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_33, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_34, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_35, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_36, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_37, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_38, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_39, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_40, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_41, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_42, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_43, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_44, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_45, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_46, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_47, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_48, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_49, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_50, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_51, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_52, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_53, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_54, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_55, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_56, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_57, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_58, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_59, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_60, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_61, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_62, // @[:@105410.4]
  input  [7:0]  io_out_rresp_bits_rdata_63, // @[:@105410.4]
  input  [31:0] io_out_rresp_bits_tag, // @[:@105410.4]
  output        io_out_wresp_ready, // @[:@105410.4]
  input         io_out_wresp_valid, // @[:@105410.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@105410.4]
);
  wire  wdataCounter_clock; // @[AXIProtocol.scala 59:28:@105620.4]
  wire  wdataCounter_reset; // @[AXIProtocol.scala 59:28:@105620.4]
  wire  wdataCounter_io_reset; // @[AXIProtocol.scala 59:28:@105620.4]
  wire  wdataCounter_io_enable; // @[AXIProtocol.scala 59:28:@105620.4]
  wire [31:0] wdataCounter_io_stride; // @[AXIProtocol.scala 59:28:@105620.4]
  wire [31:0] wdataCounter_io_out; // @[AXIProtocol.scala 59:28:@105620.4]
  wire [31:0] wdataCounter_io_next; // @[AXIProtocol.scala 59:28:@105620.4]
  reg  writeIssued; // @[AXIProtocol.scala 61:28:@105623.4]
  reg [31:0] _RAND_0;
  wire  dramCmdIssue; // @[AXIProtocol.scala 63:39:@105624.4]
  wire  dramWriteIssue; // @[AXIProtocol.scala 64:43:@105625.4]
  wire  _T_201; // @[AXIProtocol.scala 68:54:@105626.4]
  wire  wlast; // @[AXIProtocol.scala 68:30:@105627.4]
  wire  _T_203; // @[AXIProtocol.scala 72:28:@105633.6]
  wire  _GEN_0; // @[AXIProtocol.scala 72:40:@105634.6]
  wire  _GEN_1; // @[AXIProtocol.scala 70:15:@105629.4]
  wire  _T_208; // @[AXIProtocol.scala 84:55:@105643.4]
  wire  _T_210; // @[AXIProtocol.scala 84:44:@105644.4]
  Counter_112 wdataCounter ( // @[AXIProtocol.scala 59:28:@105620.4]
    .clock(wdataCounter_clock),
    .reset(wdataCounter_reset),
    .io_reset(wdataCounter_io_reset),
    .io_enable(wdataCounter_io_enable),
    .io_stride(wdataCounter_io_stride),
    .io_out(wdataCounter_io_out),
    .io_next(wdataCounter_io_next)
  );
  assign dramCmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 63:39:@105624.4]
  assign dramWriteIssue = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 64:43:@105625.4]
  assign _T_201 = wdataCounter_io_next == io_in_cmd_bits_size; // @[AXIProtocol.scala 68:54:@105626.4]
  assign wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 68:30:@105627.4]
  assign _T_203 = dramCmdIssue & io_in_cmd_bits_isWr; // @[AXIProtocol.scala 72:28:@105633.6]
  assign _GEN_0 = _T_203 ? 1'h1 : writeIssued; // @[AXIProtocol.scala 72:40:@105634.6]
  assign _GEN_1 = wlast ? 1'h0 : _GEN_0; // @[AXIProtocol.scala 70:15:@105629.4]
  assign _T_208 = writeIssued == 1'h0; // @[AXIProtocol.scala 84:55:@105643.4]
  assign _T_210 = io_in_cmd_bits_isWr ? _T_208 : 1'h1; // @[AXIProtocol.scala 84:44:@105644.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? wlast : dramCmdIssue; // @[AXIProtocol.scala 56:10:@105619.4 AXIProtocol.scala 81:19:@105641.4]
  assign io_in_wdata_ready = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 56:10:@105612.4 AXIProtocol.scala 82:21:@105642.4]
  assign io_in_rresp_valid = io_out_rresp_valid; // @[AXIProtocol.scala 56:10:@105480.4]
  assign io_in_rresp_bits_rdata_0 = io_out_rresp_bits_rdata_0; // @[AXIProtocol.scala 56:10:@105416.4]
  assign io_in_rresp_bits_rdata_1 = io_out_rresp_bits_rdata_1; // @[AXIProtocol.scala 56:10:@105417.4]
  assign io_in_rresp_bits_rdata_2 = io_out_rresp_bits_rdata_2; // @[AXIProtocol.scala 56:10:@105418.4]
  assign io_in_rresp_bits_rdata_3 = io_out_rresp_bits_rdata_3; // @[AXIProtocol.scala 56:10:@105419.4]
  assign io_in_rresp_bits_rdata_4 = io_out_rresp_bits_rdata_4; // @[AXIProtocol.scala 56:10:@105420.4]
  assign io_in_rresp_bits_rdata_5 = io_out_rresp_bits_rdata_5; // @[AXIProtocol.scala 56:10:@105421.4]
  assign io_in_rresp_bits_rdata_6 = io_out_rresp_bits_rdata_6; // @[AXIProtocol.scala 56:10:@105422.4]
  assign io_in_rresp_bits_rdata_7 = io_out_rresp_bits_rdata_7; // @[AXIProtocol.scala 56:10:@105423.4]
  assign io_in_rresp_bits_rdata_8 = io_out_rresp_bits_rdata_8; // @[AXIProtocol.scala 56:10:@105424.4]
  assign io_in_rresp_bits_rdata_9 = io_out_rresp_bits_rdata_9; // @[AXIProtocol.scala 56:10:@105425.4]
  assign io_in_rresp_bits_rdata_10 = io_out_rresp_bits_rdata_10; // @[AXIProtocol.scala 56:10:@105426.4]
  assign io_in_rresp_bits_rdata_11 = io_out_rresp_bits_rdata_11; // @[AXIProtocol.scala 56:10:@105427.4]
  assign io_in_rresp_bits_rdata_12 = io_out_rresp_bits_rdata_12; // @[AXIProtocol.scala 56:10:@105428.4]
  assign io_in_rresp_bits_rdata_13 = io_out_rresp_bits_rdata_13; // @[AXIProtocol.scala 56:10:@105429.4]
  assign io_in_rresp_bits_rdata_14 = io_out_rresp_bits_rdata_14; // @[AXIProtocol.scala 56:10:@105430.4]
  assign io_in_rresp_bits_rdata_15 = io_out_rresp_bits_rdata_15; // @[AXIProtocol.scala 56:10:@105431.4]
  assign io_in_rresp_bits_rdata_16 = io_out_rresp_bits_rdata_16; // @[AXIProtocol.scala 56:10:@105432.4]
  assign io_in_rresp_bits_rdata_17 = io_out_rresp_bits_rdata_17; // @[AXIProtocol.scala 56:10:@105433.4]
  assign io_in_rresp_bits_rdata_18 = io_out_rresp_bits_rdata_18; // @[AXIProtocol.scala 56:10:@105434.4]
  assign io_in_rresp_bits_rdata_19 = io_out_rresp_bits_rdata_19; // @[AXIProtocol.scala 56:10:@105435.4]
  assign io_in_rresp_bits_rdata_20 = io_out_rresp_bits_rdata_20; // @[AXIProtocol.scala 56:10:@105436.4]
  assign io_in_rresp_bits_rdata_21 = io_out_rresp_bits_rdata_21; // @[AXIProtocol.scala 56:10:@105437.4]
  assign io_in_rresp_bits_rdata_22 = io_out_rresp_bits_rdata_22; // @[AXIProtocol.scala 56:10:@105438.4]
  assign io_in_rresp_bits_rdata_23 = io_out_rresp_bits_rdata_23; // @[AXIProtocol.scala 56:10:@105439.4]
  assign io_in_rresp_bits_rdata_24 = io_out_rresp_bits_rdata_24; // @[AXIProtocol.scala 56:10:@105440.4]
  assign io_in_rresp_bits_rdata_25 = io_out_rresp_bits_rdata_25; // @[AXIProtocol.scala 56:10:@105441.4]
  assign io_in_rresp_bits_rdata_26 = io_out_rresp_bits_rdata_26; // @[AXIProtocol.scala 56:10:@105442.4]
  assign io_in_rresp_bits_rdata_27 = io_out_rresp_bits_rdata_27; // @[AXIProtocol.scala 56:10:@105443.4]
  assign io_in_rresp_bits_rdata_28 = io_out_rresp_bits_rdata_28; // @[AXIProtocol.scala 56:10:@105444.4]
  assign io_in_rresp_bits_rdata_29 = io_out_rresp_bits_rdata_29; // @[AXIProtocol.scala 56:10:@105445.4]
  assign io_in_rresp_bits_rdata_30 = io_out_rresp_bits_rdata_30; // @[AXIProtocol.scala 56:10:@105446.4]
  assign io_in_rresp_bits_rdata_31 = io_out_rresp_bits_rdata_31; // @[AXIProtocol.scala 56:10:@105447.4]
  assign io_in_rresp_bits_rdata_32 = io_out_rresp_bits_rdata_32; // @[AXIProtocol.scala 56:10:@105448.4]
  assign io_in_rresp_bits_rdata_33 = io_out_rresp_bits_rdata_33; // @[AXIProtocol.scala 56:10:@105449.4]
  assign io_in_rresp_bits_rdata_34 = io_out_rresp_bits_rdata_34; // @[AXIProtocol.scala 56:10:@105450.4]
  assign io_in_rresp_bits_rdata_35 = io_out_rresp_bits_rdata_35; // @[AXIProtocol.scala 56:10:@105451.4]
  assign io_in_rresp_bits_rdata_36 = io_out_rresp_bits_rdata_36; // @[AXIProtocol.scala 56:10:@105452.4]
  assign io_in_rresp_bits_rdata_37 = io_out_rresp_bits_rdata_37; // @[AXIProtocol.scala 56:10:@105453.4]
  assign io_in_rresp_bits_rdata_38 = io_out_rresp_bits_rdata_38; // @[AXIProtocol.scala 56:10:@105454.4]
  assign io_in_rresp_bits_rdata_39 = io_out_rresp_bits_rdata_39; // @[AXIProtocol.scala 56:10:@105455.4]
  assign io_in_rresp_bits_rdata_40 = io_out_rresp_bits_rdata_40; // @[AXIProtocol.scala 56:10:@105456.4]
  assign io_in_rresp_bits_rdata_41 = io_out_rresp_bits_rdata_41; // @[AXIProtocol.scala 56:10:@105457.4]
  assign io_in_rresp_bits_rdata_42 = io_out_rresp_bits_rdata_42; // @[AXIProtocol.scala 56:10:@105458.4]
  assign io_in_rresp_bits_rdata_43 = io_out_rresp_bits_rdata_43; // @[AXIProtocol.scala 56:10:@105459.4]
  assign io_in_rresp_bits_rdata_44 = io_out_rresp_bits_rdata_44; // @[AXIProtocol.scala 56:10:@105460.4]
  assign io_in_rresp_bits_rdata_45 = io_out_rresp_bits_rdata_45; // @[AXIProtocol.scala 56:10:@105461.4]
  assign io_in_rresp_bits_rdata_46 = io_out_rresp_bits_rdata_46; // @[AXIProtocol.scala 56:10:@105462.4]
  assign io_in_rresp_bits_rdata_47 = io_out_rresp_bits_rdata_47; // @[AXIProtocol.scala 56:10:@105463.4]
  assign io_in_rresp_bits_rdata_48 = io_out_rresp_bits_rdata_48; // @[AXIProtocol.scala 56:10:@105464.4]
  assign io_in_rresp_bits_rdata_49 = io_out_rresp_bits_rdata_49; // @[AXIProtocol.scala 56:10:@105465.4]
  assign io_in_rresp_bits_rdata_50 = io_out_rresp_bits_rdata_50; // @[AXIProtocol.scala 56:10:@105466.4]
  assign io_in_rresp_bits_rdata_51 = io_out_rresp_bits_rdata_51; // @[AXIProtocol.scala 56:10:@105467.4]
  assign io_in_rresp_bits_rdata_52 = io_out_rresp_bits_rdata_52; // @[AXIProtocol.scala 56:10:@105468.4]
  assign io_in_rresp_bits_rdata_53 = io_out_rresp_bits_rdata_53; // @[AXIProtocol.scala 56:10:@105469.4]
  assign io_in_rresp_bits_rdata_54 = io_out_rresp_bits_rdata_54; // @[AXIProtocol.scala 56:10:@105470.4]
  assign io_in_rresp_bits_rdata_55 = io_out_rresp_bits_rdata_55; // @[AXIProtocol.scala 56:10:@105471.4]
  assign io_in_rresp_bits_rdata_56 = io_out_rresp_bits_rdata_56; // @[AXIProtocol.scala 56:10:@105472.4]
  assign io_in_rresp_bits_rdata_57 = io_out_rresp_bits_rdata_57; // @[AXIProtocol.scala 56:10:@105473.4]
  assign io_in_rresp_bits_rdata_58 = io_out_rresp_bits_rdata_58; // @[AXIProtocol.scala 56:10:@105474.4]
  assign io_in_rresp_bits_rdata_59 = io_out_rresp_bits_rdata_59; // @[AXIProtocol.scala 56:10:@105475.4]
  assign io_in_rresp_bits_rdata_60 = io_out_rresp_bits_rdata_60; // @[AXIProtocol.scala 56:10:@105476.4]
  assign io_in_rresp_bits_rdata_61 = io_out_rresp_bits_rdata_61; // @[AXIProtocol.scala 56:10:@105477.4]
  assign io_in_rresp_bits_rdata_62 = io_out_rresp_bits_rdata_62; // @[AXIProtocol.scala 56:10:@105478.4]
  assign io_in_rresp_bits_rdata_63 = io_out_rresp_bits_rdata_63; // @[AXIProtocol.scala 56:10:@105479.4]
  assign io_in_rresp_bits_tag = io_out_rresp_bits_tag; // @[AXIProtocol.scala 56:10:@105415.4]
  assign io_in_wresp_valid = io_out_wresp_valid; // @[AXIProtocol.scala 56:10:@105413.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 56:10:@105412.4]
  assign io_out_cmd_valid = io_in_cmd_valid & _T_210; // @[AXIProtocol.scala 56:10:@105618.4 AXIProtocol.scala 84:20:@105646.4]
  assign io_out_cmd_bits_addr = io_in_cmd_bits_addr; // @[AXIProtocol.scala 56:10:@105617.4]
  assign io_out_cmd_bits_size = io_in_cmd_bits_size; // @[AXIProtocol.scala 56:10:@105616.4]
  assign io_out_cmd_bits_rawAddr = io_in_cmd_bits_rawAddr; // @[AXIProtocol.scala 56:10:@105615.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 56:10:@105614.4]
  assign io_out_cmd_bits_tag = io_in_cmd_bits_tag; // @[AXIProtocol.scala 56:10:@105613.4]
  assign io_out_wdata_valid = io_in_wdata_valid & writeIssued; // @[AXIProtocol.scala 56:10:@105611.4 AXIProtocol.scala 86:22:@105648.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 56:10:@105547.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 56:10:@105548.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 56:10:@105549.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 56:10:@105550.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 56:10:@105551.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 56:10:@105552.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 56:10:@105553.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 56:10:@105554.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 56:10:@105555.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 56:10:@105556.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 56:10:@105557.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 56:10:@105558.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 56:10:@105559.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 56:10:@105560.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 56:10:@105561.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 56:10:@105562.4]
  assign io_out_wdata_bits_wdata_16 = io_in_wdata_bits_wdata_16; // @[AXIProtocol.scala 56:10:@105563.4]
  assign io_out_wdata_bits_wdata_17 = io_in_wdata_bits_wdata_17; // @[AXIProtocol.scala 56:10:@105564.4]
  assign io_out_wdata_bits_wdata_18 = io_in_wdata_bits_wdata_18; // @[AXIProtocol.scala 56:10:@105565.4]
  assign io_out_wdata_bits_wdata_19 = io_in_wdata_bits_wdata_19; // @[AXIProtocol.scala 56:10:@105566.4]
  assign io_out_wdata_bits_wdata_20 = io_in_wdata_bits_wdata_20; // @[AXIProtocol.scala 56:10:@105567.4]
  assign io_out_wdata_bits_wdata_21 = io_in_wdata_bits_wdata_21; // @[AXIProtocol.scala 56:10:@105568.4]
  assign io_out_wdata_bits_wdata_22 = io_in_wdata_bits_wdata_22; // @[AXIProtocol.scala 56:10:@105569.4]
  assign io_out_wdata_bits_wdata_23 = io_in_wdata_bits_wdata_23; // @[AXIProtocol.scala 56:10:@105570.4]
  assign io_out_wdata_bits_wdata_24 = io_in_wdata_bits_wdata_24; // @[AXIProtocol.scala 56:10:@105571.4]
  assign io_out_wdata_bits_wdata_25 = io_in_wdata_bits_wdata_25; // @[AXIProtocol.scala 56:10:@105572.4]
  assign io_out_wdata_bits_wdata_26 = io_in_wdata_bits_wdata_26; // @[AXIProtocol.scala 56:10:@105573.4]
  assign io_out_wdata_bits_wdata_27 = io_in_wdata_bits_wdata_27; // @[AXIProtocol.scala 56:10:@105574.4]
  assign io_out_wdata_bits_wdata_28 = io_in_wdata_bits_wdata_28; // @[AXIProtocol.scala 56:10:@105575.4]
  assign io_out_wdata_bits_wdata_29 = io_in_wdata_bits_wdata_29; // @[AXIProtocol.scala 56:10:@105576.4]
  assign io_out_wdata_bits_wdata_30 = io_in_wdata_bits_wdata_30; // @[AXIProtocol.scala 56:10:@105577.4]
  assign io_out_wdata_bits_wdata_31 = io_in_wdata_bits_wdata_31; // @[AXIProtocol.scala 56:10:@105578.4]
  assign io_out_wdata_bits_wdata_32 = io_in_wdata_bits_wdata_32; // @[AXIProtocol.scala 56:10:@105579.4]
  assign io_out_wdata_bits_wdata_33 = io_in_wdata_bits_wdata_33; // @[AXIProtocol.scala 56:10:@105580.4]
  assign io_out_wdata_bits_wdata_34 = io_in_wdata_bits_wdata_34; // @[AXIProtocol.scala 56:10:@105581.4]
  assign io_out_wdata_bits_wdata_35 = io_in_wdata_bits_wdata_35; // @[AXIProtocol.scala 56:10:@105582.4]
  assign io_out_wdata_bits_wdata_36 = io_in_wdata_bits_wdata_36; // @[AXIProtocol.scala 56:10:@105583.4]
  assign io_out_wdata_bits_wdata_37 = io_in_wdata_bits_wdata_37; // @[AXIProtocol.scala 56:10:@105584.4]
  assign io_out_wdata_bits_wdata_38 = io_in_wdata_bits_wdata_38; // @[AXIProtocol.scala 56:10:@105585.4]
  assign io_out_wdata_bits_wdata_39 = io_in_wdata_bits_wdata_39; // @[AXIProtocol.scala 56:10:@105586.4]
  assign io_out_wdata_bits_wdata_40 = io_in_wdata_bits_wdata_40; // @[AXIProtocol.scala 56:10:@105587.4]
  assign io_out_wdata_bits_wdata_41 = io_in_wdata_bits_wdata_41; // @[AXIProtocol.scala 56:10:@105588.4]
  assign io_out_wdata_bits_wdata_42 = io_in_wdata_bits_wdata_42; // @[AXIProtocol.scala 56:10:@105589.4]
  assign io_out_wdata_bits_wdata_43 = io_in_wdata_bits_wdata_43; // @[AXIProtocol.scala 56:10:@105590.4]
  assign io_out_wdata_bits_wdata_44 = io_in_wdata_bits_wdata_44; // @[AXIProtocol.scala 56:10:@105591.4]
  assign io_out_wdata_bits_wdata_45 = io_in_wdata_bits_wdata_45; // @[AXIProtocol.scala 56:10:@105592.4]
  assign io_out_wdata_bits_wdata_46 = io_in_wdata_bits_wdata_46; // @[AXIProtocol.scala 56:10:@105593.4]
  assign io_out_wdata_bits_wdata_47 = io_in_wdata_bits_wdata_47; // @[AXIProtocol.scala 56:10:@105594.4]
  assign io_out_wdata_bits_wdata_48 = io_in_wdata_bits_wdata_48; // @[AXIProtocol.scala 56:10:@105595.4]
  assign io_out_wdata_bits_wdata_49 = io_in_wdata_bits_wdata_49; // @[AXIProtocol.scala 56:10:@105596.4]
  assign io_out_wdata_bits_wdata_50 = io_in_wdata_bits_wdata_50; // @[AXIProtocol.scala 56:10:@105597.4]
  assign io_out_wdata_bits_wdata_51 = io_in_wdata_bits_wdata_51; // @[AXIProtocol.scala 56:10:@105598.4]
  assign io_out_wdata_bits_wdata_52 = io_in_wdata_bits_wdata_52; // @[AXIProtocol.scala 56:10:@105599.4]
  assign io_out_wdata_bits_wdata_53 = io_in_wdata_bits_wdata_53; // @[AXIProtocol.scala 56:10:@105600.4]
  assign io_out_wdata_bits_wdata_54 = io_in_wdata_bits_wdata_54; // @[AXIProtocol.scala 56:10:@105601.4]
  assign io_out_wdata_bits_wdata_55 = io_in_wdata_bits_wdata_55; // @[AXIProtocol.scala 56:10:@105602.4]
  assign io_out_wdata_bits_wdata_56 = io_in_wdata_bits_wdata_56; // @[AXIProtocol.scala 56:10:@105603.4]
  assign io_out_wdata_bits_wdata_57 = io_in_wdata_bits_wdata_57; // @[AXIProtocol.scala 56:10:@105604.4]
  assign io_out_wdata_bits_wdata_58 = io_in_wdata_bits_wdata_58; // @[AXIProtocol.scala 56:10:@105605.4]
  assign io_out_wdata_bits_wdata_59 = io_in_wdata_bits_wdata_59; // @[AXIProtocol.scala 56:10:@105606.4]
  assign io_out_wdata_bits_wdata_60 = io_in_wdata_bits_wdata_60; // @[AXIProtocol.scala 56:10:@105607.4]
  assign io_out_wdata_bits_wdata_61 = io_in_wdata_bits_wdata_61; // @[AXIProtocol.scala 56:10:@105608.4]
  assign io_out_wdata_bits_wdata_62 = io_in_wdata_bits_wdata_62; // @[AXIProtocol.scala 56:10:@105609.4]
  assign io_out_wdata_bits_wdata_63 = io_in_wdata_bits_wdata_63; // @[AXIProtocol.scala 56:10:@105610.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 56:10:@105483.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 56:10:@105484.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 56:10:@105485.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 56:10:@105486.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 56:10:@105487.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 56:10:@105488.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 56:10:@105489.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 56:10:@105490.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 56:10:@105491.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 56:10:@105492.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 56:10:@105493.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 56:10:@105494.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 56:10:@105495.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 56:10:@105496.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 56:10:@105497.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 56:10:@105498.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 56:10:@105499.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 56:10:@105500.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 56:10:@105501.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 56:10:@105502.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 56:10:@105503.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 56:10:@105504.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 56:10:@105505.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 56:10:@105506.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 56:10:@105507.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 56:10:@105508.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 56:10:@105509.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 56:10:@105510.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 56:10:@105511.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 56:10:@105512.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 56:10:@105513.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 56:10:@105514.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 56:10:@105515.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 56:10:@105516.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 56:10:@105517.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 56:10:@105518.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 56:10:@105519.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 56:10:@105520.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 56:10:@105521.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 56:10:@105522.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 56:10:@105523.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 56:10:@105524.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 56:10:@105525.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 56:10:@105526.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 56:10:@105527.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 56:10:@105528.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 56:10:@105529.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 56:10:@105530.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 56:10:@105531.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 56:10:@105532.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 56:10:@105533.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 56:10:@105534.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 56:10:@105535.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 56:10:@105536.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 56:10:@105537.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 56:10:@105538.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 56:10:@105539.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 56:10:@105540.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 56:10:@105541.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 56:10:@105542.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 56:10:@105543.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 56:10:@105544.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 56:10:@105545.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 56:10:@105546.4]
  assign io_out_wdata_bits_wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 56:10:@105482.4 AXIProtocol.scala 87:27:@105649.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 56:10:@105481.4]
  assign io_out_wresp_ready = io_in_wresp_ready; // @[AXIProtocol.scala 56:10:@105414.4]
  assign wdataCounter_clock = clock; // @[:@105621.4]
  assign wdataCounter_reset = reset; // @[:@105622.4]
  assign wdataCounter_io_reset = dramWriteIssue & _T_201; // @[AXIProtocol.scala 76:25:@105637.4]
  assign wdataCounter_io_enable = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 77:26:@105638.4]
  assign wdataCounter_io_stride = 32'h1; // @[AXIProtocol.scala 78:26:@105639.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeIssued = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      writeIssued <= 1'h0;
    end else begin
      if (wlast) begin
        writeIssued <= 1'h0;
      end else begin
        if (_T_203) begin
          writeIssued <= 1'h1;
        end
      end
    end
  end
endmodule
module DRAMArbiter( // @[:@105651.2]
  input         clock, // @[:@105652.4]
  input         reset, // @[:@105653.4]
  input         io_enable, // @[:@105654.4]
  output        io_app_loads_0_cmd_ready, // @[:@105654.4]
  input         io_app_loads_0_cmd_valid, // @[:@105654.4]
  input  [63:0] io_app_loads_0_cmd_bits_addr, // @[:@105654.4]
  input  [31:0] io_app_loads_0_cmd_bits_size, // @[:@105654.4]
  input         io_app_loads_0_data_ready, // @[:@105654.4]
  output        io_app_loads_0_data_valid, // @[:@105654.4]
  output [31:0] io_app_loads_0_data_bits_rdata_0, // @[:@105654.4]
  output        io_app_stores_0_cmd_ready, // @[:@105654.4]
  input         io_app_stores_0_cmd_valid, // @[:@105654.4]
  input  [63:0] io_app_stores_0_cmd_bits_addr, // @[:@105654.4]
  input  [31:0] io_app_stores_0_cmd_bits_size, // @[:@105654.4]
  output        io_app_stores_0_data_ready, // @[:@105654.4]
  input         io_app_stores_0_data_valid, // @[:@105654.4]
  input  [31:0] io_app_stores_0_data_bits_wdata_0, // @[:@105654.4]
  input         io_app_stores_0_data_bits_wstrb, // @[:@105654.4]
  input         io_app_stores_0_wresp_ready, // @[:@105654.4]
  output        io_app_stores_0_wresp_valid, // @[:@105654.4]
  output        io_app_stores_0_wresp_bits, // @[:@105654.4]
  input         io_dram_cmd_ready, // @[:@105654.4]
  output        io_dram_cmd_valid, // @[:@105654.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@105654.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@105654.4]
  output [63:0] io_dram_cmd_bits_rawAddr, // @[:@105654.4]
  output        io_dram_cmd_bits_isWr, // @[:@105654.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@105654.4]
  input         io_dram_wdata_ready, // @[:@105654.4]
  output        io_dram_wdata_valid, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_0, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_1, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_2, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_3, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_4, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_5, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_6, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_7, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_8, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_9, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_10, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_11, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_12, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_13, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_14, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_15, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_16, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_17, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_18, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_19, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_20, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_21, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_22, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_23, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_24, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_25, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_26, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_27, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_28, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_29, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_30, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_31, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_32, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_33, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_34, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_35, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_36, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_37, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_38, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_39, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_40, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_41, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_42, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_43, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_44, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_45, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_46, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_47, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_48, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_49, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_50, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_51, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_52, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_53, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_54, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_55, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_56, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_57, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_58, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_59, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_60, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_61, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_62, // @[:@105654.4]
  output [7:0]  io_dram_wdata_bits_wdata_63, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@105654.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@105654.4]
  output        io_dram_wdata_bits_wlast, // @[:@105654.4]
  output        io_dram_rresp_ready, // @[:@105654.4]
  input         io_dram_rresp_valid, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_0, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_1, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_2, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_3, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_4, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_5, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_6, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_7, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_8, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_9, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_10, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_11, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_12, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_13, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_14, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_15, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_16, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_17, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_18, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_19, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_20, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_21, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_22, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_23, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_24, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_25, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_26, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_27, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_28, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_29, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_30, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_31, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_32, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_33, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_34, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_35, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_36, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_37, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_38, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_39, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_40, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_41, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_42, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_43, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_44, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_45, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_46, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_47, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_48, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_49, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_50, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_51, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_52, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_53, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_54, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_55, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_56, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_57, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_58, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_59, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_60, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_61, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_62, // @[:@105654.4]
  input  [7:0]  io_dram_rresp_bits_rdata_63, // @[:@105654.4]
  input  [31:0] io_dram_rresp_bits_tag, // @[:@105654.4]
  output        io_dram_wresp_ready, // @[:@105654.4]
  input         io_dram_wresp_valid, // @[:@105654.4]
  input  [31:0] io_dram_wresp_bits_tag, // @[:@105654.4]
  output [31:0] io_debugSignals_0, // @[:@105654.4]
  output [31:0] io_debugSignals_1, // @[:@105654.4]
  output [31:0] io_debugSignals_2, // @[:@105654.4]
  output [31:0] io_debugSignals_3, // @[:@105654.4]
  output [31:0] io_debugSignals_4, // @[:@105654.4]
  output [31:0] io_debugSignals_5, // @[:@105654.4]
  output [31:0] io_debugSignals_6, // @[:@105654.4]
  output [31:0] io_debugSignals_7, // @[:@105654.4]
  output [31:0] io_debugSignals_8, // @[:@105654.4]
  output [31:0] io_debugSignals_9, // @[:@105654.4]
  output [31:0] io_debugSignals_10, // @[:@105654.4]
  output [31:0] io_debugSignals_11, // @[:@105654.4]
  output [31:0] io_debugSignals_12, // @[:@105654.4]
  output [31:0] io_debugSignals_13, // @[:@105654.4]
  output [31:0] io_debugSignals_14, // @[:@105654.4]
  output [31:0] io_debugSignals_15, // @[:@105654.4]
  output [31:0] io_debugSignals_16, // @[:@105654.4]
  output [31:0] io_debugSignals_17, // @[:@105654.4]
  output [31:0] io_debugSignals_18, // @[:@105654.4]
  output [31:0] io_debugSignals_19, // @[:@105654.4]
  output [31:0] io_debugSignals_20, // @[:@105654.4]
  output [31:0] io_debugSignals_21, // @[:@105654.4]
  output [31:0] io_debugSignals_22, // @[:@105654.4]
  output [31:0] io_debugSignals_23, // @[:@105654.4]
  output [31:0] io_debugSignals_24, // @[:@105654.4]
  output [31:0] io_debugSignals_25, // @[:@105654.4]
  output [31:0] io_debugSignals_26, // @[:@105654.4]
  output [31:0] io_debugSignals_27, // @[:@105654.4]
  output [31:0] io_debugSignals_28, // @[:@105654.4]
  output [31:0] io_debugSignals_29, // @[:@105654.4]
  output [31:0] io_debugSignals_30, // @[:@105654.4]
  output [31:0] io_debugSignals_41 // @[:@105654.4]
);
  wire  StreamControllerLoad_clock; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire  StreamControllerLoad_reset; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire  StreamControllerLoad_io_dram_cmd_ready; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire  StreamControllerLoad_io_dram_cmd_valid; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [63:0] StreamControllerLoad_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [31:0] StreamControllerLoad_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire  StreamControllerLoad_io_dram_rresp_ready; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire  StreamControllerLoad_io_dram_rresp_valid; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_0; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_1; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_2; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_3; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_4; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_5; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_6; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_7; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_8; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_9; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_10; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_11; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_12; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_13; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_14; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_15; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_16; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_17; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_18; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_19; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_20; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_21; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_22; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_23; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_24; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_25; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_26; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_27; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_28; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_29; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_30; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_31; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_32; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_33; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_34; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_35; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_36; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_37; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_38; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_39; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_40; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_41; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_42; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_43; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_44; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_45; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_46; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_47; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_48; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_49; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_50; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_51; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_52; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_53; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_54; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_55; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_56; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_57; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_58; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_59; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_60; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_61; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_62; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [7:0] StreamControllerLoad_io_dram_rresp_bits_rdata_63; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire  StreamControllerLoad_io_load_cmd_ready; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire  StreamControllerLoad_io_load_cmd_valid; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [63:0] StreamControllerLoad_io_load_cmd_bits_addr; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [31:0] StreamControllerLoad_io_load_cmd_bits_size; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire  StreamControllerLoad_io_load_data_ready; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire  StreamControllerLoad_io_load_data_valid; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire [31:0] StreamControllerLoad_io_load_data_bits_rdata_0; // @[DRAMArbiter.scala 60:21:@106813.4]
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_16; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_17; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_18; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_19; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_20; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_21; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_22; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_23; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_24; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_25; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_26; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_27; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_28; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_29; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_30; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_31; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_32; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_33; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_34; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_35; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_36; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_37; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_38; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_39; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_40; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_41; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_42; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_43; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_44; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_45; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_46; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_47; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_48; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_49; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_50; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_51; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_52; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_53; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_54; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_55; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_56; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_57; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_58; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_59; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_60; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_61; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_62; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [7:0] StreamControllerStore_io_dram_wdata_bits_wdata_63; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@106823.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_0_rresp_valid; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_0; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_1; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_2; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_3; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_4; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_5; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_6; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_7; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_8; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_9; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_10; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_11; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_12; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_13; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_14; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_15; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_16; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_17; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_18; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_19; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_20; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_21; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_22; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_23; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_24; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_25; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_26; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_27; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_28; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_29; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_30; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_31; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_32; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_33; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_34; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_35; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_36; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_37; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_38; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_39; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_40; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_41; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_42; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_43; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_44; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_45; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_46; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_47; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_48; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_49; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_50; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_51; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_52; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_53; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_54; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_55; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_56; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_57; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_58; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_59; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_60; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_61; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_62; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_0_rresp_bits_rdata_63; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_cmd_ready; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_cmd_valid; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [63:0] StreamArbiter_io_app_1_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [31:0] StreamArbiter_io_app_1_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_ready; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_valid; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_16; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_17; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_18; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_19; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_20; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_21; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_22; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_23; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_24; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_25; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_26; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_27; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_28; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_29; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_30; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_31; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_32; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_33; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_34; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_35; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_36; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_37; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_38; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_39; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_40; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_41; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_42; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_43; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_44; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_45; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_46; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_47; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_48; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_49; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_50; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_51; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_52; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_53; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_54; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_55; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_56; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_57; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_58; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_59; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_60; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_61; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_62; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_app_1_wdata_bits_wdata_63; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wresp_ready; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_app_1_wresp_valid; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_16; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_17; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_18; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_19; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_20; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_21; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_22; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_23; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_24; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_25; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_26; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_27; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_28; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_29; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_30; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_31; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_32; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_33; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_34; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_35; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_36; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_37; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_38; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_39; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_40; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_41; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_42; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_43; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_44; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_45; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_46; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_47; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_48; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_49; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_50; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_51; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_52; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_53; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_54; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_55; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_56; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_57; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_58; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_59; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_60; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_61; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_62; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_wdata_bits_wdata_63; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_rresp_valid; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_0; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_1; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_2; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_3; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_4; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_5; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_6; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_7; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_8; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_9; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_10; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_11; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_12; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_13; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_14; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_15; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_16; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_17; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_18; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_19; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_20; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_21; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_22; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_23; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_24; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_25; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_26; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_27; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_28; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_29; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_30; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_31; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_32; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_33; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_34; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_35; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_36; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_37; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_38; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_39; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_40; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_41; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_42; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_43; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_44; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_45; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_46; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_47; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_48; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_49; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_50; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_51; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_52; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_53; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_54; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_55; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_56; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_57; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_58; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_59; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_60; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_61; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_62; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [7:0] StreamArbiter_io_dram_rresp_bits_rdata_63; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_tag; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@106837.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_16; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_17; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_18; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_19; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_20; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_21; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_22; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_23; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_24; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_25; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_26; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_27; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_28; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_29; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_30; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_31; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_32; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_33; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_34; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_35; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_36; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_37; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_38; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_39; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_40; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_41; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_42; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_43; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_44; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_45; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_46; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_47; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_48; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_49; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_50; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_51; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_52; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_53; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_54; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_55; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_56; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_57; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_58; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_59; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_60; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_61; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_62; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_wdata_bits_wdata_63; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_rresp_valid; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_0; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_1; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_2; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_3; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_4; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_5; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_6; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_7; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_8; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_9; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_10; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_11; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_12; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_13; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_14; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_15; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_16; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_17; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_18; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_19; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_20; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_21; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_22; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_23; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_24; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_25; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_26; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_27; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_28; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_29; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_30; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_31; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_32; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_33; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_34; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_35; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_36; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_37; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_38; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_39; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_40; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_41; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_42; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_43; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_44; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_45; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_46; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_47; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_48; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_49; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_50; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_51; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_52; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_53; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_54; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_55; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_56; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_57; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_58; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_59; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_60; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_61; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_62; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_in_rresp_bits_rdata_63; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_tag; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_rawAddr; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_16; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_17; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_18; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_19; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_20; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_21; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_22; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_23; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_24; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_25; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_26; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_27; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_28; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_29; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_30; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_31; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_32; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_33; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_34; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_35; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_36; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_37; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_38; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_39; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_40; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_41; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_42; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_43; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_44; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_45; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_46; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_47; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_48; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_49; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_50; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_51; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_52; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_53; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_54; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_55; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_56; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_57; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_58; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_59; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_60; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_61; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_62; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_wdata_bits_wdata_63; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_rresp_valid; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_0; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_1; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_2; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_3; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_4; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_5; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_6; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_7; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_8; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_9; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_10; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_11; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_12; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_13; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_14; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_15; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_16; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_17; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_18; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_19; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_20; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_21; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_22; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_23; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_24; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_25; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_26; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_27; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_28; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_29; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_30; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_31; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_32; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_33; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_34; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_35; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_36; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_37; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_38; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_39; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_40; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_41; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_42; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_43; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_44; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_45; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_46; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_47; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_48; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_49; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_50; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_51; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_52; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_53; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_54; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_55; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_56; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_57; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_58; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_59; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_60; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_61; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_62; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [7:0] AXICmdSplit_io_out_rresp_bits_rdata_63; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_tag; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@107673.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_rawAddr; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_16; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_17; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_18; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_19; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_20; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_21; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_22; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_23; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_24; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_25; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_26; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_27; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_28; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_29; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_30; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_31; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_32; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_33; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_34; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_35; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_36; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_37; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_38; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_39; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_40; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_41; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_42; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_43; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_44; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_45; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_46; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_47; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_48; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_49; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_50; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_51; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_52; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_53; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_54; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_55; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_56; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_57; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_58; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_59; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_60; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_61; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_62; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_wdata_bits_wdata_63; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_rresp_valid; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_0; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_1; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_2; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_3; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_4; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_5; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_6; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_7; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_8; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_9; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_10; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_11; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_12; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_13; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_14; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_15; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_16; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_17; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_18; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_19; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_20; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_21; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_22; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_23; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_24; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_25; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_26; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_27; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_28; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_29; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_30; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_31; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_32; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_33; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_34; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_35; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_36; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_37; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_38; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_39; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_40; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_41; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_42; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_43; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_44; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_45; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_46; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_47; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_48; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_49; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_50; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_51; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_52; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_53; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_54; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_55; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_56; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_57; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_58; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_59; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_60; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_61; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_62; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_in_rresp_bits_rdata_63; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_tag; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_rawAddr; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_16; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_17; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_18; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_19; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_20; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_21; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_22; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_23; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_24; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_25; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_26; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_27; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_28; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_29; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_30; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_31; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_32; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_33; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_34; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_35; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_36; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_37; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_38; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_39; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_40; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_41; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_42; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_43; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_44; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_45; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_46; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_47; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_48; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_49; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_50; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_51; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_52; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_53; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_54; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_55; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_56; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_57; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_58; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_59; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_60; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_61; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_62; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_wdata_bits_wdata_63; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_rresp_valid; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_0; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_1; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_2; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_3; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_4; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_5; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_6; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_7; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_8; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_9; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_10; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_11; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_12; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_13; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_14; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_15; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_16; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_17; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_18; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_19; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_20; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_21; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_22; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_23; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_24; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_25; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_26; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_27; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_28; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_29; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_30; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_31; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_32; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_33; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_34; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_35; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_36; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_37; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_38; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_39; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_40; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_41; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_42; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_43; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_44; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_45; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_46; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_47; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_48; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_49; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_50; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_51; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_52; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_53; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_54; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_55; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_56; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_57; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_58; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_59; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_60; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_61; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_62; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [7:0] AXICmdIssue_io_out_rresp_bits_rdata_63; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_tag; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@107884.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@107884.4]
  reg [63:0] _T_2028; // @[DRAMArbiter.scala 121:24:@108307.4]
  reg [63:0] _RAND_0;
  wire [64:0] _T_2030; // @[DRAMArbiter.scala 123:18:@108309.6]
  wire [63:0] _T_2031; // @[DRAMArbiter.scala 123:18:@108310.6]
  wire [63:0] _GEN_0; // @[DRAMArbiter.scala 122:19:@108308.4]
  wire  _T_2032; // @[DRAMArbiter.scala 139:60:@108314.4]
  wire  _T_2039; // @[DRAMArbiter.scala 140:57:@108321.4]
  reg [63:0] _T_2042; // @[DRAMArbiter.scala 121:24:@108322.4]
  reg [63:0] _RAND_1;
  wire [64:0] _T_2044; // @[DRAMArbiter.scala 123:18:@108324.6]
  wire [63:0] _T_2045; // @[DRAMArbiter.scala 123:18:@108325.6]
  wire [63:0] _GEN_2; // @[DRAMArbiter.scala 122:19:@108323.4]
  wire  _T_2046; // @[DRAMArbiter.scala 141:70:@108328.4]
  reg [63:0] _T_2049; // @[DRAMArbiter.scala 121:24:@108329.4]
  reg [63:0] _RAND_2;
  wire [64:0] _T_2051; // @[DRAMArbiter.scala 123:18:@108331.6]
  wire [63:0] _T_2052; // @[DRAMArbiter.scala 123:18:@108332.6]
  wire [63:0] _GEN_3; // @[DRAMArbiter.scala 122:19:@108330.4]
  wire  _T_2053; // @[DRAMArbiter.scala 144:52:@108336.4]
  reg [63:0] _T_2056; // @[DRAMArbiter.scala 121:24:@108337.4]
  reg [63:0] _RAND_3;
  wire [64:0] _T_2058; // @[DRAMArbiter.scala 123:18:@108339.6]
  wire [63:0] _T_2059; // @[DRAMArbiter.scala 123:18:@108340.6]
  wire [63:0] _GEN_4; // @[DRAMArbiter.scala 122:19:@108338.4]
  wire  _T_2062; // @[DRAMArbiter.scala 145:74:@108345.4]
  wire  _T_2063; // @[DRAMArbiter.scala 145:72:@108346.4]
  reg [63:0] _T_2066; // @[DRAMArbiter.scala 121:24:@108347.4]
  reg [63:0] _RAND_4;
  wire [64:0] _T_2068; // @[DRAMArbiter.scala 123:18:@108349.6]
  wire [63:0] _T_2069; // @[DRAMArbiter.scala 123:18:@108350.6]
  wire [63:0] _GEN_5; // @[DRAMArbiter.scala 122:19:@108348.4]
  wire  _T_2071; // @[DRAMArbiter.scala 146:72:@108355.4]
  reg [63:0] _T_2074; // @[DRAMArbiter.scala 121:24:@108356.4]
  reg [63:0] _RAND_5;
  wire [64:0] _T_2076; // @[DRAMArbiter.scala 123:18:@108358.6]
  wire [63:0] _T_2077; // @[DRAMArbiter.scala 123:18:@108359.6]
  wire [63:0] _GEN_6; // @[DRAMArbiter.scala 122:19:@108357.4]
  wire  _T_2078; // @[DRAMArbiter.scala 150:59:@108363.4]
  wire  _T_2079; // @[DRAMArbiter.scala 150:76:@108364.4]
  reg [63:0] _T_2082; // @[DRAMArbiter.scala 121:24:@108365.4]
  reg [63:0] _RAND_6;
  wire [64:0] _T_2084; // @[DRAMArbiter.scala 123:18:@108367.6]
  wire [63:0] _T_2085; // @[DRAMArbiter.scala 123:18:@108368.6]
  wire [63:0] _GEN_7; // @[DRAMArbiter.scala 122:19:@108366.4]
  wire  _T_2086; // @[DRAMArbiter.scala 156:60:@108372.4]
  wire  _T_2087; // @[DRAMArbiter.scala 156:78:@108373.4]
  reg [63:0] _T_2090; // @[DRAMArbiter.scala 121:24:@108374.4]
  reg [63:0] _RAND_7;
  wire [64:0] _T_2092; // @[DRAMArbiter.scala 123:18:@108376.6]
  wire [63:0] _T_2093; // @[DRAMArbiter.scala 123:18:@108377.6]
  wire [63:0] _GEN_8; // @[DRAMArbiter.scala 122:19:@108375.4]
  reg [63:0] _T_2097; // @[DRAMArbiter.scala 121:24:@108382.4]
  reg [63:0] _RAND_8;
  wire [64:0] _T_2099; // @[DRAMArbiter.scala 123:18:@108384.6]
  wire [63:0] _T_2100; // @[DRAMArbiter.scala 123:18:@108385.6]
  wire [63:0] _GEN_9; // @[DRAMArbiter.scala 122:19:@108383.4]
  wire  _T_2102; // @[DRAMArbiter.scala 161:56:@108389.4]
  wire  _T_2103; // @[DRAMArbiter.scala 161:54:@108390.4]
  reg [63:0] _T_2106; // @[DRAMArbiter.scala 121:24:@108391.4]
  reg [63:0] _RAND_9;
  wire [64:0] _T_2108; // @[DRAMArbiter.scala 123:18:@108393.6]
  wire [63:0] _T_2109; // @[DRAMArbiter.scala 123:18:@108394.6]
  wire [63:0] _GEN_10; // @[DRAMArbiter.scala 122:19:@108392.4]
  wire  _T_2111; // @[DRAMArbiter.scala 162:34:@108398.4]
  wire  _T_2112; // @[DRAMArbiter.scala 162:55:@108399.4]
  reg [63:0] _T_2115; // @[DRAMArbiter.scala 121:24:@108400.4]
  reg [63:0] _RAND_10;
  wire [64:0] _T_2117; // @[DRAMArbiter.scala 123:18:@108402.6]
  wire [63:0] _T_2118; // @[DRAMArbiter.scala 123:18:@108403.6]
  wire [63:0] _GEN_11; // @[DRAMArbiter.scala 122:19:@108401.4]
  wire [7:0] _T_2125; // @[FringeBundles.scala 132:28:@108411.4]
  wire  _T_2129; // @[DRAMArbiter.scala 165:116:@108417.4]
  wire  _T_2130; // @[DRAMArbiter.scala 165:78:@108418.4]
  reg [63:0] _T_2133; // @[DRAMArbiter.scala 121:24:@108419.4]
  reg [63:0] _RAND_11;
  wire [64:0] _T_2135; // @[DRAMArbiter.scala 123:18:@108421.6]
  wire [63:0] _T_2136; // @[DRAMArbiter.scala 123:18:@108422.6]
  wire [63:0] _GEN_12; // @[DRAMArbiter.scala 122:19:@108420.4]
  wire  _T_2137; // @[DRAMArbiter.scala 167:54:@108426.4]
  reg [63:0] _T_2140; // @[DRAMArbiter.scala 121:24:@108427.4]
  reg [63:0] _RAND_12;
  wire [64:0] _T_2142; // @[DRAMArbiter.scala 123:18:@108429.6]
  wire [63:0] _T_2143; // @[DRAMArbiter.scala 123:18:@108430.6]
  wire [63:0] _GEN_13; // @[DRAMArbiter.scala 122:19:@108428.4]
  wire  _T_2145; // @[DRAMArbiter.scala 168:56:@108434.4]
  wire  _T_2146; // @[DRAMArbiter.scala 168:54:@108435.4]
  reg [63:0] _T_2149; // @[DRAMArbiter.scala 121:24:@108436.4]
  reg [63:0] _RAND_13;
  wire [64:0] _T_2151; // @[DRAMArbiter.scala 123:18:@108438.6]
  wire [63:0] _T_2152; // @[DRAMArbiter.scala 123:18:@108439.6]
  wire [63:0] _GEN_14; // @[DRAMArbiter.scala 122:19:@108437.4]
  wire  _T_2154; // @[DRAMArbiter.scala 169:34:@108443.4]
  wire  _T_2155; // @[DRAMArbiter.scala 169:55:@108444.4]
  reg [63:0] _T_2158; // @[DRAMArbiter.scala 121:24:@108445.4]
  reg [63:0] _RAND_14;
  wire [64:0] _T_2160; // @[DRAMArbiter.scala 123:18:@108447.6]
  wire [63:0] _T_2161; // @[DRAMArbiter.scala 123:18:@108448.6]
  wire [63:0] _GEN_15; // @[DRAMArbiter.scala 122:19:@108446.4]
  wire [7:0] _T_2168; // @[FringeBundles.scala 140:28:@108456.4]
  wire  _T_2172; // @[DRAMArbiter.scala 172:116:@108462.4]
  wire  _T_2173; // @[DRAMArbiter.scala 172:78:@108463.4]
  reg [63:0] _T_2176; // @[DRAMArbiter.scala 121:24:@108464.4]
  reg [63:0] _RAND_15;
  wire [64:0] _T_2178; // @[DRAMArbiter.scala 123:18:@108466.6]
  wire [63:0] _T_2179; // @[DRAMArbiter.scala 123:18:@108467.6]
  wire [63:0] _GEN_16; // @[DRAMArbiter.scala 122:19:@108465.4]
  wire  _T_2180; // @[DRAMArbiter.scala 176:70:@108471.4]
  reg [63:0] _T_2182; // @[DRAMArbiter.scala 129:25:@108472.4]
  reg [63:0] _RAND_16;
  wire [63:0] _GEN_17; // @[DRAMArbiter.scala 130:19:@108473.4]
  reg [31:0] _T_2185; // @[DRAMArbiter.scala 129:25:@108478.4]
  reg [31:0] _RAND_17;
  wire [31:0] _GEN_18; // @[DRAMArbiter.scala 130:19:@108479.4]
  reg [7:0] _T_2188; // @[DRAMArbiter.scala 129:25:@108484.4]
  reg [31:0] _RAND_18;
  wire [7:0] _GEN_19; // @[DRAMArbiter.scala 130:19:@108485.4]
  reg  _T_2191; // @[DRAMArbiter.scala 129:25:@108490.4]
  reg [31:0] _RAND_19;
  wire  _GEN_20; // @[DRAMArbiter.scala 130:19:@108491.4]
  wire  _T_2194; // @[DRAMArbiter.scala 180:115:@108496.4]
  wire  _T_2195; // @[DRAMArbiter.scala 180:102:@108497.4]
  reg [7:0] _T_2197; // @[DRAMArbiter.scala 129:25:@108498.4]
  reg [31:0] _RAND_20;
  wire [7:0] _GEN_21; // @[DRAMArbiter.scala 130:19:@108499.4]
  reg  _T_2203; // @[DRAMArbiter.scala 129:25:@108506.4]
  reg [31:0] _RAND_21;
  wire  _GEN_22; // @[DRAMArbiter.scala 130:19:@108507.4]
  wire  _T_2206; // @[DRAMArbiter.scala 182:115:@108512.4]
  wire  _T_2207; // @[DRAMArbiter.scala 182:102:@108513.4]
  reg [7:0] _T_2209; // @[DRAMArbiter.scala 129:25:@108514.4]
  reg [31:0] _RAND_22;
  wire [7:0] _GEN_23; // @[DRAMArbiter.scala 130:19:@108515.4]
  reg  _T_2215; // @[DRAMArbiter.scala 129:25:@108522.4]
  reg [31:0] _RAND_23;
  wire  _GEN_24; // @[DRAMArbiter.scala 130:19:@108523.4]
  wire  _T_2216; // @[DRAMArbiter.scala 184:92:@108527.4]
  reg [63:0] _T_2218; // @[DRAMArbiter.scala 129:25:@108528.4]
  reg [63:0] _RAND_24;
  wire [63:0] _GEN_25; // @[DRAMArbiter.scala 130:19:@108529.4]
  reg [31:0] _T_2221; // @[DRAMArbiter.scala 129:25:@108534.4]
  reg [31:0] _RAND_25;
  wire [31:0] _GEN_26; // @[DRAMArbiter.scala 130:19:@108535.4]
  reg [31:0] _T_2224; // @[DRAMArbiter.scala 129:25:@108540.4]
  reg [31:0] _RAND_26;
  wire [31:0] _GEN_27; // @[DRAMArbiter.scala 130:19:@108541.4]
  reg  _T_2227; // @[DRAMArbiter.scala 129:25:@108546.4]
  reg [31:0] _RAND_27;
  wire  _GEN_28; // @[DRAMArbiter.scala 130:19:@108547.4]
  wire  _T_2230; // @[DRAMArbiter.scala 188:148:@108552.4]
  wire  _T_2231; // @[DRAMArbiter.scala 188:132:@108553.4]
  reg [31:0] _T_2233; // @[DRAMArbiter.scala 129:25:@108554.4]
  reg [31:0] _RAND_28;
  wire [31:0] _GEN_29; // @[DRAMArbiter.scala 130:19:@108555.4]
  reg  _T_2239; // @[DRAMArbiter.scala 129:25:@108562.4]
  reg [31:0] _RAND_29;
  wire  _GEN_30; // @[DRAMArbiter.scala 130:19:@108563.4]
  wire  _T_2242; // @[DRAMArbiter.scala 190:148:@108568.4]
  wire  _T_2243; // @[DRAMArbiter.scala 190:132:@108569.4]
  reg [31:0] _T_2245; // @[DRAMArbiter.scala 129:25:@108570.4]
  reg [31:0] _RAND_30;
  wire [31:0] _GEN_31; // @[DRAMArbiter.scala 130:19:@108571.4]
  reg  _T_2251; // @[DRAMArbiter.scala 129:25:@108578.4]
  reg [31:0] _RAND_31;
  wire  _GEN_32; // @[DRAMArbiter.scala 130:19:@108579.4]
  reg [63:0] _T_2323; // @[DRAMArbiter.scala 121:24:@108660.4]
  reg [63:0] _RAND_32;
  wire [64:0] _T_2325; // @[DRAMArbiter.scala 123:18:@108662.6]
  wire [63:0] _T_2326; // @[DRAMArbiter.scala 123:18:@108663.6]
  StreamControllerLoad StreamControllerLoad ( // @[DRAMArbiter.scala 60:21:@106813.4]
    .clock(StreamControllerLoad_clock),
    .reset(StreamControllerLoad_reset),
    .io_dram_cmd_ready(StreamControllerLoad_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerLoad_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerLoad_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerLoad_io_dram_cmd_bits_size),
    .io_dram_rresp_ready(StreamControllerLoad_io_dram_rresp_ready),
    .io_dram_rresp_valid(StreamControllerLoad_io_dram_rresp_valid),
    .io_dram_rresp_bits_rdata_0(StreamControllerLoad_io_dram_rresp_bits_rdata_0),
    .io_dram_rresp_bits_rdata_1(StreamControllerLoad_io_dram_rresp_bits_rdata_1),
    .io_dram_rresp_bits_rdata_2(StreamControllerLoad_io_dram_rresp_bits_rdata_2),
    .io_dram_rresp_bits_rdata_3(StreamControllerLoad_io_dram_rresp_bits_rdata_3),
    .io_dram_rresp_bits_rdata_4(StreamControllerLoad_io_dram_rresp_bits_rdata_4),
    .io_dram_rresp_bits_rdata_5(StreamControllerLoad_io_dram_rresp_bits_rdata_5),
    .io_dram_rresp_bits_rdata_6(StreamControllerLoad_io_dram_rresp_bits_rdata_6),
    .io_dram_rresp_bits_rdata_7(StreamControllerLoad_io_dram_rresp_bits_rdata_7),
    .io_dram_rresp_bits_rdata_8(StreamControllerLoad_io_dram_rresp_bits_rdata_8),
    .io_dram_rresp_bits_rdata_9(StreamControllerLoad_io_dram_rresp_bits_rdata_9),
    .io_dram_rresp_bits_rdata_10(StreamControllerLoad_io_dram_rresp_bits_rdata_10),
    .io_dram_rresp_bits_rdata_11(StreamControllerLoad_io_dram_rresp_bits_rdata_11),
    .io_dram_rresp_bits_rdata_12(StreamControllerLoad_io_dram_rresp_bits_rdata_12),
    .io_dram_rresp_bits_rdata_13(StreamControllerLoad_io_dram_rresp_bits_rdata_13),
    .io_dram_rresp_bits_rdata_14(StreamControllerLoad_io_dram_rresp_bits_rdata_14),
    .io_dram_rresp_bits_rdata_15(StreamControllerLoad_io_dram_rresp_bits_rdata_15),
    .io_dram_rresp_bits_rdata_16(StreamControllerLoad_io_dram_rresp_bits_rdata_16),
    .io_dram_rresp_bits_rdata_17(StreamControllerLoad_io_dram_rresp_bits_rdata_17),
    .io_dram_rresp_bits_rdata_18(StreamControllerLoad_io_dram_rresp_bits_rdata_18),
    .io_dram_rresp_bits_rdata_19(StreamControllerLoad_io_dram_rresp_bits_rdata_19),
    .io_dram_rresp_bits_rdata_20(StreamControllerLoad_io_dram_rresp_bits_rdata_20),
    .io_dram_rresp_bits_rdata_21(StreamControllerLoad_io_dram_rresp_bits_rdata_21),
    .io_dram_rresp_bits_rdata_22(StreamControllerLoad_io_dram_rresp_bits_rdata_22),
    .io_dram_rresp_bits_rdata_23(StreamControllerLoad_io_dram_rresp_bits_rdata_23),
    .io_dram_rresp_bits_rdata_24(StreamControllerLoad_io_dram_rresp_bits_rdata_24),
    .io_dram_rresp_bits_rdata_25(StreamControllerLoad_io_dram_rresp_bits_rdata_25),
    .io_dram_rresp_bits_rdata_26(StreamControllerLoad_io_dram_rresp_bits_rdata_26),
    .io_dram_rresp_bits_rdata_27(StreamControllerLoad_io_dram_rresp_bits_rdata_27),
    .io_dram_rresp_bits_rdata_28(StreamControllerLoad_io_dram_rresp_bits_rdata_28),
    .io_dram_rresp_bits_rdata_29(StreamControllerLoad_io_dram_rresp_bits_rdata_29),
    .io_dram_rresp_bits_rdata_30(StreamControllerLoad_io_dram_rresp_bits_rdata_30),
    .io_dram_rresp_bits_rdata_31(StreamControllerLoad_io_dram_rresp_bits_rdata_31),
    .io_dram_rresp_bits_rdata_32(StreamControllerLoad_io_dram_rresp_bits_rdata_32),
    .io_dram_rresp_bits_rdata_33(StreamControllerLoad_io_dram_rresp_bits_rdata_33),
    .io_dram_rresp_bits_rdata_34(StreamControllerLoad_io_dram_rresp_bits_rdata_34),
    .io_dram_rresp_bits_rdata_35(StreamControllerLoad_io_dram_rresp_bits_rdata_35),
    .io_dram_rresp_bits_rdata_36(StreamControllerLoad_io_dram_rresp_bits_rdata_36),
    .io_dram_rresp_bits_rdata_37(StreamControllerLoad_io_dram_rresp_bits_rdata_37),
    .io_dram_rresp_bits_rdata_38(StreamControllerLoad_io_dram_rresp_bits_rdata_38),
    .io_dram_rresp_bits_rdata_39(StreamControllerLoad_io_dram_rresp_bits_rdata_39),
    .io_dram_rresp_bits_rdata_40(StreamControllerLoad_io_dram_rresp_bits_rdata_40),
    .io_dram_rresp_bits_rdata_41(StreamControllerLoad_io_dram_rresp_bits_rdata_41),
    .io_dram_rresp_bits_rdata_42(StreamControllerLoad_io_dram_rresp_bits_rdata_42),
    .io_dram_rresp_bits_rdata_43(StreamControllerLoad_io_dram_rresp_bits_rdata_43),
    .io_dram_rresp_bits_rdata_44(StreamControllerLoad_io_dram_rresp_bits_rdata_44),
    .io_dram_rresp_bits_rdata_45(StreamControllerLoad_io_dram_rresp_bits_rdata_45),
    .io_dram_rresp_bits_rdata_46(StreamControllerLoad_io_dram_rresp_bits_rdata_46),
    .io_dram_rresp_bits_rdata_47(StreamControllerLoad_io_dram_rresp_bits_rdata_47),
    .io_dram_rresp_bits_rdata_48(StreamControllerLoad_io_dram_rresp_bits_rdata_48),
    .io_dram_rresp_bits_rdata_49(StreamControllerLoad_io_dram_rresp_bits_rdata_49),
    .io_dram_rresp_bits_rdata_50(StreamControllerLoad_io_dram_rresp_bits_rdata_50),
    .io_dram_rresp_bits_rdata_51(StreamControllerLoad_io_dram_rresp_bits_rdata_51),
    .io_dram_rresp_bits_rdata_52(StreamControllerLoad_io_dram_rresp_bits_rdata_52),
    .io_dram_rresp_bits_rdata_53(StreamControllerLoad_io_dram_rresp_bits_rdata_53),
    .io_dram_rresp_bits_rdata_54(StreamControllerLoad_io_dram_rresp_bits_rdata_54),
    .io_dram_rresp_bits_rdata_55(StreamControllerLoad_io_dram_rresp_bits_rdata_55),
    .io_dram_rresp_bits_rdata_56(StreamControllerLoad_io_dram_rresp_bits_rdata_56),
    .io_dram_rresp_bits_rdata_57(StreamControllerLoad_io_dram_rresp_bits_rdata_57),
    .io_dram_rresp_bits_rdata_58(StreamControllerLoad_io_dram_rresp_bits_rdata_58),
    .io_dram_rresp_bits_rdata_59(StreamControllerLoad_io_dram_rresp_bits_rdata_59),
    .io_dram_rresp_bits_rdata_60(StreamControllerLoad_io_dram_rresp_bits_rdata_60),
    .io_dram_rresp_bits_rdata_61(StreamControllerLoad_io_dram_rresp_bits_rdata_61),
    .io_dram_rresp_bits_rdata_62(StreamControllerLoad_io_dram_rresp_bits_rdata_62),
    .io_dram_rresp_bits_rdata_63(StreamControllerLoad_io_dram_rresp_bits_rdata_63),
    .io_load_cmd_ready(StreamControllerLoad_io_load_cmd_ready),
    .io_load_cmd_valid(StreamControllerLoad_io_load_cmd_valid),
    .io_load_cmd_bits_addr(StreamControllerLoad_io_load_cmd_bits_addr),
    .io_load_cmd_bits_size(StreamControllerLoad_io_load_cmd_bits_size),
    .io_load_data_ready(StreamControllerLoad_io_load_data_ready),
    .io_load_data_valid(StreamControllerLoad_io_load_data_valid),
    .io_load_data_bits_rdata_0(StreamControllerLoad_io_load_data_bits_rdata_0)
  );
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@106823.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wdata_16(StreamControllerStore_io_dram_wdata_bits_wdata_16),
    .io_dram_wdata_bits_wdata_17(StreamControllerStore_io_dram_wdata_bits_wdata_17),
    .io_dram_wdata_bits_wdata_18(StreamControllerStore_io_dram_wdata_bits_wdata_18),
    .io_dram_wdata_bits_wdata_19(StreamControllerStore_io_dram_wdata_bits_wdata_19),
    .io_dram_wdata_bits_wdata_20(StreamControllerStore_io_dram_wdata_bits_wdata_20),
    .io_dram_wdata_bits_wdata_21(StreamControllerStore_io_dram_wdata_bits_wdata_21),
    .io_dram_wdata_bits_wdata_22(StreamControllerStore_io_dram_wdata_bits_wdata_22),
    .io_dram_wdata_bits_wdata_23(StreamControllerStore_io_dram_wdata_bits_wdata_23),
    .io_dram_wdata_bits_wdata_24(StreamControllerStore_io_dram_wdata_bits_wdata_24),
    .io_dram_wdata_bits_wdata_25(StreamControllerStore_io_dram_wdata_bits_wdata_25),
    .io_dram_wdata_bits_wdata_26(StreamControllerStore_io_dram_wdata_bits_wdata_26),
    .io_dram_wdata_bits_wdata_27(StreamControllerStore_io_dram_wdata_bits_wdata_27),
    .io_dram_wdata_bits_wdata_28(StreamControllerStore_io_dram_wdata_bits_wdata_28),
    .io_dram_wdata_bits_wdata_29(StreamControllerStore_io_dram_wdata_bits_wdata_29),
    .io_dram_wdata_bits_wdata_30(StreamControllerStore_io_dram_wdata_bits_wdata_30),
    .io_dram_wdata_bits_wdata_31(StreamControllerStore_io_dram_wdata_bits_wdata_31),
    .io_dram_wdata_bits_wdata_32(StreamControllerStore_io_dram_wdata_bits_wdata_32),
    .io_dram_wdata_bits_wdata_33(StreamControllerStore_io_dram_wdata_bits_wdata_33),
    .io_dram_wdata_bits_wdata_34(StreamControllerStore_io_dram_wdata_bits_wdata_34),
    .io_dram_wdata_bits_wdata_35(StreamControllerStore_io_dram_wdata_bits_wdata_35),
    .io_dram_wdata_bits_wdata_36(StreamControllerStore_io_dram_wdata_bits_wdata_36),
    .io_dram_wdata_bits_wdata_37(StreamControllerStore_io_dram_wdata_bits_wdata_37),
    .io_dram_wdata_bits_wdata_38(StreamControllerStore_io_dram_wdata_bits_wdata_38),
    .io_dram_wdata_bits_wdata_39(StreamControllerStore_io_dram_wdata_bits_wdata_39),
    .io_dram_wdata_bits_wdata_40(StreamControllerStore_io_dram_wdata_bits_wdata_40),
    .io_dram_wdata_bits_wdata_41(StreamControllerStore_io_dram_wdata_bits_wdata_41),
    .io_dram_wdata_bits_wdata_42(StreamControllerStore_io_dram_wdata_bits_wdata_42),
    .io_dram_wdata_bits_wdata_43(StreamControllerStore_io_dram_wdata_bits_wdata_43),
    .io_dram_wdata_bits_wdata_44(StreamControllerStore_io_dram_wdata_bits_wdata_44),
    .io_dram_wdata_bits_wdata_45(StreamControllerStore_io_dram_wdata_bits_wdata_45),
    .io_dram_wdata_bits_wdata_46(StreamControllerStore_io_dram_wdata_bits_wdata_46),
    .io_dram_wdata_bits_wdata_47(StreamControllerStore_io_dram_wdata_bits_wdata_47),
    .io_dram_wdata_bits_wdata_48(StreamControllerStore_io_dram_wdata_bits_wdata_48),
    .io_dram_wdata_bits_wdata_49(StreamControllerStore_io_dram_wdata_bits_wdata_49),
    .io_dram_wdata_bits_wdata_50(StreamControllerStore_io_dram_wdata_bits_wdata_50),
    .io_dram_wdata_bits_wdata_51(StreamControllerStore_io_dram_wdata_bits_wdata_51),
    .io_dram_wdata_bits_wdata_52(StreamControllerStore_io_dram_wdata_bits_wdata_52),
    .io_dram_wdata_bits_wdata_53(StreamControllerStore_io_dram_wdata_bits_wdata_53),
    .io_dram_wdata_bits_wdata_54(StreamControllerStore_io_dram_wdata_bits_wdata_54),
    .io_dram_wdata_bits_wdata_55(StreamControllerStore_io_dram_wdata_bits_wdata_55),
    .io_dram_wdata_bits_wdata_56(StreamControllerStore_io_dram_wdata_bits_wdata_56),
    .io_dram_wdata_bits_wdata_57(StreamControllerStore_io_dram_wdata_bits_wdata_57),
    .io_dram_wdata_bits_wdata_58(StreamControllerStore_io_dram_wdata_bits_wdata_58),
    .io_dram_wdata_bits_wdata_59(StreamControllerStore_io_dram_wdata_bits_wdata_59),
    .io_dram_wdata_bits_wdata_60(StreamControllerStore_io_dram_wdata_bits_wdata_60),
    .io_dram_wdata_bits_wdata_61(StreamControllerStore_io_dram_wdata_bits_wdata_61),
    .io_dram_wdata_bits_wdata_62(StreamControllerStore_io_dram_wdata_bits_wdata_62),
    .io_dram_wdata_bits_wdata_63(StreamControllerStore_io_dram_wdata_bits_wdata_63),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@106837.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_rresp_valid(StreamArbiter_io_app_0_rresp_valid),
    .io_app_0_rresp_bits_rdata_0(StreamArbiter_io_app_0_rresp_bits_rdata_0),
    .io_app_0_rresp_bits_rdata_1(StreamArbiter_io_app_0_rresp_bits_rdata_1),
    .io_app_0_rresp_bits_rdata_2(StreamArbiter_io_app_0_rresp_bits_rdata_2),
    .io_app_0_rresp_bits_rdata_3(StreamArbiter_io_app_0_rresp_bits_rdata_3),
    .io_app_0_rresp_bits_rdata_4(StreamArbiter_io_app_0_rresp_bits_rdata_4),
    .io_app_0_rresp_bits_rdata_5(StreamArbiter_io_app_0_rresp_bits_rdata_5),
    .io_app_0_rresp_bits_rdata_6(StreamArbiter_io_app_0_rresp_bits_rdata_6),
    .io_app_0_rresp_bits_rdata_7(StreamArbiter_io_app_0_rresp_bits_rdata_7),
    .io_app_0_rresp_bits_rdata_8(StreamArbiter_io_app_0_rresp_bits_rdata_8),
    .io_app_0_rresp_bits_rdata_9(StreamArbiter_io_app_0_rresp_bits_rdata_9),
    .io_app_0_rresp_bits_rdata_10(StreamArbiter_io_app_0_rresp_bits_rdata_10),
    .io_app_0_rresp_bits_rdata_11(StreamArbiter_io_app_0_rresp_bits_rdata_11),
    .io_app_0_rresp_bits_rdata_12(StreamArbiter_io_app_0_rresp_bits_rdata_12),
    .io_app_0_rresp_bits_rdata_13(StreamArbiter_io_app_0_rresp_bits_rdata_13),
    .io_app_0_rresp_bits_rdata_14(StreamArbiter_io_app_0_rresp_bits_rdata_14),
    .io_app_0_rresp_bits_rdata_15(StreamArbiter_io_app_0_rresp_bits_rdata_15),
    .io_app_0_rresp_bits_rdata_16(StreamArbiter_io_app_0_rresp_bits_rdata_16),
    .io_app_0_rresp_bits_rdata_17(StreamArbiter_io_app_0_rresp_bits_rdata_17),
    .io_app_0_rresp_bits_rdata_18(StreamArbiter_io_app_0_rresp_bits_rdata_18),
    .io_app_0_rresp_bits_rdata_19(StreamArbiter_io_app_0_rresp_bits_rdata_19),
    .io_app_0_rresp_bits_rdata_20(StreamArbiter_io_app_0_rresp_bits_rdata_20),
    .io_app_0_rresp_bits_rdata_21(StreamArbiter_io_app_0_rresp_bits_rdata_21),
    .io_app_0_rresp_bits_rdata_22(StreamArbiter_io_app_0_rresp_bits_rdata_22),
    .io_app_0_rresp_bits_rdata_23(StreamArbiter_io_app_0_rresp_bits_rdata_23),
    .io_app_0_rresp_bits_rdata_24(StreamArbiter_io_app_0_rresp_bits_rdata_24),
    .io_app_0_rresp_bits_rdata_25(StreamArbiter_io_app_0_rresp_bits_rdata_25),
    .io_app_0_rresp_bits_rdata_26(StreamArbiter_io_app_0_rresp_bits_rdata_26),
    .io_app_0_rresp_bits_rdata_27(StreamArbiter_io_app_0_rresp_bits_rdata_27),
    .io_app_0_rresp_bits_rdata_28(StreamArbiter_io_app_0_rresp_bits_rdata_28),
    .io_app_0_rresp_bits_rdata_29(StreamArbiter_io_app_0_rresp_bits_rdata_29),
    .io_app_0_rresp_bits_rdata_30(StreamArbiter_io_app_0_rresp_bits_rdata_30),
    .io_app_0_rresp_bits_rdata_31(StreamArbiter_io_app_0_rresp_bits_rdata_31),
    .io_app_0_rresp_bits_rdata_32(StreamArbiter_io_app_0_rresp_bits_rdata_32),
    .io_app_0_rresp_bits_rdata_33(StreamArbiter_io_app_0_rresp_bits_rdata_33),
    .io_app_0_rresp_bits_rdata_34(StreamArbiter_io_app_0_rresp_bits_rdata_34),
    .io_app_0_rresp_bits_rdata_35(StreamArbiter_io_app_0_rresp_bits_rdata_35),
    .io_app_0_rresp_bits_rdata_36(StreamArbiter_io_app_0_rresp_bits_rdata_36),
    .io_app_0_rresp_bits_rdata_37(StreamArbiter_io_app_0_rresp_bits_rdata_37),
    .io_app_0_rresp_bits_rdata_38(StreamArbiter_io_app_0_rresp_bits_rdata_38),
    .io_app_0_rresp_bits_rdata_39(StreamArbiter_io_app_0_rresp_bits_rdata_39),
    .io_app_0_rresp_bits_rdata_40(StreamArbiter_io_app_0_rresp_bits_rdata_40),
    .io_app_0_rresp_bits_rdata_41(StreamArbiter_io_app_0_rresp_bits_rdata_41),
    .io_app_0_rresp_bits_rdata_42(StreamArbiter_io_app_0_rresp_bits_rdata_42),
    .io_app_0_rresp_bits_rdata_43(StreamArbiter_io_app_0_rresp_bits_rdata_43),
    .io_app_0_rresp_bits_rdata_44(StreamArbiter_io_app_0_rresp_bits_rdata_44),
    .io_app_0_rresp_bits_rdata_45(StreamArbiter_io_app_0_rresp_bits_rdata_45),
    .io_app_0_rresp_bits_rdata_46(StreamArbiter_io_app_0_rresp_bits_rdata_46),
    .io_app_0_rresp_bits_rdata_47(StreamArbiter_io_app_0_rresp_bits_rdata_47),
    .io_app_0_rresp_bits_rdata_48(StreamArbiter_io_app_0_rresp_bits_rdata_48),
    .io_app_0_rresp_bits_rdata_49(StreamArbiter_io_app_0_rresp_bits_rdata_49),
    .io_app_0_rresp_bits_rdata_50(StreamArbiter_io_app_0_rresp_bits_rdata_50),
    .io_app_0_rresp_bits_rdata_51(StreamArbiter_io_app_0_rresp_bits_rdata_51),
    .io_app_0_rresp_bits_rdata_52(StreamArbiter_io_app_0_rresp_bits_rdata_52),
    .io_app_0_rresp_bits_rdata_53(StreamArbiter_io_app_0_rresp_bits_rdata_53),
    .io_app_0_rresp_bits_rdata_54(StreamArbiter_io_app_0_rresp_bits_rdata_54),
    .io_app_0_rresp_bits_rdata_55(StreamArbiter_io_app_0_rresp_bits_rdata_55),
    .io_app_0_rresp_bits_rdata_56(StreamArbiter_io_app_0_rresp_bits_rdata_56),
    .io_app_0_rresp_bits_rdata_57(StreamArbiter_io_app_0_rresp_bits_rdata_57),
    .io_app_0_rresp_bits_rdata_58(StreamArbiter_io_app_0_rresp_bits_rdata_58),
    .io_app_0_rresp_bits_rdata_59(StreamArbiter_io_app_0_rresp_bits_rdata_59),
    .io_app_0_rresp_bits_rdata_60(StreamArbiter_io_app_0_rresp_bits_rdata_60),
    .io_app_0_rresp_bits_rdata_61(StreamArbiter_io_app_0_rresp_bits_rdata_61),
    .io_app_0_rresp_bits_rdata_62(StreamArbiter_io_app_0_rresp_bits_rdata_62),
    .io_app_0_rresp_bits_rdata_63(StreamArbiter_io_app_0_rresp_bits_rdata_63),
    .io_app_1_cmd_ready(StreamArbiter_io_app_1_cmd_ready),
    .io_app_1_cmd_valid(StreamArbiter_io_app_1_cmd_valid),
    .io_app_1_cmd_bits_addr(StreamArbiter_io_app_1_cmd_bits_addr),
    .io_app_1_cmd_bits_size(StreamArbiter_io_app_1_cmd_bits_size),
    .io_app_1_wdata_ready(StreamArbiter_io_app_1_wdata_ready),
    .io_app_1_wdata_valid(StreamArbiter_io_app_1_wdata_valid),
    .io_app_1_wdata_bits_wdata_0(StreamArbiter_io_app_1_wdata_bits_wdata_0),
    .io_app_1_wdata_bits_wdata_1(StreamArbiter_io_app_1_wdata_bits_wdata_1),
    .io_app_1_wdata_bits_wdata_2(StreamArbiter_io_app_1_wdata_bits_wdata_2),
    .io_app_1_wdata_bits_wdata_3(StreamArbiter_io_app_1_wdata_bits_wdata_3),
    .io_app_1_wdata_bits_wdata_4(StreamArbiter_io_app_1_wdata_bits_wdata_4),
    .io_app_1_wdata_bits_wdata_5(StreamArbiter_io_app_1_wdata_bits_wdata_5),
    .io_app_1_wdata_bits_wdata_6(StreamArbiter_io_app_1_wdata_bits_wdata_6),
    .io_app_1_wdata_bits_wdata_7(StreamArbiter_io_app_1_wdata_bits_wdata_7),
    .io_app_1_wdata_bits_wdata_8(StreamArbiter_io_app_1_wdata_bits_wdata_8),
    .io_app_1_wdata_bits_wdata_9(StreamArbiter_io_app_1_wdata_bits_wdata_9),
    .io_app_1_wdata_bits_wdata_10(StreamArbiter_io_app_1_wdata_bits_wdata_10),
    .io_app_1_wdata_bits_wdata_11(StreamArbiter_io_app_1_wdata_bits_wdata_11),
    .io_app_1_wdata_bits_wdata_12(StreamArbiter_io_app_1_wdata_bits_wdata_12),
    .io_app_1_wdata_bits_wdata_13(StreamArbiter_io_app_1_wdata_bits_wdata_13),
    .io_app_1_wdata_bits_wdata_14(StreamArbiter_io_app_1_wdata_bits_wdata_14),
    .io_app_1_wdata_bits_wdata_15(StreamArbiter_io_app_1_wdata_bits_wdata_15),
    .io_app_1_wdata_bits_wdata_16(StreamArbiter_io_app_1_wdata_bits_wdata_16),
    .io_app_1_wdata_bits_wdata_17(StreamArbiter_io_app_1_wdata_bits_wdata_17),
    .io_app_1_wdata_bits_wdata_18(StreamArbiter_io_app_1_wdata_bits_wdata_18),
    .io_app_1_wdata_bits_wdata_19(StreamArbiter_io_app_1_wdata_bits_wdata_19),
    .io_app_1_wdata_bits_wdata_20(StreamArbiter_io_app_1_wdata_bits_wdata_20),
    .io_app_1_wdata_bits_wdata_21(StreamArbiter_io_app_1_wdata_bits_wdata_21),
    .io_app_1_wdata_bits_wdata_22(StreamArbiter_io_app_1_wdata_bits_wdata_22),
    .io_app_1_wdata_bits_wdata_23(StreamArbiter_io_app_1_wdata_bits_wdata_23),
    .io_app_1_wdata_bits_wdata_24(StreamArbiter_io_app_1_wdata_bits_wdata_24),
    .io_app_1_wdata_bits_wdata_25(StreamArbiter_io_app_1_wdata_bits_wdata_25),
    .io_app_1_wdata_bits_wdata_26(StreamArbiter_io_app_1_wdata_bits_wdata_26),
    .io_app_1_wdata_bits_wdata_27(StreamArbiter_io_app_1_wdata_bits_wdata_27),
    .io_app_1_wdata_bits_wdata_28(StreamArbiter_io_app_1_wdata_bits_wdata_28),
    .io_app_1_wdata_bits_wdata_29(StreamArbiter_io_app_1_wdata_bits_wdata_29),
    .io_app_1_wdata_bits_wdata_30(StreamArbiter_io_app_1_wdata_bits_wdata_30),
    .io_app_1_wdata_bits_wdata_31(StreamArbiter_io_app_1_wdata_bits_wdata_31),
    .io_app_1_wdata_bits_wdata_32(StreamArbiter_io_app_1_wdata_bits_wdata_32),
    .io_app_1_wdata_bits_wdata_33(StreamArbiter_io_app_1_wdata_bits_wdata_33),
    .io_app_1_wdata_bits_wdata_34(StreamArbiter_io_app_1_wdata_bits_wdata_34),
    .io_app_1_wdata_bits_wdata_35(StreamArbiter_io_app_1_wdata_bits_wdata_35),
    .io_app_1_wdata_bits_wdata_36(StreamArbiter_io_app_1_wdata_bits_wdata_36),
    .io_app_1_wdata_bits_wdata_37(StreamArbiter_io_app_1_wdata_bits_wdata_37),
    .io_app_1_wdata_bits_wdata_38(StreamArbiter_io_app_1_wdata_bits_wdata_38),
    .io_app_1_wdata_bits_wdata_39(StreamArbiter_io_app_1_wdata_bits_wdata_39),
    .io_app_1_wdata_bits_wdata_40(StreamArbiter_io_app_1_wdata_bits_wdata_40),
    .io_app_1_wdata_bits_wdata_41(StreamArbiter_io_app_1_wdata_bits_wdata_41),
    .io_app_1_wdata_bits_wdata_42(StreamArbiter_io_app_1_wdata_bits_wdata_42),
    .io_app_1_wdata_bits_wdata_43(StreamArbiter_io_app_1_wdata_bits_wdata_43),
    .io_app_1_wdata_bits_wdata_44(StreamArbiter_io_app_1_wdata_bits_wdata_44),
    .io_app_1_wdata_bits_wdata_45(StreamArbiter_io_app_1_wdata_bits_wdata_45),
    .io_app_1_wdata_bits_wdata_46(StreamArbiter_io_app_1_wdata_bits_wdata_46),
    .io_app_1_wdata_bits_wdata_47(StreamArbiter_io_app_1_wdata_bits_wdata_47),
    .io_app_1_wdata_bits_wdata_48(StreamArbiter_io_app_1_wdata_bits_wdata_48),
    .io_app_1_wdata_bits_wdata_49(StreamArbiter_io_app_1_wdata_bits_wdata_49),
    .io_app_1_wdata_bits_wdata_50(StreamArbiter_io_app_1_wdata_bits_wdata_50),
    .io_app_1_wdata_bits_wdata_51(StreamArbiter_io_app_1_wdata_bits_wdata_51),
    .io_app_1_wdata_bits_wdata_52(StreamArbiter_io_app_1_wdata_bits_wdata_52),
    .io_app_1_wdata_bits_wdata_53(StreamArbiter_io_app_1_wdata_bits_wdata_53),
    .io_app_1_wdata_bits_wdata_54(StreamArbiter_io_app_1_wdata_bits_wdata_54),
    .io_app_1_wdata_bits_wdata_55(StreamArbiter_io_app_1_wdata_bits_wdata_55),
    .io_app_1_wdata_bits_wdata_56(StreamArbiter_io_app_1_wdata_bits_wdata_56),
    .io_app_1_wdata_bits_wdata_57(StreamArbiter_io_app_1_wdata_bits_wdata_57),
    .io_app_1_wdata_bits_wdata_58(StreamArbiter_io_app_1_wdata_bits_wdata_58),
    .io_app_1_wdata_bits_wdata_59(StreamArbiter_io_app_1_wdata_bits_wdata_59),
    .io_app_1_wdata_bits_wdata_60(StreamArbiter_io_app_1_wdata_bits_wdata_60),
    .io_app_1_wdata_bits_wdata_61(StreamArbiter_io_app_1_wdata_bits_wdata_61),
    .io_app_1_wdata_bits_wdata_62(StreamArbiter_io_app_1_wdata_bits_wdata_62),
    .io_app_1_wdata_bits_wdata_63(StreamArbiter_io_app_1_wdata_bits_wdata_63),
    .io_app_1_wdata_bits_wstrb_0(StreamArbiter_io_app_1_wdata_bits_wstrb_0),
    .io_app_1_wdata_bits_wstrb_1(StreamArbiter_io_app_1_wdata_bits_wstrb_1),
    .io_app_1_wdata_bits_wstrb_2(StreamArbiter_io_app_1_wdata_bits_wstrb_2),
    .io_app_1_wdata_bits_wstrb_3(StreamArbiter_io_app_1_wdata_bits_wstrb_3),
    .io_app_1_wdata_bits_wstrb_4(StreamArbiter_io_app_1_wdata_bits_wstrb_4),
    .io_app_1_wdata_bits_wstrb_5(StreamArbiter_io_app_1_wdata_bits_wstrb_5),
    .io_app_1_wdata_bits_wstrb_6(StreamArbiter_io_app_1_wdata_bits_wstrb_6),
    .io_app_1_wdata_bits_wstrb_7(StreamArbiter_io_app_1_wdata_bits_wstrb_7),
    .io_app_1_wdata_bits_wstrb_8(StreamArbiter_io_app_1_wdata_bits_wstrb_8),
    .io_app_1_wdata_bits_wstrb_9(StreamArbiter_io_app_1_wdata_bits_wstrb_9),
    .io_app_1_wdata_bits_wstrb_10(StreamArbiter_io_app_1_wdata_bits_wstrb_10),
    .io_app_1_wdata_bits_wstrb_11(StreamArbiter_io_app_1_wdata_bits_wstrb_11),
    .io_app_1_wdata_bits_wstrb_12(StreamArbiter_io_app_1_wdata_bits_wstrb_12),
    .io_app_1_wdata_bits_wstrb_13(StreamArbiter_io_app_1_wdata_bits_wstrb_13),
    .io_app_1_wdata_bits_wstrb_14(StreamArbiter_io_app_1_wdata_bits_wstrb_14),
    .io_app_1_wdata_bits_wstrb_15(StreamArbiter_io_app_1_wdata_bits_wstrb_15),
    .io_app_1_wdata_bits_wstrb_16(StreamArbiter_io_app_1_wdata_bits_wstrb_16),
    .io_app_1_wdata_bits_wstrb_17(StreamArbiter_io_app_1_wdata_bits_wstrb_17),
    .io_app_1_wdata_bits_wstrb_18(StreamArbiter_io_app_1_wdata_bits_wstrb_18),
    .io_app_1_wdata_bits_wstrb_19(StreamArbiter_io_app_1_wdata_bits_wstrb_19),
    .io_app_1_wdata_bits_wstrb_20(StreamArbiter_io_app_1_wdata_bits_wstrb_20),
    .io_app_1_wdata_bits_wstrb_21(StreamArbiter_io_app_1_wdata_bits_wstrb_21),
    .io_app_1_wdata_bits_wstrb_22(StreamArbiter_io_app_1_wdata_bits_wstrb_22),
    .io_app_1_wdata_bits_wstrb_23(StreamArbiter_io_app_1_wdata_bits_wstrb_23),
    .io_app_1_wdata_bits_wstrb_24(StreamArbiter_io_app_1_wdata_bits_wstrb_24),
    .io_app_1_wdata_bits_wstrb_25(StreamArbiter_io_app_1_wdata_bits_wstrb_25),
    .io_app_1_wdata_bits_wstrb_26(StreamArbiter_io_app_1_wdata_bits_wstrb_26),
    .io_app_1_wdata_bits_wstrb_27(StreamArbiter_io_app_1_wdata_bits_wstrb_27),
    .io_app_1_wdata_bits_wstrb_28(StreamArbiter_io_app_1_wdata_bits_wstrb_28),
    .io_app_1_wdata_bits_wstrb_29(StreamArbiter_io_app_1_wdata_bits_wstrb_29),
    .io_app_1_wdata_bits_wstrb_30(StreamArbiter_io_app_1_wdata_bits_wstrb_30),
    .io_app_1_wdata_bits_wstrb_31(StreamArbiter_io_app_1_wdata_bits_wstrb_31),
    .io_app_1_wdata_bits_wstrb_32(StreamArbiter_io_app_1_wdata_bits_wstrb_32),
    .io_app_1_wdata_bits_wstrb_33(StreamArbiter_io_app_1_wdata_bits_wstrb_33),
    .io_app_1_wdata_bits_wstrb_34(StreamArbiter_io_app_1_wdata_bits_wstrb_34),
    .io_app_1_wdata_bits_wstrb_35(StreamArbiter_io_app_1_wdata_bits_wstrb_35),
    .io_app_1_wdata_bits_wstrb_36(StreamArbiter_io_app_1_wdata_bits_wstrb_36),
    .io_app_1_wdata_bits_wstrb_37(StreamArbiter_io_app_1_wdata_bits_wstrb_37),
    .io_app_1_wdata_bits_wstrb_38(StreamArbiter_io_app_1_wdata_bits_wstrb_38),
    .io_app_1_wdata_bits_wstrb_39(StreamArbiter_io_app_1_wdata_bits_wstrb_39),
    .io_app_1_wdata_bits_wstrb_40(StreamArbiter_io_app_1_wdata_bits_wstrb_40),
    .io_app_1_wdata_bits_wstrb_41(StreamArbiter_io_app_1_wdata_bits_wstrb_41),
    .io_app_1_wdata_bits_wstrb_42(StreamArbiter_io_app_1_wdata_bits_wstrb_42),
    .io_app_1_wdata_bits_wstrb_43(StreamArbiter_io_app_1_wdata_bits_wstrb_43),
    .io_app_1_wdata_bits_wstrb_44(StreamArbiter_io_app_1_wdata_bits_wstrb_44),
    .io_app_1_wdata_bits_wstrb_45(StreamArbiter_io_app_1_wdata_bits_wstrb_45),
    .io_app_1_wdata_bits_wstrb_46(StreamArbiter_io_app_1_wdata_bits_wstrb_46),
    .io_app_1_wdata_bits_wstrb_47(StreamArbiter_io_app_1_wdata_bits_wstrb_47),
    .io_app_1_wdata_bits_wstrb_48(StreamArbiter_io_app_1_wdata_bits_wstrb_48),
    .io_app_1_wdata_bits_wstrb_49(StreamArbiter_io_app_1_wdata_bits_wstrb_49),
    .io_app_1_wdata_bits_wstrb_50(StreamArbiter_io_app_1_wdata_bits_wstrb_50),
    .io_app_1_wdata_bits_wstrb_51(StreamArbiter_io_app_1_wdata_bits_wstrb_51),
    .io_app_1_wdata_bits_wstrb_52(StreamArbiter_io_app_1_wdata_bits_wstrb_52),
    .io_app_1_wdata_bits_wstrb_53(StreamArbiter_io_app_1_wdata_bits_wstrb_53),
    .io_app_1_wdata_bits_wstrb_54(StreamArbiter_io_app_1_wdata_bits_wstrb_54),
    .io_app_1_wdata_bits_wstrb_55(StreamArbiter_io_app_1_wdata_bits_wstrb_55),
    .io_app_1_wdata_bits_wstrb_56(StreamArbiter_io_app_1_wdata_bits_wstrb_56),
    .io_app_1_wdata_bits_wstrb_57(StreamArbiter_io_app_1_wdata_bits_wstrb_57),
    .io_app_1_wdata_bits_wstrb_58(StreamArbiter_io_app_1_wdata_bits_wstrb_58),
    .io_app_1_wdata_bits_wstrb_59(StreamArbiter_io_app_1_wdata_bits_wstrb_59),
    .io_app_1_wdata_bits_wstrb_60(StreamArbiter_io_app_1_wdata_bits_wstrb_60),
    .io_app_1_wdata_bits_wstrb_61(StreamArbiter_io_app_1_wdata_bits_wstrb_61),
    .io_app_1_wdata_bits_wstrb_62(StreamArbiter_io_app_1_wdata_bits_wstrb_62),
    .io_app_1_wdata_bits_wstrb_63(StreamArbiter_io_app_1_wdata_bits_wstrb_63),
    .io_app_1_wresp_ready(StreamArbiter_io_app_1_wresp_ready),
    .io_app_1_wresp_valid(StreamArbiter_io_app_1_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wdata_16(StreamArbiter_io_dram_wdata_bits_wdata_16),
    .io_dram_wdata_bits_wdata_17(StreamArbiter_io_dram_wdata_bits_wdata_17),
    .io_dram_wdata_bits_wdata_18(StreamArbiter_io_dram_wdata_bits_wdata_18),
    .io_dram_wdata_bits_wdata_19(StreamArbiter_io_dram_wdata_bits_wdata_19),
    .io_dram_wdata_bits_wdata_20(StreamArbiter_io_dram_wdata_bits_wdata_20),
    .io_dram_wdata_bits_wdata_21(StreamArbiter_io_dram_wdata_bits_wdata_21),
    .io_dram_wdata_bits_wdata_22(StreamArbiter_io_dram_wdata_bits_wdata_22),
    .io_dram_wdata_bits_wdata_23(StreamArbiter_io_dram_wdata_bits_wdata_23),
    .io_dram_wdata_bits_wdata_24(StreamArbiter_io_dram_wdata_bits_wdata_24),
    .io_dram_wdata_bits_wdata_25(StreamArbiter_io_dram_wdata_bits_wdata_25),
    .io_dram_wdata_bits_wdata_26(StreamArbiter_io_dram_wdata_bits_wdata_26),
    .io_dram_wdata_bits_wdata_27(StreamArbiter_io_dram_wdata_bits_wdata_27),
    .io_dram_wdata_bits_wdata_28(StreamArbiter_io_dram_wdata_bits_wdata_28),
    .io_dram_wdata_bits_wdata_29(StreamArbiter_io_dram_wdata_bits_wdata_29),
    .io_dram_wdata_bits_wdata_30(StreamArbiter_io_dram_wdata_bits_wdata_30),
    .io_dram_wdata_bits_wdata_31(StreamArbiter_io_dram_wdata_bits_wdata_31),
    .io_dram_wdata_bits_wdata_32(StreamArbiter_io_dram_wdata_bits_wdata_32),
    .io_dram_wdata_bits_wdata_33(StreamArbiter_io_dram_wdata_bits_wdata_33),
    .io_dram_wdata_bits_wdata_34(StreamArbiter_io_dram_wdata_bits_wdata_34),
    .io_dram_wdata_bits_wdata_35(StreamArbiter_io_dram_wdata_bits_wdata_35),
    .io_dram_wdata_bits_wdata_36(StreamArbiter_io_dram_wdata_bits_wdata_36),
    .io_dram_wdata_bits_wdata_37(StreamArbiter_io_dram_wdata_bits_wdata_37),
    .io_dram_wdata_bits_wdata_38(StreamArbiter_io_dram_wdata_bits_wdata_38),
    .io_dram_wdata_bits_wdata_39(StreamArbiter_io_dram_wdata_bits_wdata_39),
    .io_dram_wdata_bits_wdata_40(StreamArbiter_io_dram_wdata_bits_wdata_40),
    .io_dram_wdata_bits_wdata_41(StreamArbiter_io_dram_wdata_bits_wdata_41),
    .io_dram_wdata_bits_wdata_42(StreamArbiter_io_dram_wdata_bits_wdata_42),
    .io_dram_wdata_bits_wdata_43(StreamArbiter_io_dram_wdata_bits_wdata_43),
    .io_dram_wdata_bits_wdata_44(StreamArbiter_io_dram_wdata_bits_wdata_44),
    .io_dram_wdata_bits_wdata_45(StreamArbiter_io_dram_wdata_bits_wdata_45),
    .io_dram_wdata_bits_wdata_46(StreamArbiter_io_dram_wdata_bits_wdata_46),
    .io_dram_wdata_bits_wdata_47(StreamArbiter_io_dram_wdata_bits_wdata_47),
    .io_dram_wdata_bits_wdata_48(StreamArbiter_io_dram_wdata_bits_wdata_48),
    .io_dram_wdata_bits_wdata_49(StreamArbiter_io_dram_wdata_bits_wdata_49),
    .io_dram_wdata_bits_wdata_50(StreamArbiter_io_dram_wdata_bits_wdata_50),
    .io_dram_wdata_bits_wdata_51(StreamArbiter_io_dram_wdata_bits_wdata_51),
    .io_dram_wdata_bits_wdata_52(StreamArbiter_io_dram_wdata_bits_wdata_52),
    .io_dram_wdata_bits_wdata_53(StreamArbiter_io_dram_wdata_bits_wdata_53),
    .io_dram_wdata_bits_wdata_54(StreamArbiter_io_dram_wdata_bits_wdata_54),
    .io_dram_wdata_bits_wdata_55(StreamArbiter_io_dram_wdata_bits_wdata_55),
    .io_dram_wdata_bits_wdata_56(StreamArbiter_io_dram_wdata_bits_wdata_56),
    .io_dram_wdata_bits_wdata_57(StreamArbiter_io_dram_wdata_bits_wdata_57),
    .io_dram_wdata_bits_wdata_58(StreamArbiter_io_dram_wdata_bits_wdata_58),
    .io_dram_wdata_bits_wdata_59(StreamArbiter_io_dram_wdata_bits_wdata_59),
    .io_dram_wdata_bits_wdata_60(StreamArbiter_io_dram_wdata_bits_wdata_60),
    .io_dram_wdata_bits_wdata_61(StreamArbiter_io_dram_wdata_bits_wdata_61),
    .io_dram_wdata_bits_wdata_62(StreamArbiter_io_dram_wdata_bits_wdata_62),
    .io_dram_wdata_bits_wdata_63(StreamArbiter_io_dram_wdata_bits_wdata_63),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_rresp_valid(StreamArbiter_io_dram_rresp_valid),
    .io_dram_rresp_bits_rdata_0(StreamArbiter_io_dram_rresp_bits_rdata_0),
    .io_dram_rresp_bits_rdata_1(StreamArbiter_io_dram_rresp_bits_rdata_1),
    .io_dram_rresp_bits_rdata_2(StreamArbiter_io_dram_rresp_bits_rdata_2),
    .io_dram_rresp_bits_rdata_3(StreamArbiter_io_dram_rresp_bits_rdata_3),
    .io_dram_rresp_bits_rdata_4(StreamArbiter_io_dram_rresp_bits_rdata_4),
    .io_dram_rresp_bits_rdata_5(StreamArbiter_io_dram_rresp_bits_rdata_5),
    .io_dram_rresp_bits_rdata_6(StreamArbiter_io_dram_rresp_bits_rdata_6),
    .io_dram_rresp_bits_rdata_7(StreamArbiter_io_dram_rresp_bits_rdata_7),
    .io_dram_rresp_bits_rdata_8(StreamArbiter_io_dram_rresp_bits_rdata_8),
    .io_dram_rresp_bits_rdata_9(StreamArbiter_io_dram_rresp_bits_rdata_9),
    .io_dram_rresp_bits_rdata_10(StreamArbiter_io_dram_rresp_bits_rdata_10),
    .io_dram_rresp_bits_rdata_11(StreamArbiter_io_dram_rresp_bits_rdata_11),
    .io_dram_rresp_bits_rdata_12(StreamArbiter_io_dram_rresp_bits_rdata_12),
    .io_dram_rresp_bits_rdata_13(StreamArbiter_io_dram_rresp_bits_rdata_13),
    .io_dram_rresp_bits_rdata_14(StreamArbiter_io_dram_rresp_bits_rdata_14),
    .io_dram_rresp_bits_rdata_15(StreamArbiter_io_dram_rresp_bits_rdata_15),
    .io_dram_rresp_bits_rdata_16(StreamArbiter_io_dram_rresp_bits_rdata_16),
    .io_dram_rresp_bits_rdata_17(StreamArbiter_io_dram_rresp_bits_rdata_17),
    .io_dram_rresp_bits_rdata_18(StreamArbiter_io_dram_rresp_bits_rdata_18),
    .io_dram_rresp_bits_rdata_19(StreamArbiter_io_dram_rresp_bits_rdata_19),
    .io_dram_rresp_bits_rdata_20(StreamArbiter_io_dram_rresp_bits_rdata_20),
    .io_dram_rresp_bits_rdata_21(StreamArbiter_io_dram_rresp_bits_rdata_21),
    .io_dram_rresp_bits_rdata_22(StreamArbiter_io_dram_rresp_bits_rdata_22),
    .io_dram_rresp_bits_rdata_23(StreamArbiter_io_dram_rresp_bits_rdata_23),
    .io_dram_rresp_bits_rdata_24(StreamArbiter_io_dram_rresp_bits_rdata_24),
    .io_dram_rresp_bits_rdata_25(StreamArbiter_io_dram_rresp_bits_rdata_25),
    .io_dram_rresp_bits_rdata_26(StreamArbiter_io_dram_rresp_bits_rdata_26),
    .io_dram_rresp_bits_rdata_27(StreamArbiter_io_dram_rresp_bits_rdata_27),
    .io_dram_rresp_bits_rdata_28(StreamArbiter_io_dram_rresp_bits_rdata_28),
    .io_dram_rresp_bits_rdata_29(StreamArbiter_io_dram_rresp_bits_rdata_29),
    .io_dram_rresp_bits_rdata_30(StreamArbiter_io_dram_rresp_bits_rdata_30),
    .io_dram_rresp_bits_rdata_31(StreamArbiter_io_dram_rresp_bits_rdata_31),
    .io_dram_rresp_bits_rdata_32(StreamArbiter_io_dram_rresp_bits_rdata_32),
    .io_dram_rresp_bits_rdata_33(StreamArbiter_io_dram_rresp_bits_rdata_33),
    .io_dram_rresp_bits_rdata_34(StreamArbiter_io_dram_rresp_bits_rdata_34),
    .io_dram_rresp_bits_rdata_35(StreamArbiter_io_dram_rresp_bits_rdata_35),
    .io_dram_rresp_bits_rdata_36(StreamArbiter_io_dram_rresp_bits_rdata_36),
    .io_dram_rresp_bits_rdata_37(StreamArbiter_io_dram_rresp_bits_rdata_37),
    .io_dram_rresp_bits_rdata_38(StreamArbiter_io_dram_rresp_bits_rdata_38),
    .io_dram_rresp_bits_rdata_39(StreamArbiter_io_dram_rresp_bits_rdata_39),
    .io_dram_rresp_bits_rdata_40(StreamArbiter_io_dram_rresp_bits_rdata_40),
    .io_dram_rresp_bits_rdata_41(StreamArbiter_io_dram_rresp_bits_rdata_41),
    .io_dram_rresp_bits_rdata_42(StreamArbiter_io_dram_rresp_bits_rdata_42),
    .io_dram_rresp_bits_rdata_43(StreamArbiter_io_dram_rresp_bits_rdata_43),
    .io_dram_rresp_bits_rdata_44(StreamArbiter_io_dram_rresp_bits_rdata_44),
    .io_dram_rresp_bits_rdata_45(StreamArbiter_io_dram_rresp_bits_rdata_45),
    .io_dram_rresp_bits_rdata_46(StreamArbiter_io_dram_rresp_bits_rdata_46),
    .io_dram_rresp_bits_rdata_47(StreamArbiter_io_dram_rresp_bits_rdata_47),
    .io_dram_rresp_bits_rdata_48(StreamArbiter_io_dram_rresp_bits_rdata_48),
    .io_dram_rresp_bits_rdata_49(StreamArbiter_io_dram_rresp_bits_rdata_49),
    .io_dram_rresp_bits_rdata_50(StreamArbiter_io_dram_rresp_bits_rdata_50),
    .io_dram_rresp_bits_rdata_51(StreamArbiter_io_dram_rresp_bits_rdata_51),
    .io_dram_rresp_bits_rdata_52(StreamArbiter_io_dram_rresp_bits_rdata_52),
    .io_dram_rresp_bits_rdata_53(StreamArbiter_io_dram_rresp_bits_rdata_53),
    .io_dram_rresp_bits_rdata_54(StreamArbiter_io_dram_rresp_bits_rdata_54),
    .io_dram_rresp_bits_rdata_55(StreamArbiter_io_dram_rresp_bits_rdata_55),
    .io_dram_rresp_bits_rdata_56(StreamArbiter_io_dram_rresp_bits_rdata_56),
    .io_dram_rresp_bits_rdata_57(StreamArbiter_io_dram_rresp_bits_rdata_57),
    .io_dram_rresp_bits_rdata_58(StreamArbiter_io_dram_rresp_bits_rdata_58),
    .io_dram_rresp_bits_rdata_59(StreamArbiter_io_dram_rresp_bits_rdata_59),
    .io_dram_rresp_bits_rdata_60(StreamArbiter_io_dram_rresp_bits_rdata_60),
    .io_dram_rresp_bits_rdata_61(StreamArbiter_io_dram_rresp_bits_rdata_61),
    .io_dram_rresp_bits_rdata_62(StreamArbiter_io_dram_rresp_bits_rdata_62),
    .io_dram_rresp_bits_rdata_63(StreamArbiter_io_dram_rresp_bits_rdata_63),
    .io_dram_rresp_bits_tag(StreamArbiter_io_dram_rresp_bits_tag),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@107673.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wdata_16(AXICmdSplit_io_in_wdata_bits_wdata_16),
    .io_in_wdata_bits_wdata_17(AXICmdSplit_io_in_wdata_bits_wdata_17),
    .io_in_wdata_bits_wdata_18(AXICmdSplit_io_in_wdata_bits_wdata_18),
    .io_in_wdata_bits_wdata_19(AXICmdSplit_io_in_wdata_bits_wdata_19),
    .io_in_wdata_bits_wdata_20(AXICmdSplit_io_in_wdata_bits_wdata_20),
    .io_in_wdata_bits_wdata_21(AXICmdSplit_io_in_wdata_bits_wdata_21),
    .io_in_wdata_bits_wdata_22(AXICmdSplit_io_in_wdata_bits_wdata_22),
    .io_in_wdata_bits_wdata_23(AXICmdSplit_io_in_wdata_bits_wdata_23),
    .io_in_wdata_bits_wdata_24(AXICmdSplit_io_in_wdata_bits_wdata_24),
    .io_in_wdata_bits_wdata_25(AXICmdSplit_io_in_wdata_bits_wdata_25),
    .io_in_wdata_bits_wdata_26(AXICmdSplit_io_in_wdata_bits_wdata_26),
    .io_in_wdata_bits_wdata_27(AXICmdSplit_io_in_wdata_bits_wdata_27),
    .io_in_wdata_bits_wdata_28(AXICmdSplit_io_in_wdata_bits_wdata_28),
    .io_in_wdata_bits_wdata_29(AXICmdSplit_io_in_wdata_bits_wdata_29),
    .io_in_wdata_bits_wdata_30(AXICmdSplit_io_in_wdata_bits_wdata_30),
    .io_in_wdata_bits_wdata_31(AXICmdSplit_io_in_wdata_bits_wdata_31),
    .io_in_wdata_bits_wdata_32(AXICmdSplit_io_in_wdata_bits_wdata_32),
    .io_in_wdata_bits_wdata_33(AXICmdSplit_io_in_wdata_bits_wdata_33),
    .io_in_wdata_bits_wdata_34(AXICmdSplit_io_in_wdata_bits_wdata_34),
    .io_in_wdata_bits_wdata_35(AXICmdSplit_io_in_wdata_bits_wdata_35),
    .io_in_wdata_bits_wdata_36(AXICmdSplit_io_in_wdata_bits_wdata_36),
    .io_in_wdata_bits_wdata_37(AXICmdSplit_io_in_wdata_bits_wdata_37),
    .io_in_wdata_bits_wdata_38(AXICmdSplit_io_in_wdata_bits_wdata_38),
    .io_in_wdata_bits_wdata_39(AXICmdSplit_io_in_wdata_bits_wdata_39),
    .io_in_wdata_bits_wdata_40(AXICmdSplit_io_in_wdata_bits_wdata_40),
    .io_in_wdata_bits_wdata_41(AXICmdSplit_io_in_wdata_bits_wdata_41),
    .io_in_wdata_bits_wdata_42(AXICmdSplit_io_in_wdata_bits_wdata_42),
    .io_in_wdata_bits_wdata_43(AXICmdSplit_io_in_wdata_bits_wdata_43),
    .io_in_wdata_bits_wdata_44(AXICmdSplit_io_in_wdata_bits_wdata_44),
    .io_in_wdata_bits_wdata_45(AXICmdSplit_io_in_wdata_bits_wdata_45),
    .io_in_wdata_bits_wdata_46(AXICmdSplit_io_in_wdata_bits_wdata_46),
    .io_in_wdata_bits_wdata_47(AXICmdSplit_io_in_wdata_bits_wdata_47),
    .io_in_wdata_bits_wdata_48(AXICmdSplit_io_in_wdata_bits_wdata_48),
    .io_in_wdata_bits_wdata_49(AXICmdSplit_io_in_wdata_bits_wdata_49),
    .io_in_wdata_bits_wdata_50(AXICmdSplit_io_in_wdata_bits_wdata_50),
    .io_in_wdata_bits_wdata_51(AXICmdSplit_io_in_wdata_bits_wdata_51),
    .io_in_wdata_bits_wdata_52(AXICmdSplit_io_in_wdata_bits_wdata_52),
    .io_in_wdata_bits_wdata_53(AXICmdSplit_io_in_wdata_bits_wdata_53),
    .io_in_wdata_bits_wdata_54(AXICmdSplit_io_in_wdata_bits_wdata_54),
    .io_in_wdata_bits_wdata_55(AXICmdSplit_io_in_wdata_bits_wdata_55),
    .io_in_wdata_bits_wdata_56(AXICmdSplit_io_in_wdata_bits_wdata_56),
    .io_in_wdata_bits_wdata_57(AXICmdSplit_io_in_wdata_bits_wdata_57),
    .io_in_wdata_bits_wdata_58(AXICmdSplit_io_in_wdata_bits_wdata_58),
    .io_in_wdata_bits_wdata_59(AXICmdSplit_io_in_wdata_bits_wdata_59),
    .io_in_wdata_bits_wdata_60(AXICmdSplit_io_in_wdata_bits_wdata_60),
    .io_in_wdata_bits_wdata_61(AXICmdSplit_io_in_wdata_bits_wdata_61),
    .io_in_wdata_bits_wdata_62(AXICmdSplit_io_in_wdata_bits_wdata_62),
    .io_in_wdata_bits_wdata_63(AXICmdSplit_io_in_wdata_bits_wdata_63),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_rresp_valid(AXICmdSplit_io_in_rresp_valid),
    .io_in_rresp_bits_rdata_0(AXICmdSplit_io_in_rresp_bits_rdata_0),
    .io_in_rresp_bits_rdata_1(AXICmdSplit_io_in_rresp_bits_rdata_1),
    .io_in_rresp_bits_rdata_2(AXICmdSplit_io_in_rresp_bits_rdata_2),
    .io_in_rresp_bits_rdata_3(AXICmdSplit_io_in_rresp_bits_rdata_3),
    .io_in_rresp_bits_rdata_4(AXICmdSplit_io_in_rresp_bits_rdata_4),
    .io_in_rresp_bits_rdata_5(AXICmdSplit_io_in_rresp_bits_rdata_5),
    .io_in_rresp_bits_rdata_6(AXICmdSplit_io_in_rresp_bits_rdata_6),
    .io_in_rresp_bits_rdata_7(AXICmdSplit_io_in_rresp_bits_rdata_7),
    .io_in_rresp_bits_rdata_8(AXICmdSplit_io_in_rresp_bits_rdata_8),
    .io_in_rresp_bits_rdata_9(AXICmdSplit_io_in_rresp_bits_rdata_9),
    .io_in_rresp_bits_rdata_10(AXICmdSplit_io_in_rresp_bits_rdata_10),
    .io_in_rresp_bits_rdata_11(AXICmdSplit_io_in_rresp_bits_rdata_11),
    .io_in_rresp_bits_rdata_12(AXICmdSplit_io_in_rresp_bits_rdata_12),
    .io_in_rresp_bits_rdata_13(AXICmdSplit_io_in_rresp_bits_rdata_13),
    .io_in_rresp_bits_rdata_14(AXICmdSplit_io_in_rresp_bits_rdata_14),
    .io_in_rresp_bits_rdata_15(AXICmdSplit_io_in_rresp_bits_rdata_15),
    .io_in_rresp_bits_rdata_16(AXICmdSplit_io_in_rresp_bits_rdata_16),
    .io_in_rresp_bits_rdata_17(AXICmdSplit_io_in_rresp_bits_rdata_17),
    .io_in_rresp_bits_rdata_18(AXICmdSplit_io_in_rresp_bits_rdata_18),
    .io_in_rresp_bits_rdata_19(AXICmdSplit_io_in_rresp_bits_rdata_19),
    .io_in_rresp_bits_rdata_20(AXICmdSplit_io_in_rresp_bits_rdata_20),
    .io_in_rresp_bits_rdata_21(AXICmdSplit_io_in_rresp_bits_rdata_21),
    .io_in_rresp_bits_rdata_22(AXICmdSplit_io_in_rresp_bits_rdata_22),
    .io_in_rresp_bits_rdata_23(AXICmdSplit_io_in_rresp_bits_rdata_23),
    .io_in_rresp_bits_rdata_24(AXICmdSplit_io_in_rresp_bits_rdata_24),
    .io_in_rresp_bits_rdata_25(AXICmdSplit_io_in_rresp_bits_rdata_25),
    .io_in_rresp_bits_rdata_26(AXICmdSplit_io_in_rresp_bits_rdata_26),
    .io_in_rresp_bits_rdata_27(AXICmdSplit_io_in_rresp_bits_rdata_27),
    .io_in_rresp_bits_rdata_28(AXICmdSplit_io_in_rresp_bits_rdata_28),
    .io_in_rresp_bits_rdata_29(AXICmdSplit_io_in_rresp_bits_rdata_29),
    .io_in_rresp_bits_rdata_30(AXICmdSplit_io_in_rresp_bits_rdata_30),
    .io_in_rresp_bits_rdata_31(AXICmdSplit_io_in_rresp_bits_rdata_31),
    .io_in_rresp_bits_rdata_32(AXICmdSplit_io_in_rresp_bits_rdata_32),
    .io_in_rresp_bits_rdata_33(AXICmdSplit_io_in_rresp_bits_rdata_33),
    .io_in_rresp_bits_rdata_34(AXICmdSplit_io_in_rresp_bits_rdata_34),
    .io_in_rresp_bits_rdata_35(AXICmdSplit_io_in_rresp_bits_rdata_35),
    .io_in_rresp_bits_rdata_36(AXICmdSplit_io_in_rresp_bits_rdata_36),
    .io_in_rresp_bits_rdata_37(AXICmdSplit_io_in_rresp_bits_rdata_37),
    .io_in_rresp_bits_rdata_38(AXICmdSplit_io_in_rresp_bits_rdata_38),
    .io_in_rresp_bits_rdata_39(AXICmdSplit_io_in_rresp_bits_rdata_39),
    .io_in_rresp_bits_rdata_40(AXICmdSplit_io_in_rresp_bits_rdata_40),
    .io_in_rresp_bits_rdata_41(AXICmdSplit_io_in_rresp_bits_rdata_41),
    .io_in_rresp_bits_rdata_42(AXICmdSplit_io_in_rresp_bits_rdata_42),
    .io_in_rresp_bits_rdata_43(AXICmdSplit_io_in_rresp_bits_rdata_43),
    .io_in_rresp_bits_rdata_44(AXICmdSplit_io_in_rresp_bits_rdata_44),
    .io_in_rresp_bits_rdata_45(AXICmdSplit_io_in_rresp_bits_rdata_45),
    .io_in_rresp_bits_rdata_46(AXICmdSplit_io_in_rresp_bits_rdata_46),
    .io_in_rresp_bits_rdata_47(AXICmdSplit_io_in_rresp_bits_rdata_47),
    .io_in_rresp_bits_rdata_48(AXICmdSplit_io_in_rresp_bits_rdata_48),
    .io_in_rresp_bits_rdata_49(AXICmdSplit_io_in_rresp_bits_rdata_49),
    .io_in_rresp_bits_rdata_50(AXICmdSplit_io_in_rresp_bits_rdata_50),
    .io_in_rresp_bits_rdata_51(AXICmdSplit_io_in_rresp_bits_rdata_51),
    .io_in_rresp_bits_rdata_52(AXICmdSplit_io_in_rresp_bits_rdata_52),
    .io_in_rresp_bits_rdata_53(AXICmdSplit_io_in_rresp_bits_rdata_53),
    .io_in_rresp_bits_rdata_54(AXICmdSplit_io_in_rresp_bits_rdata_54),
    .io_in_rresp_bits_rdata_55(AXICmdSplit_io_in_rresp_bits_rdata_55),
    .io_in_rresp_bits_rdata_56(AXICmdSplit_io_in_rresp_bits_rdata_56),
    .io_in_rresp_bits_rdata_57(AXICmdSplit_io_in_rresp_bits_rdata_57),
    .io_in_rresp_bits_rdata_58(AXICmdSplit_io_in_rresp_bits_rdata_58),
    .io_in_rresp_bits_rdata_59(AXICmdSplit_io_in_rresp_bits_rdata_59),
    .io_in_rresp_bits_rdata_60(AXICmdSplit_io_in_rresp_bits_rdata_60),
    .io_in_rresp_bits_rdata_61(AXICmdSplit_io_in_rresp_bits_rdata_61),
    .io_in_rresp_bits_rdata_62(AXICmdSplit_io_in_rresp_bits_rdata_62),
    .io_in_rresp_bits_rdata_63(AXICmdSplit_io_in_rresp_bits_rdata_63),
    .io_in_rresp_bits_tag(AXICmdSplit_io_in_rresp_bits_tag),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_rawAddr(AXICmdSplit_io_out_cmd_bits_rawAddr),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wdata_16(AXICmdSplit_io_out_wdata_bits_wdata_16),
    .io_out_wdata_bits_wdata_17(AXICmdSplit_io_out_wdata_bits_wdata_17),
    .io_out_wdata_bits_wdata_18(AXICmdSplit_io_out_wdata_bits_wdata_18),
    .io_out_wdata_bits_wdata_19(AXICmdSplit_io_out_wdata_bits_wdata_19),
    .io_out_wdata_bits_wdata_20(AXICmdSplit_io_out_wdata_bits_wdata_20),
    .io_out_wdata_bits_wdata_21(AXICmdSplit_io_out_wdata_bits_wdata_21),
    .io_out_wdata_bits_wdata_22(AXICmdSplit_io_out_wdata_bits_wdata_22),
    .io_out_wdata_bits_wdata_23(AXICmdSplit_io_out_wdata_bits_wdata_23),
    .io_out_wdata_bits_wdata_24(AXICmdSplit_io_out_wdata_bits_wdata_24),
    .io_out_wdata_bits_wdata_25(AXICmdSplit_io_out_wdata_bits_wdata_25),
    .io_out_wdata_bits_wdata_26(AXICmdSplit_io_out_wdata_bits_wdata_26),
    .io_out_wdata_bits_wdata_27(AXICmdSplit_io_out_wdata_bits_wdata_27),
    .io_out_wdata_bits_wdata_28(AXICmdSplit_io_out_wdata_bits_wdata_28),
    .io_out_wdata_bits_wdata_29(AXICmdSplit_io_out_wdata_bits_wdata_29),
    .io_out_wdata_bits_wdata_30(AXICmdSplit_io_out_wdata_bits_wdata_30),
    .io_out_wdata_bits_wdata_31(AXICmdSplit_io_out_wdata_bits_wdata_31),
    .io_out_wdata_bits_wdata_32(AXICmdSplit_io_out_wdata_bits_wdata_32),
    .io_out_wdata_bits_wdata_33(AXICmdSplit_io_out_wdata_bits_wdata_33),
    .io_out_wdata_bits_wdata_34(AXICmdSplit_io_out_wdata_bits_wdata_34),
    .io_out_wdata_bits_wdata_35(AXICmdSplit_io_out_wdata_bits_wdata_35),
    .io_out_wdata_bits_wdata_36(AXICmdSplit_io_out_wdata_bits_wdata_36),
    .io_out_wdata_bits_wdata_37(AXICmdSplit_io_out_wdata_bits_wdata_37),
    .io_out_wdata_bits_wdata_38(AXICmdSplit_io_out_wdata_bits_wdata_38),
    .io_out_wdata_bits_wdata_39(AXICmdSplit_io_out_wdata_bits_wdata_39),
    .io_out_wdata_bits_wdata_40(AXICmdSplit_io_out_wdata_bits_wdata_40),
    .io_out_wdata_bits_wdata_41(AXICmdSplit_io_out_wdata_bits_wdata_41),
    .io_out_wdata_bits_wdata_42(AXICmdSplit_io_out_wdata_bits_wdata_42),
    .io_out_wdata_bits_wdata_43(AXICmdSplit_io_out_wdata_bits_wdata_43),
    .io_out_wdata_bits_wdata_44(AXICmdSplit_io_out_wdata_bits_wdata_44),
    .io_out_wdata_bits_wdata_45(AXICmdSplit_io_out_wdata_bits_wdata_45),
    .io_out_wdata_bits_wdata_46(AXICmdSplit_io_out_wdata_bits_wdata_46),
    .io_out_wdata_bits_wdata_47(AXICmdSplit_io_out_wdata_bits_wdata_47),
    .io_out_wdata_bits_wdata_48(AXICmdSplit_io_out_wdata_bits_wdata_48),
    .io_out_wdata_bits_wdata_49(AXICmdSplit_io_out_wdata_bits_wdata_49),
    .io_out_wdata_bits_wdata_50(AXICmdSplit_io_out_wdata_bits_wdata_50),
    .io_out_wdata_bits_wdata_51(AXICmdSplit_io_out_wdata_bits_wdata_51),
    .io_out_wdata_bits_wdata_52(AXICmdSplit_io_out_wdata_bits_wdata_52),
    .io_out_wdata_bits_wdata_53(AXICmdSplit_io_out_wdata_bits_wdata_53),
    .io_out_wdata_bits_wdata_54(AXICmdSplit_io_out_wdata_bits_wdata_54),
    .io_out_wdata_bits_wdata_55(AXICmdSplit_io_out_wdata_bits_wdata_55),
    .io_out_wdata_bits_wdata_56(AXICmdSplit_io_out_wdata_bits_wdata_56),
    .io_out_wdata_bits_wdata_57(AXICmdSplit_io_out_wdata_bits_wdata_57),
    .io_out_wdata_bits_wdata_58(AXICmdSplit_io_out_wdata_bits_wdata_58),
    .io_out_wdata_bits_wdata_59(AXICmdSplit_io_out_wdata_bits_wdata_59),
    .io_out_wdata_bits_wdata_60(AXICmdSplit_io_out_wdata_bits_wdata_60),
    .io_out_wdata_bits_wdata_61(AXICmdSplit_io_out_wdata_bits_wdata_61),
    .io_out_wdata_bits_wdata_62(AXICmdSplit_io_out_wdata_bits_wdata_62),
    .io_out_wdata_bits_wdata_63(AXICmdSplit_io_out_wdata_bits_wdata_63),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_rresp_valid(AXICmdSplit_io_out_rresp_valid),
    .io_out_rresp_bits_rdata_0(AXICmdSplit_io_out_rresp_bits_rdata_0),
    .io_out_rresp_bits_rdata_1(AXICmdSplit_io_out_rresp_bits_rdata_1),
    .io_out_rresp_bits_rdata_2(AXICmdSplit_io_out_rresp_bits_rdata_2),
    .io_out_rresp_bits_rdata_3(AXICmdSplit_io_out_rresp_bits_rdata_3),
    .io_out_rresp_bits_rdata_4(AXICmdSplit_io_out_rresp_bits_rdata_4),
    .io_out_rresp_bits_rdata_5(AXICmdSplit_io_out_rresp_bits_rdata_5),
    .io_out_rresp_bits_rdata_6(AXICmdSplit_io_out_rresp_bits_rdata_6),
    .io_out_rresp_bits_rdata_7(AXICmdSplit_io_out_rresp_bits_rdata_7),
    .io_out_rresp_bits_rdata_8(AXICmdSplit_io_out_rresp_bits_rdata_8),
    .io_out_rresp_bits_rdata_9(AXICmdSplit_io_out_rresp_bits_rdata_9),
    .io_out_rresp_bits_rdata_10(AXICmdSplit_io_out_rresp_bits_rdata_10),
    .io_out_rresp_bits_rdata_11(AXICmdSplit_io_out_rresp_bits_rdata_11),
    .io_out_rresp_bits_rdata_12(AXICmdSplit_io_out_rresp_bits_rdata_12),
    .io_out_rresp_bits_rdata_13(AXICmdSplit_io_out_rresp_bits_rdata_13),
    .io_out_rresp_bits_rdata_14(AXICmdSplit_io_out_rresp_bits_rdata_14),
    .io_out_rresp_bits_rdata_15(AXICmdSplit_io_out_rresp_bits_rdata_15),
    .io_out_rresp_bits_rdata_16(AXICmdSplit_io_out_rresp_bits_rdata_16),
    .io_out_rresp_bits_rdata_17(AXICmdSplit_io_out_rresp_bits_rdata_17),
    .io_out_rresp_bits_rdata_18(AXICmdSplit_io_out_rresp_bits_rdata_18),
    .io_out_rresp_bits_rdata_19(AXICmdSplit_io_out_rresp_bits_rdata_19),
    .io_out_rresp_bits_rdata_20(AXICmdSplit_io_out_rresp_bits_rdata_20),
    .io_out_rresp_bits_rdata_21(AXICmdSplit_io_out_rresp_bits_rdata_21),
    .io_out_rresp_bits_rdata_22(AXICmdSplit_io_out_rresp_bits_rdata_22),
    .io_out_rresp_bits_rdata_23(AXICmdSplit_io_out_rresp_bits_rdata_23),
    .io_out_rresp_bits_rdata_24(AXICmdSplit_io_out_rresp_bits_rdata_24),
    .io_out_rresp_bits_rdata_25(AXICmdSplit_io_out_rresp_bits_rdata_25),
    .io_out_rresp_bits_rdata_26(AXICmdSplit_io_out_rresp_bits_rdata_26),
    .io_out_rresp_bits_rdata_27(AXICmdSplit_io_out_rresp_bits_rdata_27),
    .io_out_rresp_bits_rdata_28(AXICmdSplit_io_out_rresp_bits_rdata_28),
    .io_out_rresp_bits_rdata_29(AXICmdSplit_io_out_rresp_bits_rdata_29),
    .io_out_rresp_bits_rdata_30(AXICmdSplit_io_out_rresp_bits_rdata_30),
    .io_out_rresp_bits_rdata_31(AXICmdSplit_io_out_rresp_bits_rdata_31),
    .io_out_rresp_bits_rdata_32(AXICmdSplit_io_out_rresp_bits_rdata_32),
    .io_out_rresp_bits_rdata_33(AXICmdSplit_io_out_rresp_bits_rdata_33),
    .io_out_rresp_bits_rdata_34(AXICmdSplit_io_out_rresp_bits_rdata_34),
    .io_out_rresp_bits_rdata_35(AXICmdSplit_io_out_rresp_bits_rdata_35),
    .io_out_rresp_bits_rdata_36(AXICmdSplit_io_out_rresp_bits_rdata_36),
    .io_out_rresp_bits_rdata_37(AXICmdSplit_io_out_rresp_bits_rdata_37),
    .io_out_rresp_bits_rdata_38(AXICmdSplit_io_out_rresp_bits_rdata_38),
    .io_out_rresp_bits_rdata_39(AXICmdSplit_io_out_rresp_bits_rdata_39),
    .io_out_rresp_bits_rdata_40(AXICmdSplit_io_out_rresp_bits_rdata_40),
    .io_out_rresp_bits_rdata_41(AXICmdSplit_io_out_rresp_bits_rdata_41),
    .io_out_rresp_bits_rdata_42(AXICmdSplit_io_out_rresp_bits_rdata_42),
    .io_out_rresp_bits_rdata_43(AXICmdSplit_io_out_rresp_bits_rdata_43),
    .io_out_rresp_bits_rdata_44(AXICmdSplit_io_out_rresp_bits_rdata_44),
    .io_out_rresp_bits_rdata_45(AXICmdSplit_io_out_rresp_bits_rdata_45),
    .io_out_rresp_bits_rdata_46(AXICmdSplit_io_out_rresp_bits_rdata_46),
    .io_out_rresp_bits_rdata_47(AXICmdSplit_io_out_rresp_bits_rdata_47),
    .io_out_rresp_bits_rdata_48(AXICmdSplit_io_out_rresp_bits_rdata_48),
    .io_out_rresp_bits_rdata_49(AXICmdSplit_io_out_rresp_bits_rdata_49),
    .io_out_rresp_bits_rdata_50(AXICmdSplit_io_out_rresp_bits_rdata_50),
    .io_out_rresp_bits_rdata_51(AXICmdSplit_io_out_rresp_bits_rdata_51),
    .io_out_rresp_bits_rdata_52(AXICmdSplit_io_out_rresp_bits_rdata_52),
    .io_out_rresp_bits_rdata_53(AXICmdSplit_io_out_rresp_bits_rdata_53),
    .io_out_rresp_bits_rdata_54(AXICmdSplit_io_out_rresp_bits_rdata_54),
    .io_out_rresp_bits_rdata_55(AXICmdSplit_io_out_rresp_bits_rdata_55),
    .io_out_rresp_bits_rdata_56(AXICmdSplit_io_out_rresp_bits_rdata_56),
    .io_out_rresp_bits_rdata_57(AXICmdSplit_io_out_rresp_bits_rdata_57),
    .io_out_rresp_bits_rdata_58(AXICmdSplit_io_out_rresp_bits_rdata_58),
    .io_out_rresp_bits_rdata_59(AXICmdSplit_io_out_rresp_bits_rdata_59),
    .io_out_rresp_bits_rdata_60(AXICmdSplit_io_out_rresp_bits_rdata_60),
    .io_out_rresp_bits_rdata_61(AXICmdSplit_io_out_rresp_bits_rdata_61),
    .io_out_rresp_bits_rdata_62(AXICmdSplit_io_out_rresp_bits_rdata_62),
    .io_out_rresp_bits_rdata_63(AXICmdSplit_io_out_rresp_bits_rdata_63),
    .io_out_rresp_bits_tag(AXICmdSplit_io_out_rresp_bits_tag),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@107884.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_rawAddr(AXICmdIssue_io_in_cmd_bits_rawAddr),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wdata_16(AXICmdIssue_io_in_wdata_bits_wdata_16),
    .io_in_wdata_bits_wdata_17(AXICmdIssue_io_in_wdata_bits_wdata_17),
    .io_in_wdata_bits_wdata_18(AXICmdIssue_io_in_wdata_bits_wdata_18),
    .io_in_wdata_bits_wdata_19(AXICmdIssue_io_in_wdata_bits_wdata_19),
    .io_in_wdata_bits_wdata_20(AXICmdIssue_io_in_wdata_bits_wdata_20),
    .io_in_wdata_bits_wdata_21(AXICmdIssue_io_in_wdata_bits_wdata_21),
    .io_in_wdata_bits_wdata_22(AXICmdIssue_io_in_wdata_bits_wdata_22),
    .io_in_wdata_bits_wdata_23(AXICmdIssue_io_in_wdata_bits_wdata_23),
    .io_in_wdata_bits_wdata_24(AXICmdIssue_io_in_wdata_bits_wdata_24),
    .io_in_wdata_bits_wdata_25(AXICmdIssue_io_in_wdata_bits_wdata_25),
    .io_in_wdata_bits_wdata_26(AXICmdIssue_io_in_wdata_bits_wdata_26),
    .io_in_wdata_bits_wdata_27(AXICmdIssue_io_in_wdata_bits_wdata_27),
    .io_in_wdata_bits_wdata_28(AXICmdIssue_io_in_wdata_bits_wdata_28),
    .io_in_wdata_bits_wdata_29(AXICmdIssue_io_in_wdata_bits_wdata_29),
    .io_in_wdata_bits_wdata_30(AXICmdIssue_io_in_wdata_bits_wdata_30),
    .io_in_wdata_bits_wdata_31(AXICmdIssue_io_in_wdata_bits_wdata_31),
    .io_in_wdata_bits_wdata_32(AXICmdIssue_io_in_wdata_bits_wdata_32),
    .io_in_wdata_bits_wdata_33(AXICmdIssue_io_in_wdata_bits_wdata_33),
    .io_in_wdata_bits_wdata_34(AXICmdIssue_io_in_wdata_bits_wdata_34),
    .io_in_wdata_bits_wdata_35(AXICmdIssue_io_in_wdata_bits_wdata_35),
    .io_in_wdata_bits_wdata_36(AXICmdIssue_io_in_wdata_bits_wdata_36),
    .io_in_wdata_bits_wdata_37(AXICmdIssue_io_in_wdata_bits_wdata_37),
    .io_in_wdata_bits_wdata_38(AXICmdIssue_io_in_wdata_bits_wdata_38),
    .io_in_wdata_bits_wdata_39(AXICmdIssue_io_in_wdata_bits_wdata_39),
    .io_in_wdata_bits_wdata_40(AXICmdIssue_io_in_wdata_bits_wdata_40),
    .io_in_wdata_bits_wdata_41(AXICmdIssue_io_in_wdata_bits_wdata_41),
    .io_in_wdata_bits_wdata_42(AXICmdIssue_io_in_wdata_bits_wdata_42),
    .io_in_wdata_bits_wdata_43(AXICmdIssue_io_in_wdata_bits_wdata_43),
    .io_in_wdata_bits_wdata_44(AXICmdIssue_io_in_wdata_bits_wdata_44),
    .io_in_wdata_bits_wdata_45(AXICmdIssue_io_in_wdata_bits_wdata_45),
    .io_in_wdata_bits_wdata_46(AXICmdIssue_io_in_wdata_bits_wdata_46),
    .io_in_wdata_bits_wdata_47(AXICmdIssue_io_in_wdata_bits_wdata_47),
    .io_in_wdata_bits_wdata_48(AXICmdIssue_io_in_wdata_bits_wdata_48),
    .io_in_wdata_bits_wdata_49(AXICmdIssue_io_in_wdata_bits_wdata_49),
    .io_in_wdata_bits_wdata_50(AXICmdIssue_io_in_wdata_bits_wdata_50),
    .io_in_wdata_bits_wdata_51(AXICmdIssue_io_in_wdata_bits_wdata_51),
    .io_in_wdata_bits_wdata_52(AXICmdIssue_io_in_wdata_bits_wdata_52),
    .io_in_wdata_bits_wdata_53(AXICmdIssue_io_in_wdata_bits_wdata_53),
    .io_in_wdata_bits_wdata_54(AXICmdIssue_io_in_wdata_bits_wdata_54),
    .io_in_wdata_bits_wdata_55(AXICmdIssue_io_in_wdata_bits_wdata_55),
    .io_in_wdata_bits_wdata_56(AXICmdIssue_io_in_wdata_bits_wdata_56),
    .io_in_wdata_bits_wdata_57(AXICmdIssue_io_in_wdata_bits_wdata_57),
    .io_in_wdata_bits_wdata_58(AXICmdIssue_io_in_wdata_bits_wdata_58),
    .io_in_wdata_bits_wdata_59(AXICmdIssue_io_in_wdata_bits_wdata_59),
    .io_in_wdata_bits_wdata_60(AXICmdIssue_io_in_wdata_bits_wdata_60),
    .io_in_wdata_bits_wdata_61(AXICmdIssue_io_in_wdata_bits_wdata_61),
    .io_in_wdata_bits_wdata_62(AXICmdIssue_io_in_wdata_bits_wdata_62),
    .io_in_wdata_bits_wdata_63(AXICmdIssue_io_in_wdata_bits_wdata_63),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_rresp_valid(AXICmdIssue_io_in_rresp_valid),
    .io_in_rresp_bits_rdata_0(AXICmdIssue_io_in_rresp_bits_rdata_0),
    .io_in_rresp_bits_rdata_1(AXICmdIssue_io_in_rresp_bits_rdata_1),
    .io_in_rresp_bits_rdata_2(AXICmdIssue_io_in_rresp_bits_rdata_2),
    .io_in_rresp_bits_rdata_3(AXICmdIssue_io_in_rresp_bits_rdata_3),
    .io_in_rresp_bits_rdata_4(AXICmdIssue_io_in_rresp_bits_rdata_4),
    .io_in_rresp_bits_rdata_5(AXICmdIssue_io_in_rresp_bits_rdata_5),
    .io_in_rresp_bits_rdata_6(AXICmdIssue_io_in_rresp_bits_rdata_6),
    .io_in_rresp_bits_rdata_7(AXICmdIssue_io_in_rresp_bits_rdata_7),
    .io_in_rresp_bits_rdata_8(AXICmdIssue_io_in_rresp_bits_rdata_8),
    .io_in_rresp_bits_rdata_9(AXICmdIssue_io_in_rresp_bits_rdata_9),
    .io_in_rresp_bits_rdata_10(AXICmdIssue_io_in_rresp_bits_rdata_10),
    .io_in_rresp_bits_rdata_11(AXICmdIssue_io_in_rresp_bits_rdata_11),
    .io_in_rresp_bits_rdata_12(AXICmdIssue_io_in_rresp_bits_rdata_12),
    .io_in_rresp_bits_rdata_13(AXICmdIssue_io_in_rresp_bits_rdata_13),
    .io_in_rresp_bits_rdata_14(AXICmdIssue_io_in_rresp_bits_rdata_14),
    .io_in_rresp_bits_rdata_15(AXICmdIssue_io_in_rresp_bits_rdata_15),
    .io_in_rresp_bits_rdata_16(AXICmdIssue_io_in_rresp_bits_rdata_16),
    .io_in_rresp_bits_rdata_17(AXICmdIssue_io_in_rresp_bits_rdata_17),
    .io_in_rresp_bits_rdata_18(AXICmdIssue_io_in_rresp_bits_rdata_18),
    .io_in_rresp_bits_rdata_19(AXICmdIssue_io_in_rresp_bits_rdata_19),
    .io_in_rresp_bits_rdata_20(AXICmdIssue_io_in_rresp_bits_rdata_20),
    .io_in_rresp_bits_rdata_21(AXICmdIssue_io_in_rresp_bits_rdata_21),
    .io_in_rresp_bits_rdata_22(AXICmdIssue_io_in_rresp_bits_rdata_22),
    .io_in_rresp_bits_rdata_23(AXICmdIssue_io_in_rresp_bits_rdata_23),
    .io_in_rresp_bits_rdata_24(AXICmdIssue_io_in_rresp_bits_rdata_24),
    .io_in_rresp_bits_rdata_25(AXICmdIssue_io_in_rresp_bits_rdata_25),
    .io_in_rresp_bits_rdata_26(AXICmdIssue_io_in_rresp_bits_rdata_26),
    .io_in_rresp_bits_rdata_27(AXICmdIssue_io_in_rresp_bits_rdata_27),
    .io_in_rresp_bits_rdata_28(AXICmdIssue_io_in_rresp_bits_rdata_28),
    .io_in_rresp_bits_rdata_29(AXICmdIssue_io_in_rresp_bits_rdata_29),
    .io_in_rresp_bits_rdata_30(AXICmdIssue_io_in_rresp_bits_rdata_30),
    .io_in_rresp_bits_rdata_31(AXICmdIssue_io_in_rresp_bits_rdata_31),
    .io_in_rresp_bits_rdata_32(AXICmdIssue_io_in_rresp_bits_rdata_32),
    .io_in_rresp_bits_rdata_33(AXICmdIssue_io_in_rresp_bits_rdata_33),
    .io_in_rresp_bits_rdata_34(AXICmdIssue_io_in_rresp_bits_rdata_34),
    .io_in_rresp_bits_rdata_35(AXICmdIssue_io_in_rresp_bits_rdata_35),
    .io_in_rresp_bits_rdata_36(AXICmdIssue_io_in_rresp_bits_rdata_36),
    .io_in_rresp_bits_rdata_37(AXICmdIssue_io_in_rresp_bits_rdata_37),
    .io_in_rresp_bits_rdata_38(AXICmdIssue_io_in_rresp_bits_rdata_38),
    .io_in_rresp_bits_rdata_39(AXICmdIssue_io_in_rresp_bits_rdata_39),
    .io_in_rresp_bits_rdata_40(AXICmdIssue_io_in_rresp_bits_rdata_40),
    .io_in_rresp_bits_rdata_41(AXICmdIssue_io_in_rresp_bits_rdata_41),
    .io_in_rresp_bits_rdata_42(AXICmdIssue_io_in_rresp_bits_rdata_42),
    .io_in_rresp_bits_rdata_43(AXICmdIssue_io_in_rresp_bits_rdata_43),
    .io_in_rresp_bits_rdata_44(AXICmdIssue_io_in_rresp_bits_rdata_44),
    .io_in_rresp_bits_rdata_45(AXICmdIssue_io_in_rresp_bits_rdata_45),
    .io_in_rresp_bits_rdata_46(AXICmdIssue_io_in_rresp_bits_rdata_46),
    .io_in_rresp_bits_rdata_47(AXICmdIssue_io_in_rresp_bits_rdata_47),
    .io_in_rresp_bits_rdata_48(AXICmdIssue_io_in_rresp_bits_rdata_48),
    .io_in_rresp_bits_rdata_49(AXICmdIssue_io_in_rresp_bits_rdata_49),
    .io_in_rresp_bits_rdata_50(AXICmdIssue_io_in_rresp_bits_rdata_50),
    .io_in_rresp_bits_rdata_51(AXICmdIssue_io_in_rresp_bits_rdata_51),
    .io_in_rresp_bits_rdata_52(AXICmdIssue_io_in_rresp_bits_rdata_52),
    .io_in_rresp_bits_rdata_53(AXICmdIssue_io_in_rresp_bits_rdata_53),
    .io_in_rresp_bits_rdata_54(AXICmdIssue_io_in_rresp_bits_rdata_54),
    .io_in_rresp_bits_rdata_55(AXICmdIssue_io_in_rresp_bits_rdata_55),
    .io_in_rresp_bits_rdata_56(AXICmdIssue_io_in_rresp_bits_rdata_56),
    .io_in_rresp_bits_rdata_57(AXICmdIssue_io_in_rresp_bits_rdata_57),
    .io_in_rresp_bits_rdata_58(AXICmdIssue_io_in_rresp_bits_rdata_58),
    .io_in_rresp_bits_rdata_59(AXICmdIssue_io_in_rresp_bits_rdata_59),
    .io_in_rresp_bits_rdata_60(AXICmdIssue_io_in_rresp_bits_rdata_60),
    .io_in_rresp_bits_rdata_61(AXICmdIssue_io_in_rresp_bits_rdata_61),
    .io_in_rresp_bits_rdata_62(AXICmdIssue_io_in_rresp_bits_rdata_62),
    .io_in_rresp_bits_rdata_63(AXICmdIssue_io_in_rresp_bits_rdata_63),
    .io_in_rresp_bits_tag(AXICmdIssue_io_in_rresp_bits_tag),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_rawAddr(AXICmdIssue_io_out_cmd_bits_rawAddr),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wdata_16(AXICmdIssue_io_out_wdata_bits_wdata_16),
    .io_out_wdata_bits_wdata_17(AXICmdIssue_io_out_wdata_bits_wdata_17),
    .io_out_wdata_bits_wdata_18(AXICmdIssue_io_out_wdata_bits_wdata_18),
    .io_out_wdata_bits_wdata_19(AXICmdIssue_io_out_wdata_bits_wdata_19),
    .io_out_wdata_bits_wdata_20(AXICmdIssue_io_out_wdata_bits_wdata_20),
    .io_out_wdata_bits_wdata_21(AXICmdIssue_io_out_wdata_bits_wdata_21),
    .io_out_wdata_bits_wdata_22(AXICmdIssue_io_out_wdata_bits_wdata_22),
    .io_out_wdata_bits_wdata_23(AXICmdIssue_io_out_wdata_bits_wdata_23),
    .io_out_wdata_bits_wdata_24(AXICmdIssue_io_out_wdata_bits_wdata_24),
    .io_out_wdata_bits_wdata_25(AXICmdIssue_io_out_wdata_bits_wdata_25),
    .io_out_wdata_bits_wdata_26(AXICmdIssue_io_out_wdata_bits_wdata_26),
    .io_out_wdata_bits_wdata_27(AXICmdIssue_io_out_wdata_bits_wdata_27),
    .io_out_wdata_bits_wdata_28(AXICmdIssue_io_out_wdata_bits_wdata_28),
    .io_out_wdata_bits_wdata_29(AXICmdIssue_io_out_wdata_bits_wdata_29),
    .io_out_wdata_bits_wdata_30(AXICmdIssue_io_out_wdata_bits_wdata_30),
    .io_out_wdata_bits_wdata_31(AXICmdIssue_io_out_wdata_bits_wdata_31),
    .io_out_wdata_bits_wdata_32(AXICmdIssue_io_out_wdata_bits_wdata_32),
    .io_out_wdata_bits_wdata_33(AXICmdIssue_io_out_wdata_bits_wdata_33),
    .io_out_wdata_bits_wdata_34(AXICmdIssue_io_out_wdata_bits_wdata_34),
    .io_out_wdata_bits_wdata_35(AXICmdIssue_io_out_wdata_bits_wdata_35),
    .io_out_wdata_bits_wdata_36(AXICmdIssue_io_out_wdata_bits_wdata_36),
    .io_out_wdata_bits_wdata_37(AXICmdIssue_io_out_wdata_bits_wdata_37),
    .io_out_wdata_bits_wdata_38(AXICmdIssue_io_out_wdata_bits_wdata_38),
    .io_out_wdata_bits_wdata_39(AXICmdIssue_io_out_wdata_bits_wdata_39),
    .io_out_wdata_bits_wdata_40(AXICmdIssue_io_out_wdata_bits_wdata_40),
    .io_out_wdata_bits_wdata_41(AXICmdIssue_io_out_wdata_bits_wdata_41),
    .io_out_wdata_bits_wdata_42(AXICmdIssue_io_out_wdata_bits_wdata_42),
    .io_out_wdata_bits_wdata_43(AXICmdIssue_io_out_wdata_bits_wdata_43),
    .io_out_wdata_bits_wdata_44(AXICmdIssue_io_out_wdata_bits_wdata_44),
    .io_out_wdata_bits_wdata_45(AXICmdIssue_io_out_wdata_bits_wdata_45),
    .io_out_wdata_bits_wdata_46(AXICmdIssue_io_out_wdata_bits_wdata_46),
    .io_out_wdata_bits_wdata_47(AXICmdIssue_io_out_wdata_bits_wdata_47),
    .io_out_wdata_bits_wdata_48(AXICmdIssue_io_out_wdata_bits_wdata_48),
    .io_out_wdata_bits_wdata_49(AXICmdIssue_io_out_wdata_bits_wdata_49),
    .io_out_wdata_bits_wdata_50(AXICmdIssue_io_out_wdata_bits_wdata_50),
    .io_out_wdata_bits_wdata_51(AXICmdIssue_io_out_wdata_bits_wdata_51),
    .io_out_wdata_bits_wdata_52(AXICmdIssue_io_out_wdata_bits_wdata_52),
    .io_out_wdata_bits_wdata_53(AXICmdIssue_io_out_wdata_bits_wdata_53),
    .io_out_wdata_bits_wdata_54(AXICmdIssue_io_out_wdata_bits_wdata_54),
    .io_out_wdata_bits_wdata_55(AXICmdIssue_io_out_wdata_bits_wdata_55),
    .io_out_wdata_bits_wdata_56(AXICmdIssue_io_out_wdata_bits_wdata_56),
    .io_out_wdata_bits_wdata_57(AXICmdIssue_io_out_wdata_bits_wdata_57),
    .io_out_wdata_bits_wdata_58(AXICmdIssue_io_out_wdata_bits_wdata_58),
    .io_out_wdata_bits_wdata_59(AXICmdIssue_io_out_wdata_bits_wdata_59),
    .io_out_wdata_bits_wdata_60(AXICmdIssue_io_out_wdata_bits_wdata_60),
    .io_out_wdata_bits_wdata_61(AXICmdIssue_io_out_wdata_bits_wdata_61),
    .io_out_wdata_bits_wdata_62(AXICmdIssue_io_out_wdata_bits_wdata_62),
    .io_out_wdata_bits_wdata_63(AXICmdIssue_io_out_wdata_bits_wdata_63),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_rresp_valid(AXICmdIssue_io_out_rresp_valid),
    .io_out_rresp_bits_rdata_0(AXICmdIssue_io_out_rresp_bits_rdata_0),
    .io_out_rresp_bits_rdata_1(AXICmdIssue_io_out_rresp_bits_rdata_1),
    .io_out_rresp_bits_rdata_2(AXICmdIssue_io_out_rresp_bits_rdata_2),
    .io_out_rresp_bits_rdata_3(AXICmdIssue_io_out_rresp_bits_rdata_3),
    .io_out_rresp_bits_rdata_4(AXICmdIssue_io_out_rresp_bits_rdata_4),
    .io_out_rresp_bits_rdata_5(AXICmdIssue_io_out_rresp_bits_rdata_5),
    .io_out_rresp_bits_rdata_6(AXICmdIssue_io_out_rresp_bits_rdata_6),
    .io_out_rresp_bits_rdata_7(AXICmdIssue_io_out_rresp_bits_rdata_7),
    .io_out_rresp_bits_rdata_8(AXICmdIssue_io_out_rresp_bits_rdata_8),
    .io_out_rresp_bits_rdata_9(AXICmdIssue_io_out_rresp_bits_rdata_9),
    .io_out_rresp_bits_rdata_10(AXICmdIssue_io_out_rresp_bits_rdata_10),
    .io_out_rresp_bits_rdata_11(AXICmdIssue_io_out_rresp_bits_rdata_11),
    .io_out_rresp_bits_rdata_12(AXICmdIssue_io_out_rresp_bits_rdata_12),
    .io_out_rresp_bits_rdata_13(AXICmdIssue_io_out_rresp_bits_rdata_13),
    .io_out_rresp_bits_rdata_14(AXICmdIssue_io_out_rresp_bits_rdata_14),
    .io_out_rresp_bits_rdata_15(AXICmdIssue_io_out_rresp_bits_rdata_15),
    .io_out_rresp_bits_rdata_16(AXICmdIssue_io_out_rresp_bits_rdata_16),
    .io_out_rresp_bits_rdata_17(AXICmdIssue_io_out_rresp_bits_rdata_17),
    .io_out_rresp_bits_rdata_18(AXICmdIssue_io_out_rresp_bits_rdata_18),
    .io_out_rresp_bits_rdata_19(AXICmdIssue_io_out_rresp_bits_rdata_19),
    .io_out_rresp_bits_rdata_20(AXICmdIssue_io_out_rresp_bits_rdata_20),
    .io_out_rresp_bits_rdata_21(AXICmdIssue_io_out_rresp_bits_rdata_21),
    .io_out_rresp_bits_rdata_22(AXICmdIssue_io_out_rresp_bits_rdata_22),
    .io_out_rresp_bits_rdata_23(AXICmdIssue_io_out_rresp_bits_rdata_23),
    .io_out_rresp_bits_rdata_24(AXICmdIssue_io_out_rresp_bits_rdata_24),
    .io_out_rresp_bits_rdata_25(AXICmdIssue_io_out_rresp_bits_rdata_25),
    .io_out_rresp_bits_rdata_26(AXICmdIssue_io_out_rresp_bits_rdata_26),
    .io_out_rresp_bits_rdata_27(AXICmdIssue_io_out_rresp_bits_rdata_27),
    .io_out_rresp_bits_rdata_28(AXICmdIssue_io_out_rresp_bits_rdata_28),
    .io_out_rresp_bits_rdata_29(AXICmdIssue_io_out_rresp_bits_rdata_29),
    .io_out_rresp_bits_rdata_30(AXICmdIssue_io_out_rresp_bits_rdata_30),
    .io_out_rresp_bits_rdata_31(AXICmdIssue_io_out_rresp_bits_rdata_31),
    .io_out_rresp_bits_rdata_32(AXICmdIssue_io_out_rresp_bits_rdata_32),
    .io_out_rresp_bits_rdata_33(AXICmdIssue_io_out_rresp_bits_rdata_33),
    .io_out_rresp_bits_rdata_34(AXICmdIssue_io_out_rresp_bits_rdata_34),
    .io_out_rresp_bits_rdata_35(AXICmdIssue_io_out_rresp_bits_rdata_35),
    .io_out_rresp_bits_rdata_36(AXICmdIssue_io_out_rresp_bits_rdata_36),
    .io_out_rresp_bits_rdata_37(AXICmdIssue_io_out_rresp_bits_rdata_37),
    .io_out_rresp_bits_rdata_38(AXICmdIssue_io_out_rresp_bits_rdata_38),
    .io_out_rresp_bits_rdata_39(AXICmdIssue_io_out_rresp_bits_rdata_39),
    .io_out_rresp_bits_rdata_40(AXICmdIssue_io_out_rresp_bits_rdata_40),
    .io_out_rresp_bits_rdata_41(AXICmdIssue_io_out_rresp_bits_rdata_41),
    .io_out_rresp_bits_rdata_42(AXICmdIssue_io_out_rresp_bits_rdata_42),
    .io_out_rresp_bits_rdata_43(AXICmdIssue_io_out_rresp_bits_rdata_43),
    .io_out_rresp_bits_rdata_44(AXICmdIssue_io_out_rresp_bits_rdata_44),
    .io_out_rresp_bits_rdata_45(AXICmdIssue_io_out_rresp_bits_rdata_45),
    .io_out_rresp_bits_rdata_46(AXICmdIssue_io_out_rresp_bits_rdata_46),
    .io_out_rresp_bits_rdata_47(AXICmdIssue_io_out_rresp_bits_rdata_47),
    .io_out_rresp_bits_rdata_48(AXICmdIssue_io_out_rresp_bits_rdata_48),
    .io_out_rresp_bits_rdata_49(AXICmdIssue_io_out_rresp_bits_rdata_49),
    .io_out_rresp_bits_rdata_50(AXICmdIssue_io_out_rresp_bits_rdata_50),
    .io_out_rresp_bits_rdata_51(AXICmdIssue_io_out_rresp_bits_rdata_51),
    .io_out_rresp_bits_rdata_52(AXICmdIssue_io_out_rresp_bits_rdata_52),
    .io_out_rresp_bits_rdata_53(AXICmdIssue_io_out_rresp_bits_rdata_53),
    .io_out_rresp_bits_rdata_54(AXICmdIssue_io_out_rresp_bits_rdata_54),
    .io_out_rresp_bits_rdata_55(AXICmdIssue_io_out_rresp_bits_rdata_55),
    .io_out_rresp_bits_rdata_56(AXICmdIssue_io_out_rresp_bits_rdata_56),
    .io_out_rresp_bits_rdata_57(AXICmdIssue_io_out_rresp_bits_rdata_57),
    .io_out_rresp_bits_rdata_58(AXICmdIssue_io_out_rresp_bits_rdata_58),
    .io_out_rresp_bits_rdata_59(AXICmdIssue_io_out_rresp_bits_rdata_59),
    .io_out_rresp_bits_rdata_60(AXICmdIssue_io_out_rresp_bits_rdata_60),
    .io_out_rresp_bits_rdata_61(AXICmdIssue_io_out_rresp_bits_rdata_61),
    .io_out_rresp_bits_rdata_62(AXICmdIssue_io_out_rresp_bits_rdata_62),
    .io_out_rresp_bits_rdata_63(AXICmdIssue_io_out_rresp_bits_rdata_63),
    .io_out_rresp_bits_tag(AXICmdIssue_io_out_rresp_bits_tag),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign _T_2030 = _T_2028 + 64'h1; // @[DRAMArbiter.scala 123:18:@108309.6]
  assign _T_2031 = _T_2028 + 64'h1; // @[DRAMArbiter.scala 123:18:@108310.6]
  assign _GEN_0 = io_enable ? _T_2031 : _T_2028; // @[DRAMArbiter.scala 122:19:@108308.4]
  assign _T_2032 = io_dram_rresp_valid & io_dram_rresp_ready; // @[DRAMArbiter.scala 139:60:@108314.4]
  assign _T_2039 = io_dram_wdata_valid & io_dram_wdata_ready; // @[DRAMArbiter.scala 140:57:@108321.4]
  assign _T_2044 = _T_2042 + 64'h1; // @[DRAMArbiter.scala 123:18:@108324.6]
  assign _T_2045 = _T_2042 + 64'h1; // @[DRAMArbiter.scala 123:18:@108325.6]
  assign _GEN_2 = _T_2039 ? _T_2045 : _T_2042; // @[DRAMArbiter.scala 122:19:@108323.4]
  assign _T_2046 = io_app_stores_0_data_valid & io_app_stores_0_data_ready; // @[DRAMArbiter.scala 141:70:@108328.4]
  assign _T_2051 = _T_2049 + 64'h1; // @[DRAMArbiter.scala 123:18:@108331.6]
  assign _T_2052 = _T_2049 + 64'h1; // @[DRAMArbiter.scala 123:18:@108332.6]
  assign _GEN_3 = _T_2046 ? _T_2052 : _T_2049; // @[DRAMArbiter.scala 122:19:@108330.4]
  assign _T_2053 = io_dram_cmd_ready & io_dram_cmd_valid; // @[DRAMArbiter.scala 144:52:@108336.4]
  assign _T_2058 = _T_2056 + 64'h1; // @[DRAMArbiter.scala 123:18:@108339.6]
  assign _T_2059 = _T_2056 + 64'h1; // @[DRAMArbiter.scala 123:18:@108340.6]
  assign _GEN_4 = _T_2053 ? _T_2059 : _T_2056; // @[DRAMArbiter.scala 122:19:@108338.4]
  assign _T_2062 = io_dram_cmd_bits_isWr == 1'h0; // @[DRAMArbiter.scala 145:74:@108345.4]
  assign _T_2063 = _T_2053 & _T_2062; // @[DRAMArbiter.scala 145:72:@108346.4]
  assign _T_2068 = _T_2066 + 64'h1; // @[DRAMArbiter.scala 123:18:@108349.6]
  assign _T_2069 = _T_2066 + 64'h1; // @[DRAMArbiter.scala 123:18:@108350.6]
  assign _GEN_5 = _T_2063 ? _T_2069 : _T_2066; // @[DRAMArbiter.scala 122:19:@108348.4]
  assign _T_2071 = _T_2053 & io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 146:72:@108355.4]
  assign _T_2076 = _T_2074 + 64'h1; // @[DRAMArbiter.scala 123:18:@108358.6]
  assign _T_2077 = _T_2074 + 64'h1; // @[DRAMArbiter.scala 123:18:@108359.6]
  assign _GEN_6 = _T_2071 ? _T_2077 : _T_2074; // @[DRAMArbiter.scala 122:19:@108357.4]
  assign _T_2078 = io_enable & io_app_loads_0_cmd_valid; // @[DRAMArbiter.scala 150:59:@108363.4]
  assign _T_2079 = _T_2078 & io_app_loads_0_cmd_ready; // @[DRAMArbiter.scala 150:76:@108364.4]
  assign _T_2084 = _T_2082 + 64'h1; // @[DRAMArbiter.scala 123:18:@108367.6]
  assign _T_2085 = _T_2082 + 64'h1; // @[DRAMArbiter.scala 123:18:@108368.6]
  assign _GEN_7 = _T_2079 ? _T_2085 : _T_2082; // @[DRAMArbiter.scala 122:19:@108366.4]
  assign _T_2086 = io_enable & io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 156:60:@108372.4]
  assign _T_2087 = _T_2086 & io_app_stores_0_cmd_ready; // @[DRAMArbiter.scala 156:78:@108373.4]
  assign _T_2092 = _T_2090 + 64'h1; // @[DRAMArbiter.scala 123:18:@108376.6]
  assign _T_2093 = _T_2090 + 64'h1; // @[DRAMArbiter.scala 123:18:@108377.6]
  assign _GEN_8 = _T_2087 ? _T_2093 : _T_2090; // @[DRAMArbiter.scala 122:19:@108375.4]
  assign _T_2099 = _T_2097 + 64'h1; // @[DRAMArbiter.scala 123:18:@108384.6]
  assign _T_2100 = _T_2097 + 64'h1; // @[DRAMArbiter.scala 123:18:@108385.6]
  assign _GEN_9 = _T_2032 ? _T_2100 : _T_2097; // @[DRAMArbiter.scala 122:19:@108383.4]
  assign _T_2102 = io_dram_rresp_ready == 1'h0; // @[DRAMArbiter.scala 161:56:@108389.4]
  assign _T_2103 = io_dram_rresp_valid & _T_2102; // @[DRAMArbiter.scala 161:54:@108390.4]
  assign _T_2108 = _T_2106 + 64'h1; // @[DRAMArbiter.scala 123:18:@108393.6]
  assign _T_2109 = _T_2106 + 64'h1; // @[DRAMArbiter.scala 123:18:@108394.6]
  assign _GEN_10 = _T_2103 ? _T_2109 : _T_2106; // @[DRAMArbiter.scala 122:19:@108392.4]
  assign _T_2111 = io_dram_rresp_valid == 1'h0; // @[DRAMArbiter.scala 162:34:@108398.4]
  assign _T_2112 = _T_2111 & io_dram_rresp_ready; // @[DRAMArbiter.scala 162:55:@108399.4]
  assign _T_2117 = _T_2115 + 64'h1; // @[DRAMArbiter.scala 123:18:@108402.6]
  assign _T_2118 = _T_2115 + 64'h1; // @[DRAMArbiter.scala 123:18:@108403.6]
  assign _GEN_11 = _T_2112 ? _T_2118 : _T_2115; // @[DRAMArbiter.scala 122:19:@108401.4]
  assign _T_2125 = io_dram_rresp_bits_tag[7:0]; // @[FringeBundles.scala 132:28:@108411.4]
  assign _T_2129 = _T_2125 == 8'h0; // @[DRAMArbiter.scala 165:116:@108417.4]
  assign _T_2130 = _T_2032 & _T_2129; // @[DRAMArbiter.scala 165:78:@108418.4]
  assign _T_2135 = _T_2133 + 64'h1; // @[DRAMArbiter.scala 123:18:@108421.6]
  assign _T_2136 = _T_2133 + 64'h1; // @[DRAMArbiter.scala 123:18:@108422.6]
  assign _GEN_12 = _T_2130 ? _T_2136 : _T_2133; // @[DRAMArbiter.scala 122:19:@108420.4]
  assign _T_2137 = io_dram_wresp_valid & io_dram_wresp_ready; // @[DRAMArbiter.scala 167:54:@108426.4]
  assign _T_2142 = _T_2140 + 64'h1; // @[DRAMArbiter.scala 123:18:@108429.6]
  assign _T_2143 = _T_2140 + 64'h1; // @[DRAMArbiter.scala 123:18:@108430.6]
  assign _GEN_13 = _T_2137 ? _T_2143 : _T_2140; // @[DRAMArbiter.scala 122:19:@108428.4]
  assign _T_2145 = io_dram_wresp_ready == 1'h0; // @[DRAMArbiter.scala 168:56:@108434.4]
  assign _T_2146 = io_dram_wresp_valid & _T_2145; // @[DRAMArbiter.scala 168:54:@108435.4]
  assign _T_2151 = _T_2149 + 64'h1; // @[DRAMArbiter.scala 123:18:@108438.6]
  assign _T_2152 = _T_2149 + 64'h1; // @[DRAMArbiter.scala 123:18:@108439.6]
  assign _GEN_14 = _T_2146 ? _T_2152 : _T_2149; // @[DRAMArbiter.scala 122:19:@108437.4]
  assign _T_2154 = io_dram_wresp_valid == 1'h0; // @[DRAMArbiter.scala 169:34:@108443.4]
  assign _T_2155 = _T_2154 & io_dram_wresp_ready; // @[DRAMArbiter.scala 169:55:@108444.4]
  assign _T_2160 = _T_2158 + 64'h1; // @[DRAMArbiter.scala 123:18:@108447.6]
  assign _T_2161 = _T_2158 + 64'h1; // @[DRAMArbiter.scala 123:18:@108448.6]
  assign _GEN_15 = _T_2155 ? _T_2161 : _T_2158; // @[DRAMArbiter.scala 122:19:@108446.4]
  assign _T_2168 = io_dram_wresp_bits_tag[7:0]; // @[FringeBundles.scala 140:28:@108456.4]
  assign _T_2172 = _T_2168 == 8'h1; // @[DRAMArbiter.scala 172:116:@108462.4]
  assign _T_2173 = _T_2137 & _T_2172; // @[DRAMArbiter.scala 172:78:@108463.4]
  assign _T_2178 = _T_2176 + 64'h1; // @[DRAMArbiter.scala 123:18:@108466.6]
  assign _T_2179 = _T_2176 + 64'h1; // @[DRAMArbiter.scala 123:18:@108467.6]
  assign _GEN_16 = _T_2173 ? _T_2179 : _T_2176; // @[DRAMArbiter.scala 122:19:@108465.4]
  assign _T_2180 = io_dram_cmd_valid & io_dram_cmd_ready; // @[DRAMArbiter.scala 176:70:@108471.4]
  assign _GEN_17 = _T_2180 ? io_dram_cmd_bits_addr : _T_2182; // @[DRAMArbiter.scala 130:19:@108473.4]
  assign _GEN_18 = _T_2180 ? io_dram_cmd_bits_size : _T_2185; // @[DRAMArbiter.scala 130:19:@108479.4]
  assign _GEN_19 = _T_2039 ? io_dram_wdata_bits_wdata_0 : _T_2188; // @[DRAMArbiter.scala 130:19:@108485.4]
  assign _GEN_20 = _T_2039 ? io_dram_wdata_bits_wstrb_0 : _T_2191; // @[DRAMArbiter.scala 130:19:@108491.4]
  assign _T_2194 = _T_2042 == 64'h0; // @[DRAMArbiter.scala 180:115:@108496.4]
  assign _T_2195 = _T_2039 & _T_2194; // @[DRAMArbiter.scala 180:102:@108497.4]
  assign _GEN_21 = _T_2195 ? io_dram_wdata_bits_wdata_0 : _T_2197; // @[DRAMArbiter.scala 130:19:@108499.4]
  assign _GEN_22 = _T_2195 ? io_dram_wdata_bits_wstrb_0 : _T_2203; // @[DRAMArbiter.scala 130:19:@108507.4]
  assign _T_2206 = _T_2042 == 64'h1; // @[DRAMArbiter.scala 182:115:@108512.4]
  assign _T_2207 = _T_2039 & _T_2206; // @[DRAMArbiter.scala 182:102:@108513.4]
  assign _GEN_23 = _T_2207 ? io_dram_wdata_bits_wdata_0 : _T_2209; // @[DRAMArbiter.scala 130:19:@108515.4]
  assign _GEN_24 = _T_2207 ? io_dram_wdata_bits_wstrb_0 : _T_2215; // @[DRAMArbiter.scala 130:19:@108523.4]
  assign _T_2216 = io_app_stores_0_cmd_valid & io_app_stores_0_cmd_ready; // @[DRAMArbiter.scala 184:92:@108527.4]
  assign _GEN_25 = _T_2216 ? io_app_stores_0_cmd_bits_addr : _T_2218; // @[DRAMArbiter.scala 130:19:@108529.4]
  assign _GEN_26 = _T_2216 ? io_app_stores_0_cmd_bits_size : _T_2221; // @[DRAMArbiter.scala 130:19:@108535.4]
  assign _GEN_27 = _T_2046 ? io_app_stores_0_data_bits_wdata_0 : _T_2224; // @[DRAMArbiter.scala 130:19:@108541.4]
  assign _GEN_28 = _T_2046 ? io_app_stores_0_data_bits_wstrb : _T_2227; // @[DRAMArbiter.scala 130:19:@108547.4]
  assign _T_2230 = _T_2049 == 64'h0; // @[DRAMArbiter.scala 188:148:@108552.4]
  assign _T_2231 = _T_2046 & _T_2230; // @[DRAMArbiter.scala 188:132:@108553.4]
  assign _GEN_29 = _T_2231 ? io_app_stores_0_data_bits_wdata_0 : _T_2233; // @[DRAMArbiter.scala 130:19:@108555.4]
  assign _GEN_30 = _T_2231 ? io_app_stores_0_data_bits_wstrb : _T_2239; // @[DRAMArbiter.scala 130:19:@108563.4]
  assign _T_2242 = _T_2049 == 64'h1; // @[DRAMArbiter.scala 190:148:@108568.4]
  assign _T_2243 = _T_2046 & _T_2242; // @[DRAMArbiter.scala 190:132:@108569.4]
  assign _GEN_31 = _T_2243 ? io_app_stores_0_data_bits_wdata_0 : _T_2245; // @[DRAMArbiter.scala 130:19:@108571.4]
  assign _GEN_32 = _T_2243 ? io_app_stores_0_data_bits_wstrb : _T_2251; // @[DRAMArbiter.scala 130:19:@108579.4]
  assign _T_2325 = _T_2323 + 64'h1; // @[DRAMArbiter.scala 123:18:@108662.6]
  assign _T_2326 = _T_2323 + 64'h1; // @[DRAMArbiter.scala 123:18:@108663.6]
  assign io_app_loads_0_cmd_ready = StreamControllerLoad_io_load_cmd_ready; // @[DRAMArbiter.scala 61:17:@106822.4]
  assign io_app_loads_0_data_valid = StreamControllerLoad_io_load_data_valid; // @[DRAMArbiter.scala 61:17:@106817.4]
  assign io_app_loads_0_data_bits_rdata_0 = StreamControllerLoad_io_load_data_bits_rdata_0; // @[DRAMArbiter.scala 61:17:@106816.4]
  assign io_app_stores_0_cmd_ready = StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 68:18:@106836.4]
  assign io_app_stores_0_data_ready = StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 68:18:@106832.4]
  assign io_app_stores_0_wresp_valid = StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 68:18:@106827.4]
  assign io_app_stores_0_wresp_bits = StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 68:18:@106826.4]
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@108301.4 DRAMArbiter.scala 100:23:@108304.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@108300.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@108299.4]
  assign io_dram_cmd_bits_rawAddr = AXICmdIssue_io_out_cmd_bits_rawAddr; // @[DRAMArbiter.scala 99:13:@108298.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@108297.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@108296.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@108294.4 DRAMArbiter.scala 101:25:@108306.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@108230.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@108231.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@108232.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@108233.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@108234.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@108235.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@108236.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@108237.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@108238.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@108239.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@108240.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@108241.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@108242.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@108243.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@108244.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@108245.4]
  assign io_dram_wdata_bits_wdata_16 = AXICmdIssue_io_out_wdata_bits_wdata_16; // @[DRAMArbiter.scala 99:13:@108246.4]
  assign io_dram_wdata_bits_wdata_17 = AXICmdIssue_io_out_wdata_bits_wdata_17; // @[DRAMArbiter.scala 99:13:@108247.4]
  assign io_dram_wdata_bits_wdata_18 = AXICmdIssue_io_out_wdata_bits_wdata_18; // @[DRAMArbiter.scala 99:13:@108248.4]
  assign io_dram_wdata_bits_wdata_19 = AXICmdIssue_io_out_wdata_bits_wdata_19; // @[DRAMArbiter.scala 99:13:@108249.4]
  assign io_dram_wdata_bits_wdata_20 = AXICmdIssue_io_out_wdata_bits_wdata_20; // @[DRAMArbiter.scala 99:13:@108250.4]
  assign io_dram_wdata_bits_wdata_21 = AXICmdIssue_io_out_wdata_bits_wdata_21; // @[DRAMArbiter.scala 99:13:@108251.4]
  assign io_dram_wdata_bits_wdata_22 = AXICmdIssue_io_out_wdata_bits_wdata_22; // @[DRAMArbiter.scala 99:13:@108252.4]
  assign io_dram_wdata_bits_wdata_23 = AXICmdIssue_io_out_wdata_bits_wdata_23; // @[DRAMArbiter.scala 99:13:@108253.4]
  assign io_dram_wdata_bits_wdata_24 = AXICmdIssue_io_out_wdata_bits_wdata_24; // @[DRAMArbiter.scala 99:13:@108254.4]
  assign io_dram_wdata_bits_wdata_25 = AXICmdIssue_io_out_wdata_bits_wdata_25; // @[DRAMArbiter.scala 99:13:@108255.4]
  assign io_dram_wdata_bits_wdata_26 = AXICmdIssue_io_out_wdata_bits_wdata_26; // @[DRAMArbiter.scala 99:13:@108256.4]
  assign io_dram_wdata_bits_wdata_27 = AXICmdIssue_io_out_wdata_bits_wdata_27; // @[DRAMArbiter.scala 99:13:@108257.4]
  assign io_dram_wdata_bits_wdata_28 = AXICmdIssue_io_out_wdata_bits_wdata_28; // @[DRAMArbiter.scala 99:13:@108258.4]
  assign io_dram_wdata_bits_wdata_29 = AXICmdIssue_io_out_wdata_bits_wdata_29; // @[DRAMArbiter.scala 99:13:@108259.4]
  assign io_dram_wdata_bits_wdata_30 = AXICmdIssue_io_out_wdata_bits_wdata_30; // @[DRAMArbiter.scala 99:13:@108260.4]
  assign io_dram_wdata_bits_wdata_31 = AXICmdIssue_io_out_wdata_bits_wdata_31; // @[DRAMArbiter.scala 99:13:@108261.4]
  assign io_dram_wdata_bits_wdata_32 = AXICmdIssue_io_out_wdata_bits_wdata_32; // @[DRAMArbiter.scala 99:13:@108262.4]
  assign io_dram_wdata_bits_wdata_33 = AXICmdIssue_io_out_wdata_bits_wdata_33; // @[DRAMArbiter.scala 99:13:@108263.4]
  assign io_dram_wdata_bits_wdata_34 = AXICmdIssue_io_out_wdata_bits_wdata_34; // @[DRAMArbiter.scala 99:13:@108264.4]
  assign io_dram_wdata_bits_wdata_35 = AXICmdIssue_io_out_wdata_bits_wdata_35; // @[DRAMArbiter.scala 99:13:@108265.4]
  assign io_dram_wdata_bits_wdata_36 = AXICmdIssue_io_out_wdata_bits_wdata_36; // @[DRAMArbiter.scala 99:13:@108266.4]
  assign io_dram_wdata_bits_wdata_37 = AXICmdIssue_io_out_wdata_bits_wdata_37; // @[DRAMArbiter.scala 99:13:@108267.4]
  assign io_dram_wdata_bits_wdata_38 = AXICmdIssue_io_out_wdata_bits_wdata_38; // @[DRAMArbiter.scala 99:13:@108268.4]
  assign io_dram_wdata_bits_wdata_39 = AXICmdIssue_io_out_wdata_bits_wdata_39; // @[DRAMArbiter.scala 99:13:@108269.4]
  assign io_dram_wdata_bits_wdata_40 = AXICmdIssue_io_out_wdata_bits_wdata_40; // @[DRAMArbiter.scala 99:13:@108270.4]
  assign io_dram_wdata_bits_wdata_41 = AXICmdIssue_io_out_wdata_bits_wdata_41; // @[DRAMArbiter.scala 99:13:@108271.4]
  assign io_dram_wdata_bits_wdata_42 = AXICmdIssue_io_out_wdata_bits_wdata_42; // @[DRAMArbiter.scala 99:13:@108272.4]
  assign io_dram_wdata_bits_wdata_43 = AXICmdIssue_io_out_wdata_bits_wdata_43; // @[DRAMArbiter.scala 99:13:@108273.4]
  assign io_dram_wdata_bits_wdata_44 = AXICmdIssue_io_out_wdata_bits_wdata_44; // @[DRAMArbiter.scala 99:13:@108274.4]
  assign io_dram_wdata_bits_wdata_45 = AXICmdIssue_io_out_wdata_bits_wdata_45; // @[DRAMArbiter.scala 99:13:@108275.4]
  assign io_dram_wdata_bits_wdata_46 = AXICmdIssue_io_out_wdata_bits_wdata_46; // @[DRAMArbiter.scala 99:13:@108276.4]
  assign io_dram_wdata_bits_wdata_47 = AXICmdIssue_io_out_wdata_bits_wdata_47; // @[DRAMArbiter.scala 99:13:@108277.4]
  assign io_dram_wdata_bits_wdata_48 = AXICmdIssue_io_out_wdata_bits_wdata_48; // @[DRAMArbiter.scala 99:13:@108278.4]
  assign io_dram_wdata_bits_wdata_49 = AXICmdIssue_io_out_wdata_bits_wdata_49; // @[DRAMArbiter.scala 99:13:@108279.4]
  assign io_dram_wdata_bits_wdata_50 = AXICmdIssue_io_out_wdata_bits_wdata_50; // @[DRAMArbiter.scala 99:13:@108280.4]
  assign io_dram_wdata_bits_wdata_51 = AXICmdIssue_io_out_wdata_bits_wdata_51; // @[DRAMArbiter.scala 99:13:@108281.4]
  assign io_dram_wdata_bits_wdata_52 = AXICmdIssue_io_out_wdata_bits_wdata_52; // @[DRAMArbiter.scala 99:13:@108282.4]
  assign io_dram_wdata_bits_wdata_53 = AXICmdIssue_io_out_wdata_bits_wdata_53; // @[DRAMArbiter.scala 99:13:@108283.4]
  assign io_dram_wdata_bits_wdata_54 = AXICmdIssue_io_out_wdata_bits_wdata_54; // @[DRAMArbiter.scala 99:13:@108284.4]
  assign io_dram_wdata_bits_wdata_55 = AXICmdIssue_io_out_wdata_bits_wdata_55; // @[DRAMArbiter.scala 99:13:@108285.4]
  assign io_dram_wdata_bits_wdata_56 = AXICmdIssue_io_out_wdata_bits_wdata_56; // @[DRAMArbiter.scala 99:13:@108286.4]
  assign io_dram_wdata_bits_wdata_57 = AXICmdIssue_io_out_wdata_bits_wdata_57; // @[DRAMArbiter.scala 99:13:@108287.4]
  assign io_dram_wdata_bits_wdata_58 = AXICmdIssue_io_out_wdata_bits_wdata_58; // @[DRAMArbiter.scala 99:13:@108288.4]
  assign io_dram_wdata_bits_wdata_59 = AXICmdIssue_io_out_wdata_bits_wdata_59; // @[DRAMArbiter.scala 99:13:@108289.4]
  assign io_dram_wdata_bits_wdata_60 = AXICmdIssue_io_out_wdata_bits_wdata_60; // @[DRAMArbiter.scala 99:13:@108290.4]
  assign io_dram_wdata_bits_wdata_61 = AXICmdIssue_io_out_wdata_bits_wdata_61; // @[DRAMArbiter.scala 99:13:@108291.4]
  assign io_dram_wdata_bits_wdata_62 = AXICmdIssue_io_out_wdata_bits_wdata_62; // @[DRAMArbiter.scala 99:13:@108292.4]
  assign io_dram_wdata_bits_wdata_63 = AXICmdIssue_io_out_wdata_bits_wdata_63; // @[DRAMArbiter.scala 99:13:@108293.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@108166.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@108167.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@108168.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@108169.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@108170.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@108171.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@108172.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@108173.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@108174.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@108175.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@108176.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@108177.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@108178.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@108179.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@108180.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@108181.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@108182.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@108183.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@108184.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@108185.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@108186.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@108187.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@108188.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@108189.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@108190.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@108191.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@108192.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@108193.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@108194.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@108195.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@108196.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@108197.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@108198.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@108199.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@108200.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@108201.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@108202.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@108203.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@108204.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@108205.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@108206.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@108207.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@108208.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@108209.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@108210.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@108211.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@108212.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@108213.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@108214.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@108215.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@108216.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@108217.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@108218.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@108219.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@108220.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@108221.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@108222.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@108223.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@108224.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@108225.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@108226.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@108227.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@108228.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@108229.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@108165.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@108164.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@108097.4]
  assign io_debugSignals_0 = _T_2028[31:0]; // @[DRAMArbiter.scala 111:39:@108313.4]
  assign io_debugSignals_1 = _T_2042[31:0]; // @[DRAMArbiter.scala 111:39:@108335.4]
  assign io_debugSignals_2 = _T_2056[31:0]; // @[DRAMArbiter.scala 111:39:@108343.4]
  assign io_debugSignals_3 = _T_2066[31:0]; // @[DRAMArbiter.scala 111:39:@108353.4]
  assign io_debugSignals_4 = _T_2074[31:0]; // @[DRAMArbiter.scala 111:39:@108362.4]
  assign io_debugSignals_5 = _T_2082[31:0]; // @[DRAMArbiter.scala 111:39:@108371.4]
  assign io_debugSignals_6 = _T_2090[31:0]; // @[DRAMArbiter.scala 111:39:@108380.4]
  assign io_debugSignals_7 = _T_2097[31:0]; // @[DRAMArbiter.scala 111:39:@108388.4]
  assign io_debugSignals_8 = _T_2106[31:0]; // @[DRAMArbiter.scala 111:39:@108397.4]
  assign io_debugSignals_9 = _T_2115[31:0]; // @[DRAMArbiter.scala 111:39:@108406.4]
  assign io_debugSignals_10 = _T_2133[31:0]; // @[DRAMArbiter.scala 111:39:@108425.4]
  assign io_debugSignals_11 = _T_2140[31:0]; // @[DRAMArbiter.scala 111:39:@108433.4]
  assign io_debugSignals_12 = _T_2149[31:0]; // @[DRAMArbiter.scala 111:39:@108442.4]
  assign io_debugSignals_13 = _T_2158[31:0]; // @[DRAMArbiter.scala 111:39:@108451.4]
  assign io_debugSignals_14 = _T_2176[31:0]; // @[DRAMArbiter.scala 111:39:@108470.4]
  assign io_debugSignals_15 = _T_2182[31:0]; // @[DRAMArbiter.scala 111:39:@108476.4]
  assign io_debugSignals_16 = _T_2185; // @[DRAMArbiter.scala 111:39:@108482.4]
  assign io_debugSignals_17 = {{24'd0}, _T_2188}; // @[DRAMArbiter.scala 111:39:@108488.4]
  assign io_debugSignals_18 = {{31'd0}, _T_2191}; // @[DRAMArbiter.scala 111:39:@108494.4]
  assign io_debugSignals_19 = {{24'd0}, _T_2197}; // @[DRAMArbiter.scala 111:39:@108502.4]
  assign io_debugSignals_20 = {{31'd0}, _T_2203}; // @[DRAMArbiter.scala 111:39:@108510.4]
  assign io_debugSignals_21 = {{24'd0}, _T_2209}; // @[DRAMArbiter.scala 111:39:@108518.4]
  assign io_debugSignals_22 = {{31'd0}, _T_2215}; // @[DRAMArbiter.scala 111:39:@108526.4]
  assign io_debugSignals_23 = _T_2218[31:0]; // @[DRAMArbiter.scala 111:39:@108532.4]
  assign io_debugSignals_24 = _T_2221; // @[DRAMArbiter.scala 111:39:@108538.4]
  assign io_debugSignals_25 = _T_2224; // @[DRAMArbiter.scala 111:39:@108544.4]
  assign io_debugSignals_26 = {{31'd0}, _T_2227}; // @[DRAMArbiter.scala 111:39:@108550.4]
  assign io_debugSignals_27 = _T_2233; // @[DRAMArbiter.scala 111:39:@108558.4]
  assign io_debugSignals_28 = {{31'd0}, _T_2239}; // @[DRAMArbiter.scala 111:39:@108566.4]
  assign io_debugSignals_29 = _T_2245; // @[DRAMArbiter.scala 111:39:@108574.4]
  assign io_debugSignals_30 = {{31'd0}, _T_2251}; // @[DRAMArbiter.scala 111:39:@108582.4]
  assign io_debugSignals_41 = _T_2323[31:0]; // @[DRAMArbiter.scala 111:39:@108666.4]
  assign StreamControllerLoad_clock = clock; // @[:@106814.4]
  assign StreamControllerLoad_reset = reset; // @[:@106815.4]
  assign StreamControllerLoad_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@107048.4]
  assign StreamControllerLoad_io_dram_rresp_valid = StreamArbiter_io_app_0_rresp_valid; // @[DRAMArbiter.scala 87:32:@106909.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_0 = StreamArbiter_io_app_0_rresp_bits_rdata_0; // @[DRAMArbiter.scala 87:32:@106845.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_1 = StreamArbiter_io_app_0_rresp_bits_rdata_1; // @[DRAMArbiter.scala 87:32:@106846.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_2 = StreamArbiter_io_app_0_rresp_bits_rdata_2; // @[DRAMArbiter.scala 87:32:@106847.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_3 = StreamArbiter_io_app_0_rresp_bits_rdata_3; // @[DRAMArbiter.scala 87:32:@106848.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_4 = StreamArbiter_io_app_0_rresp_bits_rdata_4; // @[DRAMArbiter.scala 87:32:@106849.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_5 = StreamArbiter_io_app_0_rresp_bits_rdata_5; // @[DRAMArbiter.scala 87:32:@106850.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_6 = StreamArbiter_io_app_0_rresp_bits_rdata_6; // @[DRAMArbiter.scala 87:32:@106851.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_7 = StreamArbiter_io_app_0_rresp_bits_rdata_7; // @[DRAMArbiter.scala 87:32:@106852.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_8 = StreamArbiter_io_app_0_rresp_bits_rdata_8; // @[DRAMArbiter.scala 87:32:@106853.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_9 = StreamArbiter_io_app_0_rresp_bits_rdata_9; // @[DRAMArbiter.scala 87:32:@106854.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_10 = StreamArbiter_io_app_0_rresp_bits_rdata_10; // @[DRAMArbiter.scala 87:32:@106855.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_11 = StreamArbiter_io_app_0_rresp_bits_rdata_11; // @[DRAMArbiter.scala 87:32:@106856.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_12 = StreamArbiter_io_app_0_rresp_bits_rdata_12; // @[DRAMArbiter.scala 87:32:@106857.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_13 = StreamArbiter_io_app_0_rresp_bits_rdata_13; // @[DRAMArbiter.scala 87:32:@106858.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_14 = StreamArbiter_io_app_0_rresp_bits_rdata_14; // @[DRAMArbiter.scala 87:32:@106859.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_15 = StreamArbiter_io_app_0_rresp_bits_rdata_15; // @[DRAMArbiter.scala 87:32:@106860.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_16 = StreamArbiter_io_app_0_rresp_bits_rdata_16; // @[DRAMArbiter.scala 87:32:@106861.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_17 = StreamArbiter_io_app_0_rresp_bits_rdata_17; // @[DRAMArbiter.scala 87:32:@106862.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_18 = StreamArbiter_io_app_0_rresp_bits_rdata_18; // @[DRAMArbiter.scala 87:32:@106863.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_19 = StreamArbiter_io_app_0_rresp_bits_rdata_19; // @[DRAMArbiter.scala 87:32:@106864.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_20 = StreamArbiter_io_app_0_rresp_bits_rdata_20; // @[DRAMArbiter.scala 87:32:@106865.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_21 = StreamArbiter_io_app_0_rresp_bits_rdata_21; // @[DRAMArbiter.scala 87:32:@106866.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_22 = StreamArbiter_io_app_0_rresp_bits_rdata_22; // @[DRAMArbiter.scala 87:32:@106867.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_23 = StreamArbiter_io_app_0_rresp_bits_rdata_23; // @[DRAMArbiter.scala 87:32:@106868.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_24 = StreamArbiter_io_app_0_rresp_bits_rdata_24; // @[DRAMArbiter.scala 87:32:@106869.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_25 = StreamArbiter_io_app_0_rresp_bits_rdata_25; // @[DRAMArbiter.scala 87:32:@106870.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_26 = StreamArbiter_io_app_0_rresp_bits_rdata_26; // @[DRAMArbiter.scala 87:32:@106871.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_27 = StreamArbiter_io_app_0_rresp_bits_rdata_27; // @[DRAMArbiter.scala 87:32:@106872.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_28 = StreamArbiter_io_app_0_rresp_bits_rdata_28; // @[DRAMArbiter.scala 87:32:@106873.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_29 = StreamArbiter_io_app_0_rresp_bits_rdata_29; // @[DRAMArbiter.scala 87:32:@106874.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_30 = StreamArbiter_io_app_0_rresp_bits_rdata_30; // @[DRAMArbiter.scala 87:32:@106875.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_31 = StreamArbiter_io_app_0_rresp_bits_rdata_31; // @[DRAMArbiter.scala 87:32:@106876.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_32 = StreamArbiter_io_app_0_rresp_bits_rdata_32; // @[DRAMArbiter.scala 87:32:@106877.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_33 = StreamArbiter_io_app_0_rresp_bits_rdata_33; // @[DRAMArbiter.scala 87:32:@106878.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_34 = StreamArbiter_io_app_0_rresp_bits_rdata_34; // @[DRAMArbiter.scala 87:32:@106879.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_35 = StreamArbiter_io_app_0_rresp_bits_rdata_35; // @[DRAMArbiter.scala 87:32:@106880.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_36 = StreamArbiter_io_app_0_rresp_bits_rdata_36; // @[DRAMArbiter.scala 87:32:@106881.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_37 = StreamArbiter_io_app_0_rresp_bits_rdata_37; // @[DRAMArbiter.scala 87:32:@106882.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_38 = StreamArbiter_io_app_0_rresp_bits_rdata_38; // @[DRAMArbiter.scala 87:32:@106883.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_39 = StreamArbiter_io_app_0_rresp_bits_rdata_39; // @[DRAMArbiter.scala 87:32:@106884.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_40 = StreamArbiter_io_app_0_rresp_bits_rdata_40; // @[DRAMArbiter.scala 87:32:@106885.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_41 = StreamArbiter_io_app_0_rresp_bits_rdata_41; // @[DRAMArbiter.scala 87:32:@106886.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_42 = StreamArbiter_io_app_0_rresp_bits_rdata_42; // @[DRAMArbiter.scala 87:32:@106887.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_43 = StreamArbiter_io_app_0_rresp_bits_rdata_43; // @[DRAMArbiter.scala 87:32:@106888.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_44 = StreamArbiter_io_app_0_rresp_bits_rdata_44; // @[DRAMArbiter.scala 87:32:@106889.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_45 = StreamArbiter_io_app_0_rresp_bits_rdata_45; // @[DRAMArbiter.scala 87:32:@106890.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_46 = StreamArbiter_io_app_0_rresp_bits_rdata_46; // @[DRAMArbiter.scala 87:32:@106891.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_47 = StreamArbiter_io_app_0_rresp_bits_rdata_47; // @[DRAMArbiter.scala 87:32:@106892.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_48 = StreamArbiter_io_app_0_rresp_bits_rdata_48; // @[DRAMArbiter.scala 87:32:@106893.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_49 = StreamArbiter_io_app_0_rresp_bits_rdata_49; // @[DRAMArbiter.scala 87:32:@106894.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_50 = StreamArbiter_io_app_0_rresp_bits_rdata_50; // @[DRAMArbiter.scala 87:32:@106895.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_51 = StreamArbiter_io_app_0_rresp_bits_rdata_51; // @[DRAMArbiter.scala 87:32:@106896.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_52 = StreamArbiter_io_app_0_rresp_bits_rdata_52; // @[DRAMArbiter.scala 87:32:@106897.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_53 = StreamArbiter_io_app_0_rresp_bits_rdata_53; // @[DRAMArbiter.scala 87:32:@106898.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_54 = StreamArbiter_io_app_0_rresp_bits_rdata_54; // @[DRAMArbiter.scala 87:32:@106899.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_55 = StreamArbiter_io_app_0_rresp_bits_rdata_55; // @[DRAMArbiter.scala 87:32:@106900.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_56 = StreamArbiter_io_app_0_rresp_bits_rdata_56; // @[DRAMArbiter.scala 87:32:@106901.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_57 = StreamArbiter_io_app_0_rresp_bits_rdata_57; // @[DRAMArbiter.scala 87:32:@106902.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_58 = StreamArbiter_io_app_0_rresp_bits_rdata_58; // @[DRAMArbiter.scala 87:32:@106903.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_59 = StreamArbiter_io_app_0_rresp_bits_rdata_59; // @[DRAMArbiter.scala 87:32:@106904.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_60 = StreamArbiter_io_app_0_rresp_bits_rdata_60; // @[DRAMArbiter.scala 87:32:@106905.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_61 = StreamArbiter_io_app_0_rresp_bits_rdata_61; // @[DRAMArbiter.scala 87:32:@106906.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_62 = StreamArbiter_io_app_0_rresp_bits_rdata_62; // @[DRAMArbiter.scala 87:32:@106907.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_63 = StreamArbiter_io_app_0_rresp_bits_rdata_63; // @[DRAMArbiter.scala 87:32:@106908.4]
  assign StreamControllerLoad_io_load_cmd_valid = io_app_loads_0_cmd_valid; // @[DRAMArbiter.scala 61:17:@106821.4]
  assign StreamControllerLoad_io_load_cmd_bits_addr = io_app_loads_0_cmd_bits_addr; // @[DRAMArbiter.scala 61:17:@106820.4]
  assign StreamControllerLoad_io_load_cmd_bits_size = io_app_loads_0_cmd_bits_size; // @[DRAMArbiter.scala 61:17:@106819.4]
  assign StreamControllerLoad_io_load_data_ready = io_app_loads_0_data_ready; // @[DRAMArbiter.scala 61:17:@106818.4]
  assign StreamControllerStore_clock = clock; // @[:@106824.4]
  assign StreamControllerStore_reset = reset; // @[:@106825.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_1_cmd_ready; // @[DRAMArbiter.scala 87:32:@107256.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_1_wdata_ready; // @[DRAMArbiter.scala 87:32:@107249.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_1_wresp_valid; // @[DRAMArbiter.scala 87:32:@107050.4]
  assign StreamControllerStore_io_store_cmd_valid = io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 68:18:@106835.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = io_app_stores_0_cmd_bits_addr; // @[DRAMArbiter.scala 68:18:@106834.4]
  assign StreamControllerStore_io_store_cmd_bits_size = io_app_stores_0_cmd_bits_size; // @[DRAMArbiter.scala 68:18:@106833.4]
  assign StreamControllerStore_io_store_data_valid = io_app_stores_0_data_valid; // @[DRAMArbiter.scala 68:18:@106831.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = io_app_stores_0_data_bits_wdata_0; // @[DRAMArbiter.scala 68:18:@106830.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = io_app_stores_0_data_bits_wstrb; // @[DRAMArbiter.scala 68:18:@106829.4]
  assign StreamControllerStore_io_store_wresp_ready = io_app_stores_0_wresp_ready; // @[DRAMArbiter.scala 68:18:@106828.4]
  assign StreamArbiter_clock = clock; // @[:@106838.4]
  assign StreamArbiter_reset = reset; // @[:@106839.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerLoad_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@107463.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerLoad_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@107462.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerLoad_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@107461.4]
  assign StreamArbiter_io_app_0_rresp_ready = StreamControllerLoad_io_dram_rresp_ready; // @[DRAMArbiter.scala 87:22:@107326.4]
  assign StreamArbiter_io_app_1_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@107671.4]
  assign StreamArbiter_io_app_1_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@107670.4]
  assign StreamArbiter_io_app_1_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@107669.4]
  assign StreamArbiter_io_app_1_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@107664.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@107600.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@107601.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@107602.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@107603.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@107604.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@107605.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@107606.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@107607.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@107608.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@107609.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@107610.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@107611.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@107612.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@107613.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@107614.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@107615.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_16 = StreamControllerStore_io_dram_wdata_bits_wdata_16; // @[DRAMArbiter.scala 87:22:@107616.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_17 = StreamControllerStore_io_dram_wdata_bits_wdata_17; // @[DRAMArbiter.scala 87:22:@107617.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_18 = StreamControllerStore_io_dram_wdata_bits_wdata_18; // @[DRAMArbiter.scala 87:22:@107618.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_19 = StreamControllerStore_io_dram_wdata_bits_wdata_19; // @[DRAMArbiter.scala 87:22:@107619.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_20 = StreamControllerStore_io_dram_wdata_bits_wdata_20; // @[DRAMArbiter.scala 87:22:@107620.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_21 = StreamControllerStore_io_dram_wdata_bits_wdata_21; // @[DRAMArbiter.scala 87:22:@107621.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_22 = StreamControllerStore_io_dram_wdata_bits_wdata_22; // @[DRAMArbiter.scala 87:22:@107622.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_23 = StreamControllerStore_io_dram_wdata_bits_wdata_23; // @[DRAMArbiter.scala 87:22:@107623.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_24 = StreamControllerStore_io_dram_wdata_bits_wdata_24; // @[DRAMArbiter.scala 87:22:@107624.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_25 = StreamControllerStore_io_dram_wdata_bits_wdata_25; // @[DRAMArbiter.scala 87:22:@107625.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_26 = StreamControllerStore_io_dram_wdata_bits_wdata_26; // @[DRAMArbiter.scala 87:22:@107626.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_27 = StreamControllerStore_io_dram_wdata_bits_wdata_27; // @[DRAMArbiter.scala 87:22:@107627.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_28 = StreamControllerStore_io_dram_wdata_bits_wdata_28; // @[DRAMArbiter.scala 87:22:@107628.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_29 = StreamControllerStore_io_dram_wdata_bits_wdata_29; // @[DRAMArbiter.scala 87:22:@107629.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_30 = StreamControllerStore_io_dram_wdata_bits_wdata_30; // @[DRAMArbiter.scala 87:22:@107630.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_31 = StreamControllerStore_io_dram_wdata_bits_wdata_31; // @[DRAMArbiter.scala 87:22:@107631.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_32 = StreamControllerStore_io_dram_wdata_bits_wdata_32; // @[DRAMArbiter.scala 87:22:@107632.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_33 = StreamControllerStore_io_dram_wdata_bits_wdata_33; // @[DRAMArbiter.scala 87:22:@107633.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_34 = StreamControllerStore_io_dram_wdata_bits_wdata_34; // @[DRAMArbiter.scala 87:22:@107634.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_35 = StreamControllerStore_io_dram_wdata_bits_wdata_35; // @[DRAMArbiter.scala 87:22:@107635.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_36 = StreamControllerStore_io_dram_wdata_bits_wdata_36; // @[DRAMArbiter.scala 87:22:@107636.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_37 = StreamControllerStore_io_dram_wdata_bits_wdata_37; // @[DRAMArbiter.scala 87:22:@107637.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_38 = StreamControllerStore_io_dram_wdata_bits_wdata_38; // @[DRAMArbiter.scala 87:22:@107638.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_39 = StreamControllerStore_io_dram_wdata_bits_wdata_39; // @[DRAMArbiter.scala 87:22:@107639.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_40 = StreamControllerStore_io_dram_wdata_bits_wdata_40; // @[DRAMArbiter.scala 87:22:@107640.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_41 = StreamControllerStore_io_dram_wdata_bits_wdata_41; // @[DRAMArbiter.scala 87:22:@107641.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_42 = StreamControllerStore_io_dram_wdata_bits_wdata_42; // @[DRAMArbiter.scala 87:22:@107642.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_43 = StreamControllerStore_io_dram_wdata_bits_wdata_43; // @[DRAMArbiter.scala 87:22:@107643.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_44 = StreamControllerStore_io_dram_wdata_bits_wdata_44; // @[DRAMArbiter.scala 87:22:@107644.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_45 = StreamControllerStore_io_dram_wdata_bits_wdata_45; // @[DRAMArbiter.scala 87:22:@107645.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_46 = StreamControllerStore_io_dram_wdata_bits_wdata_46; // @[DRAMArbiter.scala 87:22:@107646.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_47 = StreamControllerStore_io_dram_wdata_bits_wdata_47; // @[DRAMArbiter.scala 87:22:@107647.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_48 = StreamControllerStore_io_dram_wdata_bits_wdata_48; // @[DRAMArbiter.scala 87:22:@107648.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_49 = StreamControllerStore_io_dram_wdata_bits_wdata_49; // @[DRAMArbiter.scala 87:22:@107649.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_50 = StreamControllerStore_io_dram_wdata_bits_wdata_50; // @[DRAMArbiter.scala 87:22:@107650.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_51 = StreamControllerStore_io_dram_wdata_bits_wdata_51; // @[DRAMArbiter.scala 87:22:@107651.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_52 = StreamControllerStore_io_dram_wdata_bits_wdata_52; // @[DRAMArbiter.scala 87:22:@107652.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_53 = StreamControllerStore_io_dram_wdata_bits_wdata_53; // @[DRAMArbiter.scala 87:22:@107653.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_54 = StreamControllerStore_io_dram_wdata_bits_wdata_54; // @[DRAMArbiter.scala 87:22:@107654.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_55 = StreamControllerStore_io_dram_wdata_bits_wdata_55; // @[DRAMArbiter.scala 87:22:@107655.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_56 = StreamControllerStore_io_dram_wdata_bits_wdata_56; // @[DRAMArbiter.scala 87:22:@107656.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_57 = StreamControllerStore_io_dram_wdata_bits_wdata_57; // @[DRAMArbiter.scala 87:22:@107657.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_58 = StreamControllerStore_io_dram_wdata_bits_wdata_58; // @[DRAMArbiter.scala 87:22:@107658.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_59 = StreamControllerStore_io_dram_wdata_bits_wdata_59; // @[DRAMArbiter.scala 87:22:@107659.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_60 = StreamControllerStore_io_dram_wdata_bits_wdata_60; // @[DRAMArbiter.scala 87:22:@107660.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_61 = StreamControllerStore_io_dram_wdata_bits_wdata_61; // @[DRAMArbiter.scala 87:22:@107661.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_62 = StreamControllerStore_io_dram_wdata_bits_wdata_62; // @[DRAMArbiter.scala 87:22:@107662.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_63 = StreamControllerStore_io_dram_wdata_bits_wdata_63; // @[DRAMArbiter.scala 87:22:@107663.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@107536.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@107537.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@107538.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@107539.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@107540.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@107541.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@107542.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@107543.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@107544.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@107545.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@107546.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@107547.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@107548.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@107549.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@107550.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@107551.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@107552.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@107553.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@107554.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@107555.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@107556.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@107557.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@107558.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@107559.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@107560.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@107561.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@107562.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@107563.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@107564.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@107565.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@107566.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@107567.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@107568.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@107569.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@107570.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@107571.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@107572.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@107573.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@107574.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@107575.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@107576.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@107577.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@107578.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@107579.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@107580.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@107581.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@107582.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@107583.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@107584.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@107585.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@107586.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@107587.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@107588.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@107589.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@107590.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@107591.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@107592.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@107593.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@107594.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@107595.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@107596.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@107597.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@107598.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@107599.4]
  assign StreamArbiter_io_app_1_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@107467.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@107883.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@107876.4]
  assign StreamArbiter_io_dram_rresp_valid = AXICmdSplit_io_in_rresp_valid; // @[DRAMArbiter.scala 95:20:@107744.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_0 = AXICmdSplit_io_in_rresp_bits_rdata_0; // @[DRAMArbiter.scala 95:20:@107680.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_1 = AXICmdSplit_io_in_rresp_bits_rdata_1; // @[DRAMArbiter.scala 95:20:@107681.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_2 = AXICmdSplit_io_in_rresp_bits_rdata_2; // @[DRAMArbiter.scala 95:20:@107682.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_3 = AXICmdSplit_io_in_rresp_bits_rdata_3; // @[DRAMArbiter.scala 95:20:@107683.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_4 = AXICmdSplit_io_in_rresp_bits_rdata_4; // @[DRAMArbiter.scala 95:20:@107684.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_5 = AXICmdSplit_io_in_rresp_bits_rdata_5; // @[DRAMArbiter.scala 95:20:@107685.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_6 = AXICmdSplit_io_in_rresp_bits_rdata_6; // @[DRAMArbiter.scala 95:20:@107686.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_7 = AXICmdSplit_io_in_rresp_bits_rdata_7; // @[DRAMArbiter.scala 95:20:@107687.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_8 = AXICmdSplit_io_in_rresp_bits_rdata_8; // @[DRAMArbiter.scala 95:20:@107688.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_9 = AXICmdSplit_io_in_rresp_bits_rdata_9; // @[DRAMArbiter.scala 95:20:@107689.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_10 = AXICmdSplit_io_in_rresp_bits_rdata_10; // @[DRAMArbiter.scala 95:20:@107690.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_11 = AXICmdSplit_io_in_rresp_bits_rdata_11; // @[DRAMArbiter.scala 95:20:@107691.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_12 = AXICmdSplit_io_in_rresp_bits_rdata_12; // @[DRAMArbiter.scala 95:20:@107692.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_13 = AXICmdSplit_io_in_rresp_bits_rdata_13; // @[DRAMArbiter.scala 95:20:@107693.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_14 = AXICmdSplit_io_in_rresp_bits_rdata_14; // @[DRAMArbiter.scala 95:20:@107694.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_15 = AXICmdSplit_io_in_rresp_bits_rdata_15; // @[DRAMArbiter.scala 95:20:@107695.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_16 = AXICmdSplit_io_in_rresp_bits_rdata_16; // @[DRAMArbiter.scala 95:20:@107696.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_17 = AXICmdSplit_io_in_rresp_bits_rdata_17; // @[DRAMArbiter.scala 95:20:@107697.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_18 = AXICmdSplit_io_in_rresp_bits_rdata_18; // @[DRAMArbiter.scala 95:20:@107698.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_19 = AXICmdSplit_io_in_rresp_bits_rdata_19; // @[DRAMArbiter.scala 95:20:@107699.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_20 = AXICmdSplit_io_in_rresp_bits_rdata_20; // @[DRAMArbiter.scala 95:20:@107700.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_21 = AXICmdSplit_io_in_rresp_bits_rdata_21; // @[DRAMArbiter.scala 95:20:@107701.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_22 = AXICmdSplit_io_in_rresp_bits_rdata_22; // @[DRAMArbiter.scala 95:20:@107702.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_23 = AXICmdSplit_io_in_rresp_bits_rdata_23; // @[DRAMArbiter.scala 95:20:@107703.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_24 = AXICmdSplit_io_in_rresp_bits_rdata_24; // @[DRAMArbiter.scala 95:20:@107704.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_25 = AXICmdSplit_io_in_rresp_bits_rdata_25; // @[DRAMArbiter.scala 95:20:@107705.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_26 = AXICmdSplit_io_in_rresp_bits_rdata_26; // @[DRAMArbiter.scala 95:20:@107706.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_27 = AXICmdSplit_io_in_rresp_bits_rdata_27; // @[DRAMArbiter.scala 95:20:@107707.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_28 = AXICmdSplit_io_in_rresp_bits_rdata_28; // @[DRAMArbiter.scala 95:20:@107708.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_29 = AXICmdSplit_io_in_rresp_bits_rdata_29; // @[DRAMArbiter.scala 95:20:@107709.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_30 = AXICmdSplit_io_in_rresp_bits_rdata_30; // @[DRAMArbiter.scala 95:20:@107710.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_31 = AXICmdSplit_io_in_rresp_bits_rdata_31; // @[DRAMArbiter.scala 95:20:@107711.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_32 = AXICmdSplit_io_in_rresp_bits_rdata_32; // @[DRAMArbiter.scala 95:20:@107712.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_33 = AXICmdSplit_io_in_rresp_bits_rdata_33; // @[DRAMArbiter.scala 95:20:@107713.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_34 = AXICmdSplit_io_in_rresp_bits_rdata_34; // @[DRAMArbiter.scala 95:20:@107714.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_35 = AXICmdSplit_io_in_rresp_bits_rdata_35; // @[DRAMArbiter.scala 95:20:@107715.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_36 = AXICmdSplit_io_in_rresp_bits_rdata_36; // @[DRAMArbiter.scala 95:20:@107716.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_37 = AXICmdSplit_io_in_rresp_bits_rdata_37; // @[DRAMArbiter.scala 95:20:@107717.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_38 = AXICmdSplit_io_in_rresp_bits_rdata_38; // @[DRAMArbiter.scala 95:20:@107718.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_39 = AXICmdSplit_io_in_rresp_bits_rdata_39; // @[DRAMArbiter.scala 95:20:@107719.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_40 = AXICmdSplit_io_in_rresp_bits_rdata_40; // @[DRAMArbiter.scala 95:20:@107720.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_41 = AXICmdSplit_io_in_rresp_bits_rdata_41; // @[DRAMArbiter.scala 95:20:@107721.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_42 = AXICmdSplit_io_in_rresp_bits_rdata_42; // @[DRAMArbiter.scala 95:20:@107722.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_43 = AXICmdSplit_io_in_rresp_bits_rdata_43; // @[DRAMArbiter.scala 95:20:@107723.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_44 = AXICmdSplit_io_in_rresp_bits_rdata_44; // @[DRAMArbiter.scala 95:20:@107724.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_45 = AXICmdSplit_io_in_rresp_bits_rdata_45; // @[DRAMArbiter.scala 95:20:@107725.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_46 = AXICmdSplit_io_in_rresp_bits_rdata_46; // @[DRAMArbiter.scala 95:20:@107726.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_47 = AXICmdSplit_io_in_rresp_bits_rdata_47; // @[DRAMArbiter.scala 95:20:@107727.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_48 = AXICmdSplit_io_in_rresp_bits_rdata_48; // @[DRAMArbiter.scala 95:20:@107728.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_49 = AXICmdSplit_io_in_rresp_bits_rdata_49; // @[DRAMArbiter.scala 95:20:@107729.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_50 = AXICmdSplit_io_in_rresp_bits_rdata_50; // @[DRAMArbiter.scala 95:20:@107730.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_51 = AXICmdSplit_io_in_rresp_bits_rdata_51; // @[DRAMArbiter.scala 95:20:@107731.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_52 = AXICmdSplit_io_in_rresp_bits_rdata_52; // @[DRAMArbiter.scala 95:20:@107732.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_53 = AXICmdSplit_io_in_rresp_bits_rdata_53; // @[DRAMArbiter.scala 95:20:@107733.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_54 = AXICmdSplit_io_in_rresp_bits_rdata_54; // @[DRAMArbiter.scala 95:20:@107734.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_55 = AXICmdSplit_io_in_rresp_bits_rdata_55; // @[DRAMArbiter.scala 95:20:@107735.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_56 = AXICmdSplit_io_in_rresp_bits_rdata_56; // @[DRAMArbiter.scala 95:20:@107736.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_57 = AXICmdSplit_io_in_rresp_bits_rdata_57; // @[DRAMArbiter.scala 95:20:@107737.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_58 = AXICmdSplit_io_in_rresp_bits_rdata_58; // @[DRAMArbiter.scala 95:20:@107738.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_59 = AXICmdSplit_io_in_rresp_bits_rdata_59; // @[DRAMArbiter.scala 95:20:@107739.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_60 = AXICmdSplit_io_in_rresp_bits_rdata_60; // @[DRAMArbiter.scala 95:20:@107740.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_61 = AXICmdSplit_io_in_rresp_bits_rdata_61; // @[DRAMArbiter.scala 95:20:@107741.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_62 = AXICmdSplit_io_in_rresp_bits_rdata_62; // @[DRAMArbiter.scala 95:20:@107742.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_63 = AXICmdSplit_io_in_rresp_bits_rdata_63; // @[DRAMArbiter.scala 95:20:@107743.4]
  assign StreamArbiter_io_dram_rresp_bits_tag = AXICmdSplit_io_in_rresp_bits_tag; // @[DRAMArbiter.scala 95:20:@107679.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@107677.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@107676.4]
  assign AXICmdSplit_clock = clock; // @[:@107674.4]
  assign AXICmdSplit_reset = reset; // @[:@107675.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@107882.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@107881.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@107880.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@107878.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@107877.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@107875.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@107811.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@107812.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@107813.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@107814.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@107815.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@107816.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@107817.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@107818.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@107819.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@107820.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@107821.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@107822.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@107823.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@107824.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@107825.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@107826.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_16 = StreamArbiter_io_dram_wdata_bits_wdata_16; // @[DRAMArbiter.scala 95:20:@107827.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_17 = StreamArbiter_io_dram_wdata_bits_wdata_17; // @[DRAMArbiter.scala 95:20:@107828.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_18 = StreamArbiter_io_dram_wdata_bits_wdata_18; // @[DRAMArbiter.scala 95:20:@107829.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_19 = StreamArbiter_io_dram_wdata_bits_wdata_19; // @[DRAMArbiter.scala 95:20:@107830.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_20 = StreamArbiter_io_dram_wdata_bits_wdata_20; // @[DRAMArbiter.scala 95:20:@107831.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_21 = StreamArbiter_io_dram_wdata_bits_wdata_21; // @[DRAMArbiter.scala 95:20:@107832.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_22 = StreamArbiter_io_dram_wdata_bits_wdata_22; // @[DRAMArbiter.scala 95:20:@107833.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_23 = StreamArbiter_io_dram_wdata_bits_wdata_23; // @[DRAMArbiter.scala 95:20:@107834.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_24 = StreamArbiter_io_dram_wdata_bits_wdata_24; // @[DRAMArbiter.scala 95:20:@107835.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_25 = StreamArbiter_io_dram_wdata_bits_wdata_25; // @[DRAMArbiter.scala 95:20:@107836.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_26 = StreamArbiter_io_dram_wdata_bits_wdata_26; // @[DRAMArbiter.scala 95:20:@107837.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_27 = StreamArbiter_io_dram_wdata_bits_wdata_27; // @[DRAMArbiter.scala 95:20:@107838.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_28 = StreamArbiter_io_dram_wdata_bits_wdata_28; // @[DRAMArbiter.scala 95:20:@107839.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_29 = StreamArbiter_io_dram_wdata_bits_wdata_29; // @[DRAMArbiter.scala 95:20:@107840.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_30 = StreamArbiter_io_dram_wdata_bits_wdata_30; // @[DRAMArbiter.scala 95:20:@107841.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_31 = StreamArbiter_io_dram_wdata_bits_wdata_31; // @[DRAMArbiter.scala 95:20:@107842.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_32 = StreamArbiter_io_dram_wdata_bits_wdata_32; // @[DRAMArbiter.scala 95:20:@107843.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_33 = StreamArbiter_io_dram_wdata_bits_wdata_33; // @[DRAMArbiter.scala 95:20:@107844.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_34 = StreamArbiter_io_dram_wdata_bits_wdata_34; // @[DRAMArbiter.scala 95:20:@107845.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_35 = StreamArbiter_io_dram_wdata_bits_wdata_35; // @[DRAMArbiter.scala 95:20:@107846.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_36 = StreamArbiter_io_dram_wdata_bits_wdata_36; // @[DRAMArbiter.scala 95:20:@107847.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_37 = StreamArbiter_io_dram_wdata_bits_wdata_37; // @[DRAMArbiter.scala 95:20:@107848.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_38 = StreamArbiter_io_dram_wdata_bits_wdata_38; // @[DRAMArbiter.scala 95:20:@107849.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_39 = StreamArbiter_io_dram_wdata_bits_wdata_39; // @[DRAMArbiter.scala 95:20:@107850.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_40 = StreamArbiter_io_dram_wdata_bits_wdata_40; // @[DRAMArbiter.scala 95:20:@107851.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_41 = StreamArbiter_io_dram_wdata_bits_wdata_41; // @[DRAMArbiter.scala 95:20:@107852.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_42 = StreamArbiter_io_dram_wdata_bits_wdata_42; // @[DRAMArbiter.scala 95:20:@107853.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_43 = StreamArbiter_io_dram_wdata_bits_wdata_43; // @[DRAMArbiter.scala 95:20:@107854.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_44 = StreamArbiter_io_dram_wdata_bits_wdata_44; // @[DRAMArbiter.scala 95:20:@107855.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_45 = StreamArbiter_io_dram_wdata_bits_wdata_45; // @[DRAMArbiter.scala 95:20:@107856.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_46 = StreamArbiter_io_dram_wdata_bits_wdata_46; // @[DRAMArbiter.scala 95:20:@107857.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_47 = StreamArbiter_io_dram_wdata_bits_wdata_47; // @[DRAMArbiter.scala 95:20:@107858.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_48 = StreamArbiter_io_dram_wdata_bits_wdata_48; // @[DRAMArbiter.scala 95:20:@107859.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_49 = StreamArbiter_io_dram_wdata_bits_wdata_49; // @[DRAMArbiter.scala 95:20:@107860.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_50 = StreamArbiter_io_dram_wdata_bits_wdata_50; // @[DRAMArbiter.scala 95:20:@107861.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_51 = StreamArbiter_io_dram_wdata_bits_wdata_51; // @[DRAMArbiter.scala 95:20:@107862.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_52 = StreamArbiter_io_dram_wdata_bits_wdata_52; // @[DRAMArbiter.scala 95:20:@107863.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_53 = StreamArbiter_io_dram_wdata_bits_wdata_53; // @[DRAMArbiter.scala 95:20:@107864.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_54 = StreamArbiter_io_dram_wdata_bits_wdata_54; // @[DRAMArbiter.scala 95:20:@107865.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_55 = StreamArbiter_io_dram_wdata_bits_wdata_55; // @[DRAMArbiter.scala 95:20:@107866.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_56 = StreamArbiter_io_dram_wdata_bits_wdata_56; // @[DRAMArbiter.scala 95:20:@107867.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_57 = StreamArbiter_io_dram_wdata_bits_wdata_57; // @[DRAMArbiter.scala 95:20:@107868.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_58 = StreamArbiter_io_dram_wdata_bits_wdata_58; // @[DRAMArbiter.scala 95:20:@107869.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_59 = StreamArbiter_io_dram_wdata_bits_wdata_59; // @[DRAMArbiter.scala 95:20:@107870.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_60 = StreamArbiter_io_dram_wdata_bits_wdata_60; // @[DRAMArbiter.scala 95:20:@107871.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_61 = StreamArbiter_io_dram_wdata_bits_wdata_61; // @[DRAMArbiter.scala 95:20:@107872.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_62 = StreamArbiter_io_dram_wdata_bits_wdata_62; // @[DRAMArbiter.scala 95:20:@107873.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_63 = StreamArbiter_io_dram_wdata_bits_wdata_63; // @[DRAMArbiter.scala 95:20:@107874.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@107747.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@107748.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@107749.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@107750.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@107751.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@107752.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@107753.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@107754.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@107755.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@107756.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@107757.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@107758.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@107759.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@107760.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@107761.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@107762.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@107763.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@107764.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@107765.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@107766.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@107767.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@107768.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@107769.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@107770.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@107771.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@107772.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@107773.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@107774.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@107775.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@107776.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@107777.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@107778.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@107779.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@107780.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@107781.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@107782.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@107783.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@107784.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@107785.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@107786.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@107787.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@107788.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@107789.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@107790.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@107791.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@107792.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@107793.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@107794.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@107795.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@107796.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@107797.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@107798.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@107799.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@107800.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@107801.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@107802.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@107803.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@107804.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@107805.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@107806.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@107807.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@107808.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@107809.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@107810.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@107745.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@107678.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@108094.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@108087.4]
  assign AXICmdSplit_io_out_rresp_valid = AXICmdIssue_io_in_rresp_valid; // @[DRAMArbiter.scala 98:20:@107955.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_0 = AXICmdIssue_io_in_rresp_bits_rdata_0; // @[DRAMArbiter.scala 98:20:@107891.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_1 = AXICmdIssue_io_in_rresp_bits_rdata_1; // @[DRAMArbiter.scala 98:20:@107892.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_2 = AXICmdIssue_io_in_rresp_bits_rdata_2; // @[DRAMArbiter.scala 98:20:@107893.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_3 = AXICmdIssue_io_in_rresp_bits_rdata_3; // @[DRAMArbiter.scala 98:20:@107894.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_4 = AXICmdIssue_io_in_rresp_bits_rdata_4; // @[DRAMArbiter.scala 98:20:@107895.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_5 = AXICmdIssue_io_in_rresp_bits_rdata_5; // @[DRAMArbiter.scala 98:20:@107896.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_6 = AXICmdIssue_io_in_rresp_bits_rdata_6; // @[DRAMArbiter.scala 98:20:@107897.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_7 = AXICmdIssue_io_in_rresp_bits_rdata_7; // @[DRAMArbiter.scala 98:20:@107898.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_8 = AXICmdIssue_io_in_rresp_bits_rdata_8; // @[DRAMArbiter.scala 98:20:@107899.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_9 = AXICmdIssue_io_in_rresp_bits_rdata_9; // @[DRAMArbiter.scala 98:20:@107900.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_10 = AXICmdIssue_io_in_rresp_bits_rdata_10; // @[DRAMArbiter.scala 98:20:@107901.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_11 = AXICmdIssue_io_in_rresp_bits_rdata_11; // @[DRAMArbiter.scala 98:20:@107902.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_12 = AXICmdIssue_io_in_rresp_bits_rdata_12; // @[DRAMArbiter.scala 98:20:@107903.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_13 = AXICmdIssue_io_in_rresp_bits_rdata_13; // @[DRAMArbiter.scala 98:20:@107904.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_14 = AXICmdIssue_io_in_rresp_bits_rdata_14; // @[DRAMArbiter.scala 98:20:@107905.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_15 = AXICmdIssue_io_in_rresp_bits_rdata_15; // @[DRAMArbiter.scala 98:20:@107906.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_16 = AXICmdIssue_io_in_rresp_bits_rdata_16; // @[DRAMArbiter.scala 98:20:@107907.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_17 = AXICmdIssue_io_in_rresp_bits_rdata_17; // @[DRAMArbiter.scala 98:20:@107908.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_18 = AXICmdIssue_io_in_rresp_bits_rdata_18; // @[DRAMArbiter.scala 98:20:@107909.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_19 = AXICmdIssue_io_in_rresp_bits_rdata_19; // @[DRAMArbiter.scala 98:20:@107910.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_20 = AXICmdIssue_io_in_rresp_bits_rdata_20; // @[DRAMArbiter.scala 98:20:@107911.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_21 = AXICmdIssue_io_in_rresp_bits_rdata_21; // @[DRAMArbiter.scala 98:20:@107912.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_22 = AXICmdIssue_io_in_rresp_bits_rdata_22; // @[DRAMArbiter.scala 98:20:@107913.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_23 = AXICmdIssue_io_in_rresp_bits_rdata_23; // @[DRAMArbiter.scala 98:20:@107914.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_24 = AXICmdIssue_io_in_rresp_bits_rdata_24; // @[DRAMArbiter.scala 98:20:@107915.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_25 = AXICmdIssue_io_in_rresp_bits_rdata_25; // @[DRAMArbiter.scala 98:20:@107916.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_26 = AXICmdIssue_io_in_rresp_bits_rdata_26; // @[DRAMArbiter.scala 98:20:@107917.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_27 = AXICmdIssue_io_in_rresp_bits_rdata_27; // @[DRAMArbiter.scala 98:20:@107918.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_28 = AXICmdIssue_io_in_rresp_bits_rdata_28; // @[DRAMArbiter.scala 98:20:@107919.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_29 = AXICmdIssue_io_in_rresp_bits_rdata_29; // @[DRAMArbiter.scala 98:20:@107920.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_30 = AXICmdIssue_io_in_rresp_bits_rdata_30; // @[DRAMArbiter.scala 98:20:@107921.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_31 = AXICmdIssue_io_in_rresp_bits_rdata_31; // @[DRAMArbiter.scala 98:20:@107922.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_32 = AXICmdIssue_io_in_rresp_bits_rdata_32; // @[DRAMArbiter.scala 98:20:@107923.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_33 = AXICmdIssue_io_in_rresp_bits_rdata_33; // @[DRAMArbiter.scala 98:20:@107924.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_34 = AXICmdIssue_io_in_rresp_bits_rdata_34; // @[DRAMArbiter.scala 98:20:@107925.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_35 = AXICmdIssue_io_in_rresp_bits_rdata_35; // @[DRAMArbiter.scala 98:20:@107926.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_36 = AXICmdIssue_io_in_rresp_bits_rdata_36; // @[DRAMArbiter.scala 98:20:@107927.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_37 = AXICmdIssue_io_in_rresp_bits_rdata_37; // @[DRAMArbiter.scala 98:20:@107928.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_38 = AXICmdIssue_io_in_rresp_bits_rdata_38; // @[DRAMArbiter.scala 98:20:@107929.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_39 = AXICmdIssue_io_in_rresp_bits_rdata_39; // @[DRAMArbiter.scala 98:20:@107930.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_40 = AXICmdIssue_io_in_rresp_bits_rdata_40; // @[DRAMArbiter.scala 98:20:@107931.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_41 = AXICmdIssue_io_in_rresp_bits_rdata_41; // @[DRAMArbiter.scala 98:20:@107932.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_42 = AXICmdIssue_io_in_rresp_bits_rdata_42; // @[DRAMArbiter.scala 98:20:@107933.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_43 = AXICmdIssue_io_in_rresp_bits_rdata_43; // @[DRAMArbiter.scala 98:20:@107934.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_44 = AXICmdIssue_io_in_rresp_bits_rdata_44; // @[DRAMArbiter.scala 98:20:@107935.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_45 = AXICmdIssue_io_in_rresp_bits_rdata_45; // @[DRAMArbiter.scala 98:20:@107936.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_46 = AXICmdIssue_io_in_rresp_bits_rdata_46; // @[DRAMArbiter.scala 98:20:@107937.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_47 = AXICmdIssue_io_in_rresp_bits_rdata_47; // @[DRAMArbiter.scala 98:20:@107938.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_48 = AXICmdIssue_io_in_rresp_bits_rdata_48; // @[DRAMArbiter.scala 98:20:@107939.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_49 = AXICmdIssue_io_in_rresp_bits_rdata_49; // @[DRAMArbiter.scala 98:20:@107940.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_50 = AXICmdIssue_io_in_rresp_bits_rdata_50; // @[DRAMArbiter.scala 98:20:@107941.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_51 = AXICmdIssue_io_in_rresp_bits_rdata_51; // @[DRAMArbiter.scala 98:20:@107942.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_52 = AXICmdIssue_io_in_rresp_bits_rdata_52; // @[DRAMArbiter.scala 98:20:@107943.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_53 = AXICmdIssue_io_in_rresp_bits_rdata_53; // @[DRAMArbiter.scala 98:20:@107944.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_54 = AXICmdIssue_io_in_rresp_bits_rdata_54; // @[DRAMArbiter.scala 98:20:@107945.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_55 = AXICmdIssue_io_in_rresp_bits_rdata_55; // @[DRAMArbiter.scala 98:20:@107946.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_56 = AXICmdIssue_io_in_rresp_bits_rdata_56; // @[DRAMArbiter.scala 98:20:@107947.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_57 = AXICmdIssue_io_in_rresp_bits_rdata_57; // @[DRAMArbiter.scala 98:20:@107948.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_58 = AXICmdIssue_io_in_rresp_bits_rdata_58; // @[DRAMArbiter.scala 98:20:@107949.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_59 = AXICmdIssue_io_in_rresp_bits_rdata_59; // @[DRAMArbiter.scala 98:20:@107950.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_60 = AXICmdIssue_io_in_rresp_bits_rdata_60; // @[DRAMArbiter.scala 98:20:@107951.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_61 = AXICmdIssue_io_in_rresp_bits_rdata_61; // @[DRAMArbiter.scala 98:20:@107952.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_62 = AXICmdIssue_io_in_rresp_bits_rdata_62; // @[DRAMArbiter.scala 98:20:@107953.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_63 = AXICmdIssue_io_in_rresp_bits_rdata_63; // @[DRAMArbiter.scala 98:20:@107954.4]
  assign AXICmdSplit_io_out_rresp_bits_tag = AXICmdIssue_io_in_rresp_bits_tag; // @[DRAMArbiter.scala 98:20:@107890.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@107888.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@107887.4]
  assign AXICmdIssue_clock = clock; // @[:@107885.4]
  assign AXICmdIssue_reset = reset; // @[:@107886.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@108093.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@108092.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@108091.4]
  assign AXICmdIssue_io_in_cmd_bits_rawAddr = AXICmdSplit_io_out_cmd_bits_rawAddr; // @[DRAMArbiter.scala 98:20:@108090.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@108089.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@108088.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@108086.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@108022.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@108023.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@108024.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@108025.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@108026.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@108027.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@108028.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@108029.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@108030.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@108031.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@108032.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@108033.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@108034.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@108035.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@108036.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@108037.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_16 = AXICmdSplit_io_out_wdata_bits_wdata_16; // @[DRAMArbiter.scala 98:20:@108038.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_17 = AXICmdSplit_io_out_wdata_bits_wdata_17; // @[DRAMArbiter.scala 98:20:@108039.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_18 = AXICmdSplit_io_out_wdata_bits_wdata_18; // @[DRAMArbiter.scala 98:20:@108040.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_19 = AXICmdSplit_io_out_wdata_bits_wdata_19; // @[DRAMArbiter.scala 98:20:@108041.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_20 = AXICmdSplit_io_out_wdata_bits_wdata_20; // @[DRAMArbiter.scala 98:20:@108042.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_21 = AXICmdSplit_io_out_wdata_bits_wdata_21; // @[DRAMArbiter.scala 98:20:@108043.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_22 = AXICmdSplit_io_out_wdata_bits_wdata_22; // @[DRAMArbiter.scala 98:20:@108044.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_23 = AXICmdSplit_io_out_wdata_bits_wdata_23; // @[DRAMArbiter.scala 98:20:@108045.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_24 = AXICmdSplit_io_out_wdata_bits_wdata_24; // @[DRAMArbiter.scala 98:20:@108046.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_25 = AXICmdSplit_io_out_wdata_bits_wdata_25; // @[DRAMArbiter.scala 98:20:@108047.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_26 = AXICmdSplit_io_out_wdata_bits_wdata_26; // @[DRAMArbiter.scala 98:20:@108048.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_27 = AXICmdSplit_io_out_wdata_bits_wdata_27; // @[DRAMArbiter.scala 98:20:@108049.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_28 = AXICmdSplit_io_out_wdata_bits_wdata_28; // @[DRAMArbiter.scala 98:20:@108050.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_29 = AXICmdSplit_io_out_wdata_bits_wdata_29; // @[DRAMArbiter.scala 98:20:@108051.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_30 = AXICmdSplit_io_out_wdata_bits_wdata_30; // @[DRAMArbiter.scala 98:20:@108052.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_31 = AXICmdSplit_io_out_wdata_bits_wdata_31; // @[DRAMArbiter.scala 98:20:@108053.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_32 = AXICmdSplit_io_out_wdata_bits_wdata_32; // @[DRAMArbiter.scala 98:20:@108054.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_33 = AXICmdSplit_io_out_wdata_bits_wdata_33; // @[DRAMArbiter.scala 98:20:@108055.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_34 = AXICmdSplit_io_out_wdata_bits_wdata_34; // @[DRAMArbiter.scala 98:20:@108056.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_35 = AXICmdSplit_io_out_wdata_bits_wdata_35; // @[DRAMArbiter.scala 98:20:@108057.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_36 = AXICmdSplit_io_out_wdata_bits_wdata_36; // @[DRAMArbiter.scala 98:20:@108058.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_37 = AXICmdSplit_io_out_wdata_bits_wdata_37; // @[DRAMArbiter.scala 98:20:@108059.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_38 = AXICmdSplit_io_out_wdata_bits_wdata_38; // @[DRAMArbiter.scala 98:20:@108060.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_39 = AXICmdSplit_io_out_wdata_bits_wdata_39; // @[DRAMArbiter.scala 98:20:@108061.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_40 = AXICmdSplit_io_out_wdata_bits_wdata_40; // @[DRAMArbiter.scala 98:20:@108062.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_41 = AXICmdSplit_io_out_wdata_bits_wdata_41; // @[DRAMArbiter.scala 98:20:@108063.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_42 = AXICmdSplit_io_out_wdata_bits_wdata_42; // @[DRAMArbiter.scala 98:20:@108064.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_43 = AXICmdSplit_io_out_wdata_bits_wdata_43; // @[DRAMArbiter.scala 98:20:@108065.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_44 = AXICmdSplit_io_out_wdata_bits_wdata_44; // @[DRAMArbiter.scala 98:20:@108066.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_45 = AXICmdSplit_io_out_wdata_bits_wdata_45; // @[DRAMArbiter.scala 98:20:@108067.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_46 = AXICmdSplit_io_out_wdata_bits_wdata_46; // @[DRAMArbiter.scala 98:20:@108068.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_47 = AXICmdSplit_io_out_wdata_bits_wdata_47; // @[DRAMArbiter.scala 98:20:@108069.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_48 = AXICmdSplit_io_out_wdata_bits_wdata_48; // @[DRAMArbiter.scala 98:20:@108070.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_49 = AXICmdSplit_io_out_wdata_bits_wdata_49; // @[DRAMArbiter.scala 98:20:@108071.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_50 = AXICmdSplit_io_out_wdata_bits_wdata_50; // @[DRAMArbiter.scala 98:20:@108072.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_51 = AXICmdSplit_io_out_wdata_bits_wdata_51; // @[DRAMArbiter.scala 98:20:@108073.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_52 = AXICmdSplit_io_out_wdata_bits_wdata_52; // @[DRAMArbiter.scala 98:20:@108074.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_53 = AXICmdSplit_io_out_wdata_bits_wdata_53; // @[DRAMArbiter.scala 98:20:@108075.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_54 = AXICmdSplit_io_out_wdata_bits_wdata_54; // @[DRAMArbiter.scala 98:20:@108076.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_55 = AXICmdSplit_io_out_wdata_bits_wdata_55; // @[DRAMArbiter.scala 98:20:@108077.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_56 = AXICmdSplit_io_out_wdata_bits_wdata_56; // @[DRAMArbiter.scala 98:20:@108078.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_57 = AXICmdSplit_io_out_wdata_bits_wdata_57; // @[DRAMArbiter.scala 98:20:@108079.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_58 = AXICmdSplit_io_out_wdata_bits_wdata_58; // @[DRAMArbiter.scala 98:20:@108080.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_59 = AXICmdSplit_io_out_wdata_bits_wdata_59; // @[DRAMArbiter.scala 98:20:@108081.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_60 = AXICmdSplit_io_out_wdata_bits_wdata_60; // @[DRAMArbiter.scala 98:20:@108082.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_61 = AXICmdSplit_io_out_wdata_bits_wdata_61; // @[DRAMArbiter.scala 98:20:@108083.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_62 = AXICmdSplit_io_out_wdata_bits_wdata_62; // @[DRAMArbiter.scala 98:20:@108084.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_63 = AXICmdSplit_io_out_wdata_bits_wdata_63; // @[DRAMArbiter.scala 98:20:@108085.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@107958.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@107959.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@107960.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@107961.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@107962.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@107963.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@107964.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@107965.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@107966.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@107967.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@107968.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@107969.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@107970.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@107971.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@107972.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@107973.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@107974.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@107975.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@107976.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@107977.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@107978.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@107979.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@107980.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@107981.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@107982.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@107983.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@107984.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@107985.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@107986.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@107987.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@107988.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@107989.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@107990.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@107991.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@107992.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@107993.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@107994.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@107995.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@107996.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@107997.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@107998.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@107999.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@108000.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@108001.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@108002.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@108003.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@108004.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@108005.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@108006.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@108007.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@108008.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@108009.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@108010.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@108011.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@108012.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@108013.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@108014.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@108015.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@108016.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@108017.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@108018.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@108019.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@108020.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@108021.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@107956.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@107889.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@108302.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@108295.4]
  assign AXICmdIssue_io_out_rresp_valid = io_dram_rresp_valid; // @[DRAMArbiter.scala 99:13:@108163.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_0 = io_dram_rresp_bits_rdata_0; // @[DRAMArbiter.scala 99:13:@108099.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_1 = io_dram_rresp_bits_rdata_1; // @[DRAMArbiter.scala 99:13:@108100.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_2 = io_dram_rresp_bits_rdata_2; // @[DRAMArbiter.scala 99:13:@108101.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_3 = io_dram_rresp_bits_rdata_3; // @[DRAMArbiter.scala 99:13:@108102.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_4 = io_dram_rresp_bits_rdata_4; // @[DRAMArbiter.scala 99:13:@108103.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_5 = io_dram_rresp_bits_rdata_5; // @[DRAMArbiter.scala 99:13:@108104.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_6 = io_dram_rresp_bits_rdata_6; // @[DRAMArbiter.scala 99:13:@108105.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_7 = io_dram_rresp_bits_rdata_7; // @[DRAMArbiter.scala 99:13:@108106.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_8 = io_dram_rresp_bits_rdata_8; // @[DRAMArbiter.scala 99:13:@108107.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_9 = io_dram_rresp_bits_rdata_9; // @[DRAMArbiter.scala 99:13:@108108.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_10 = io_dram_rresp_bits_rdata_10; // @[DRAMArbiter.scala 99:13:@108109.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_11 = io_dram_rresp_bits_rdata_11; // @[DRAMArbiter.scala 99:13:@108110.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_12 = io_dram_rresp_bits_rdata_12; // @[DRAMArbiter.scala 99:13:@108111.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_13 = io_dram_rresp_bits_rdata_13; // @[DRAMArbiter.scala 99:13:@108112.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_14 = io_dram_rresp_bits_rdata_14; // @[DRAMArbiter.scala 99:13:@108113.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_15 = io_dram_rresp_bits_rdata_15; // @[DRAMArbiter.scala 99:13:@108114.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_16 = io_dram_rresp_bits_rdata_16; // @[DRAMArbiter.scala 99:13:@108115.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_17 = io_dram_rresp_bits_rdata_17; // @[DRAMArbiter.scala 99:13:@108116.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_18 = io_dram_rresp_bits_rdata_18; // @[DRAMArbiter.scala 99:13:@108117.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_19 = io_dram_rresp_bits_rdata_19; // @[DRAMArbiter.scala 99:13:@108118.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_20 = io_dram_rresp_bits_rdata_20; // @[DRAMArbiter.scala 99:13:@108119.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_21 = io_dram_rresp_bits_rdata_21; // @[DRAMArbiter.scala 99:13:@108120.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_22 = io_dram_rresp_bits_rdata_22; // @[DRAMArbiter.scala 99:13:@108121.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_23 = io_dram_rresp_bits_rdata_23; // @[DRAMArbiter.scala 99:13:@108122.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_24 = io_dram_rresp_bits_rdata_24; // @[DRAMArbiter.scala 99:13:@108123.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_25 = io_dram_rresp_bits_rdata_25; // @[DRAMArbiter.scala 99:13:@108124.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_26 = io_dram_rresp_bits_rdata_26; // @[DRAMArbiter.scala 99:13:@108125.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_27 = io_dram_rresp_bits_rdata_27; // @[DRAMArbiter.scala 99:13:@108126.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_28 = io_dram_rresp_bits_rdata_28; // @[DRAMArbiter.scala 99:13:@108127.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_29 = io_dram_rresp_bits_rdata_29; // @[DRAMArbiter.scala 99:13:@108128.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_30 = io_dram_rresp_bits_rdata_30; // @[DRAMArbiter.scala 99:13:@108129.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_31 = io_dram_rresp_bits_rdata_31; // @[DRAMArbiter.scala 99:13:@108130.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_32 = io_dram_rresp_bits_rdata_32; // @[DRAMArbiter.scala 99:13:@108131.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_33 = io_dram_rresp_bits_rdata_33; // @[DRAMArbiter.scala 99:13:@108132.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_34 = io_dram_rresp_bits_rdata_34; // @[DRAMArbiter.scala 99:13:@108133.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_35 = io_dram_rresp_bits_rdata_35; // @[DRAMArbiter.scala 99:13:@108134.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_36 = io_dram_rresp_bits_rdata_36; // @[DRAMArbiter.scala 99:13:@108135.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_37 = io_dram_rresp_bits_rdata_37; // @[DRAMArbiter.scala 99:13:@108136.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_38 = io_dram_rresp_bits_rdata_38; // @[DRAMArbiter.scala 99:13:@108137.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_39 = io_dram_rresp_bits_rdata_39; // @[DRAMArbiter.scala 99:13:@108138.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_40 = io_dram_rresp_bits_rdata_40; // @[DRAMArbiter.scala 99:13:@108139.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_41 = io_dram_rresp_bits_rdata_41; // @[DRAMArbiter.scala 99:13:@108140.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_42 = io_dram_rresp_bits_rdata_42; // @[DRAMArbiter.scala 99:13:@108141.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_43 = io_dram_rresp_bits_rdata_43; // @[DRAMArbiter.scala 99:13:@108142.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_44 = io_dram_rresp_bits_rdata_44; // @[DRAMArbiter.scala 99:13:@108143.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_45 = io_dram_rresp_bits_rdata_45; // @[DRAMArbiter.scala 99:13:@108144.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_46 = io_dram_rresp_bits_rdata_46; // @[DRAMArbiter.scala 99:13:@108145.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_47 = io_dram_rresp_bits_rdata_47; // @[DRAMArbiter.scala 99:13:@108146.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_48 = io_dram_rresp_bits_rdata_48; // @[DRAMArbiter.scala 99:13:@108147.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_49 = io_dram_rresp_bits_rdata_49; // @[DRAMArbiter.scala 99:13:@108148.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_50 = io_dram_rresp_bits_rdata_50; // @[DRAMArbiter.scala 99:13:@108149.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_51 = io_dram_rresp_bits_rdata_51; // @[DRAMArbiter.scala 99:13:@108150.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_52 = io_dram_rresp_bits_rdata_52; // @[DRAMArbiter.scala 99:13:@108151.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_53 = io_dram_rresp_bits_rdata_53; // @[DRAMArbiter.scala 99:13:@108152.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_54 = io_dram_rresp_bits_rdata_54; // @[DRAMArbiter.scala 99:13:@108153.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_55 = io_dram_rresp_bits_rdata_55; // @[DRAMArbiter.scala 99:13:@108154.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_56 = io_dram_rresp_bits_rdata_56; // @[DRAMArbiter.scala 99:13:@108155.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_57 = io_dram_rresp_bits_rdata_57; // @[DRAMArbiter.scala 99:13:@108156.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_58 = io_dram_rresp_bits_rdata_58; // @[DRAMArbiter.scala 99:13:@108157.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_59 = io_dram_rresp_bits_rdata_59; // @[DRAMArbiter.scala 99:13:@108158.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_60 = io_dram_rresp_bits_rdata_60; // @[DRAMArbiter.scala 99:13:@108159.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_61 = io_dram_rresp_bits_rdata_61; // @[DRAMArbiter.scala 99:13:@108160.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_62 = io_dram_rresp_bits_rdata_62; // @[DRAMArbiter.scala 99:13:@108161.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_63 = io_dram_rresp_bits_rdata_63; // @[DRAMArbiter.scala 99:13:@108162.4]
  assign AXICmdIssue_io_out_rresp_bits_tag = io_dram_rresp_bits_tag; // @[DRAMArbiter.scala 99:13:@108098.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@108096.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@108095.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_2028 = _RAND_0[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  _T_2042 = _RAND_1[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  _T_2049 = _RAND_2[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  _T_2056 = _RAND_3[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  _T_2066 = _RAND_4[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  _T_2074 = _RAND_5[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {2{`RANDOM}};
  _T_2082 = _RAND_6[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{`RANDOM}};
  _T_2090 = _RAND_7[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{`RANDOM}};
  _T_2097 = _RAND_8[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{`RANDOM}};
  _T_2106 = _RAND_9[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  _T_2115 = _RAND_10[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  _T_2133 = _RAND_11[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  _T_2140 = _RAND_12[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  _T_2149 = _RAND_13[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {2{`RANDOM}};
  _T_2158 = _RAND_14[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {2{`RANDOM}};
  _T_2176 = _RAND_15[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {2{`RANDOM}};
  _T_2182 = _RAND_16[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_2185 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_2188 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_2191 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_2197 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_2203 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_2209 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_2215 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {2{`RANDOM}};
  _T_2218 = _RAND_24[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_2221 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_2224 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_2227 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_2233 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_2239 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_2245 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_2251 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {2{`RANDOM}};
  _T_2323 = _RAND_32[63:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_2028 <= 64'h0;
    end else begin
      if (io_enable) begin
        _T_2028 <= _T_2031;
      end
    end
    if (reset) begin
      _T_2042 <= 64'h0;
    end else begin
      if (_T_2039) begin
        _T_2042 <= _T_2045;
      end
    end
    if (reset) begin
      _T_2049 <= 64'h0;
    end else begin
      if (_T_2046) begin
        _T_2049 <= _T_2052;
      end
    end
    if (reset) begin
      _T_2056 <= 64'h0;
    end else begin
      if (_T_2053) begin
        _T_2056 <= _T_2059;
      end
    end
    if (reset) begin
      _T_2066 <= 64'h0;
    end else begin
      if (_T_2063) begin
        _T_2066 <= _T_2069;
      end
    end
    if (reset) begin
      _T_2074 <= 64'h0;
    end else begin
      if (_T_2071) begin
        _T_2074 <= _T_2077;
      end
    end
    if (reset) begin
      _T_2082 <= 64'h0;
    end else begin
      if (_T_2079) begin
        _T_2082 <= _T_2085;
      end
    end
    if (reset) begin
      _T_2090 <= 64'h0;
    end else begin
      if (_T_2087) begin
        _T_2090 <= _T_2093;
      end
    end
    if (reset) begin
      _T_2097 <= 64'h0;
    end else begin
      if (_T_2032) begin
        _T_2097 <= _T_2100;
      end
    end
    if (reset) begin
      _T_2106 <= 64'h0;
    end else begin
      if (_T_2103) begin
        _T_2106 <= _T_2109;
      end
    end
    if (reset) begin
      _T_2115 <= 64'h0;
    end else begin
      if (_T_2112) begin
        _T_2115 <= _T_2118;
      end
    end
    if (reset) begin
      _T_2133 <= 64'h0;
    end else begin
      if (_T_2130) begin
        _T_2133 <= _T_2136;
      end
    end
    if (reset) begin
      _T_2140 <= 64'h0;
    end else begin
      if (_T_2137) begin
        _T_2140 <= _T_2143;
      end
    end
    if (reset) begin
      _T_2149 <= 64'h0;
    end else begin
      if (_T_2146) begin
        _T_2149 <= _T_2152;
      end
    end
    if (reset) begin
      _T_2158 <= 64'h0;
    end else begin
      if (_T_2155) begin
        _T_2158 <= _T_2161;
      end
    end
    if (reset) begin
      _T_2176 <= 64'h0;
    end else begin
      if (_T_2173) begin
        _T_2176 <= _T_2179;
      end
    end
    if (reset) begin
      _T_2182 <= io_dram_cmd_bits_addr;
    end else begin
      if (_T_2180) begin
        _T_2182 <= io_dram_cmd_bits_addr;
      end
    end
    if (reset) begin
      _T_2185 <= io_dram_cmd_bits_size;
    end else begin
      if (_T_2180) begin
        _T_2185 <= io_dram_cmd_bits_size;
      end
    end
    if (reset) begin
      _T_2188 <= io_dram_wdata_bits_wdata_0;
    end else begin
      if (_T_2039) begin
        _T_2188 <= io_dram_wdata_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_2191 <= io_dram_wdata_bits_wstrb_0;
    end else begin
      if (_T_2039) begin
        _T_2191 <= io_dram_wdata_bits_wstrb_0;
      end
    end
    if (reset) begin
      _T_2197 <= io_dram_wdata_bits_wdata_0;
    end else begin
      if (_T_2195) begin
        _T_2197 <= io_dram_wdata_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_2203 <= io_dram_wdata_bits_wstrb_0;
    end else begin
      if (_T_2195) begin
        _T_2203 <= io_dram_wdata_bits_wstrb_0;
      end
    end
    if (reset) begin
      _T_2209 <= io_dram_wdata_bits_wdata_0;
    end else begin
      if (_T_2207) begin
        _T_2209 <= io_dram_wdata_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_2215 <= io_dram_wdata_bits_wstrb_0;
    end else begin
      if (_T_2207) begin
        _T_2215 <= io_dram_wdata_bits_wstrb_0;
      end
    end
    if (reset) begin
      _T_2218 <= io_app_stores_0_cmd_bits_addr;
    end else begin
      if (_T_2216) begin
        _T_2218 <= io_app_stores_0_cmd_bits_addr;
      end
    end
    if (reset) begin
      _T_2221 <= io_app_stores_0_cmd_bits_size;
    end else begin
      if (_T_2216) begin
        _T_2221 <= io_app_stores_0_cmd_bits_size;
      end
    end
    if (reset) begin
      _T_2224 <= io_app_stores_0_data_bits_wdata_0;
    end else begin
      if (_T_2046) begin
        _T_2224 <= io_app_stores_0_data_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_2227 <= io_app_stores_0_data_bits_wstrb;
    end else begin
      if (_T_2046) begin
        _T_2227 <= io_app_stores_0_data_bits_wstrb;
      end
    end
    if (reset) begin
      _T_2233 <= io_app_stores_0_data_bits_wdata_0;
    end else begin
      if (_T_2231) begin
        _T_2233 <= io_app_stores_0_data_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_2239 <= io_app_stores_0_data_bits_wstrb;
    end else begin
      if (_T_2231) begin
        _T_2239 <= io_app_stores_0_data_bits_wstrb;
      end
    end
    if (reset) begin
      _T_2245 <= io_app_stores_0_data_bits_wdata_0;
    end else begin
      if (_T_2243) begin
        _T_2245 <= io_app_stores_0_data_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_2251 <= io_app_stores_0_data_bits_wstrb;
    end else begin
      if (_T_2243) begin
        _T_2251 <= io_app_stores_0_data_bits_wstrb;
      end
    end
    if (reset) begin
      _T_2323 <= 64'h0;
    end else begin
      _T_2323 <= _T_2326;
    end
  end
endmodule
module DRAMHeap( // @[:@108769.2]
  input         io_accel_0_req_valid, // @[:@108772.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@108772.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@108772.4]
  output        io_accel_0_resp_valid, // @[:@108772.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@108772.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@108772.4]
  output        io_host_0_req_valid, // @[:@108772.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@108772.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@108772.4]
  input         io_host_0_resp_valid, // @[:@108772.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@108772.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@108772.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@108779.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@108781.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@108780.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@108776.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@108775.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@108774.4]
endmodule
module FringeFF( // @[:@108815.2]
  input         clock, // @[:@108816.4]
  input         reset, // @[:@108817.4]
  input  [63:0] io_in, // @[:@108818.4]
  input         io_reset, // @[:@108818.4]
  output [63:0] io_out, // @[:@108818.4]
  input         io_enable // @[:@108818.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@108821.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@108821.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@108821.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@108821.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@108821.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@108826.4 package.scala 96:25:@108827.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@108832.6]
  RetimeWrapper_38 RetimeWrapper ( // @[package.scala 93:22:@108821.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@108826.4 package.scala 96:25:@108827.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@108832.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@108838.4]
  assign RetimeWrapper_clock = clock; // @[:@108822.4]
  assign RetimeWrapper_reset = reset; // @[:@108823.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@108825.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@108824.4]
endmodule
module MuxN_2( // @[:@140817.2]
  input  [63:0] io_ins_0, // @[:@140820.4]
  input  [63:0] io_ins_1, // @[:@140820.4]
  input  [63:0] io_ins_2, // @[:@140820.4]
  input  [63:0] io_ins_3, // @[:@140820.4]
  input  [63:0] io_ins_4, // @[:@140820.4]
  input  [63:0] io_ins_5, // @[:@140820.4]
  input  [63:0] io_ins_6, // @[:@140820.4]
  input  [63:0] io_ins_7, // @[:@140820.4]
  input  [63:0] io_ins_8, // @[:@140820.4]
  input  [63:0] io_ins_9, // @[:@140820.4]
  input  [63:0] io_ins_10, // @[:@140820.4]
  input  [63:0] io_ins_11, // @[:@140820.4]
  input  [63:0] io_ins_12, // @[:@140820.4]
  input  [63:0] io_ins_13, // @[:@140820.4]
  input  [63:0] io_ins_14, // @[:@140820.4]
  input  [63:0] io_ins_15, // @[:@140820.4]
  input  [63:0] io_ins_16, // @[:@140820.4]
  input  [63:0] io_ins_17, // @[:@140820.4]
  input  [63:0] io_ins_18, // @[:@140820.4]
  input  [63:0] io_ins_19, // @[:@140820.4]
  input  [63:0] io_ins_20, // @[:@140820.4]
  input  [63:0] io_ins_21, // @[:@140820.4]
  input  [63:0] io_ins_22, // @[:@140820.4]
  input  [63:0] io_ins_23, // @[:@140820.4]
  input  [63:0] io_ins_24, // @[:@140820.4]
  input  [63:0] io_ins_25, // @[:@140820.4]
  input  [63:0] io_ins_26, // @[:@140820.4]
  input  [63:0] io_ins_27, // @[:@140820.4]
  input  [63:0] io_ins_28, // @[:@140820.4]
  input  [63:0] io_ins_29, // @[:@140820.4]
  input  [63:0] io_ins_30, // @[:@140820.4]
  input  [63:0] io_ins_31, // @[:@140820.4]
  input  [63:0] io_ins_32, // @[:@140820.4]
  input  [63:0] io_ins_33, // @[:@140820.4]
  input  [63:0] io_ins_34, // @[:@140820.4]
  input  [63:0] io_ins_35, // @[:@140820.4]
  input  [63:0] io_ins_36, // @[:@140820.4]
  input  [63:0] io_ins_37, // @[:@140820.4]
  input  [63:0] io_ins_38, // @[:@140820.4]
  input  [63:0] io_ins_39, // @[:@140820.4]
  input  [63:0] io_ins_40, // @[:@140820.4]
  input  [63:0] io_ins_41, // @[:@140820.4]
  input  [63:0] io_ins_42, // @[:@140820.4]
  input  [63:0] io_ins_43, // @[:@140820.4]
  input  [63:0] io_ins_44, // @[:@140820.4]
  input  [63:0] io_ins_45, // @[:@140820.4]
  input  [63:0] io_ins_46, // @[:@140820.4]
  input  [63:0] io_ins_47, // @[:@140820.4]
  input  [63:0] io_ins_48, // @[:@140820.4]
  input  [63:0] io_ins_49, // @[:@140820.4]
  input  [63:0] io_ins_50, // @[:@140820.4]
  input  [63:0] io_ins_51, // @[:@140820.4]
  input  [63:0] io_ins_52, // @[:@140820.4]
  input  [63:0] io_ins_53, // @[:@140820.4]
  input  [63:0] io_ins_54, // @[:@140820.4]
  input  [63:0] io_ins_55, // @[:@140820.4]
  input  [63:0] io_ins_56, // @[:@140820.4]
  input  [63:0] io_ins_57, // @[:@140820.4]
  input  [63:0] io_ins_58, // @[:@140820.4]
  input  [63:0] io_ins_59, // @[:@140820.4]
  input  [63:0] io_ins_60, // @[:@140820.4]
  input  [63:0] io_ins_61, // @[:@140820.4]
  input  [63:0] io_ins_62, // @[:@140820.4]
  input  [63:0] io_ins_63, // @[:@140820.4]
  input  [63:0] io_ins_64, // @[:@140820.4]
  input  [63:0] io_ins_65, // @[:@140820.4]
  input  [63:0] io_ins_66, // @[:@140820.4]
  input  [63:0] io_ins_67, // @[:@140820.4]
  input  [63:0] io_ins_68, // @[:@140820.4]
  input  [63:0] io_ins_69, // @[:@140820.4]
  input  [63:0] io_ins_70, // @[:@140820.4]
  input  [63:0] io_ins_71, // @[:@140820.4]
  input  [63:0] io_ins_72, // @[:@140820.4]
  input  [63:0] io_ins_73, // @[:@140820.4]
  input  [63:0] io_ins_74, // @[:@140820.4]
  input  [63:0] io_ins_75, // @[:@140820.4]
  input  [63:0] io_ins_76, // @[:@140820.4]
  input  [63:0] io_ins_77, // @[:@140820.4]
  input  [63:0] io_ins_78, // @[:@140820.4]
  input  [63:0] io_ins_79, // @[:@140820.4]
  input  [63:0] io_ins_80, // @[:@140820.4]
  input  [63:0] io_ins_81, // @[:@140820.4]
  input  [63:0] io_ins_82, // @[:@140820.4]
  input  [63:0] io_ins_83, // @[:@140820.4]
  input  [63:0] io_ins_84, // @[:@140820.4]
  input  [63:0] io_ins_85, // @[:@140820.4]
  input  [63:0] io_ins_86, // @[:@140820.4]
  input  [63:0] io_ins_87, // @[:@140820.4]
  input  [63:0] io_ins_88, // @[:@140820.4]
  input  [63:0] io_ins_89, // @[:@140820.4]
  input  [63:0] io_ins_90, // @[:@140820.4]
  input  [63:0] io_ins_91, // @[:@140820.4]
  input  [63:0] io_ins_92, // @[:@140820.4]
  input  [63:0] io_ins_93, // @[:@140820.4]
  input  [63:0] io_ins_94, // @[:@140820.4]
  input  [63:0] io_ins_95, // @[:@140820.4]
  input  [63:0] io_ins_96, // @[:@140820.4]
  input  [63:0] io_ins_97, // @[:@140820.4]
  input  [63:0] io_ins_98, // @[:@140820.4]
  input  [63:0] io_ins_99, // @[:@140820.4]
  input  [63:0] io_ins_100, // @[:@140820.4]
  input  [63:0] io_ins_101, // @[:@140820.4]
  input  [63:0] io_ins_102, // @[:@140820.4]
  input  [63:0] io_ins_103, // @[:@140820.4]
  input  [63:0] io_ins_104, // @[:@140820.4]
  input  [63:0] io_ins_105, // @[:@140820.4]
  input  [63:0] io_ins_106, // @[:@140820.4]
  input  [63:0] io_ins_107, // @[:@140820.4]
  input  [63:0] io_ins_108, // @[:@140820.4]
  input  [63:0] io_ins_109, // @[:@140820.4]
  input  [63:0] io_ins_110, // @[:@140820.4]
  input  [63:0] io_ins_111, // @[:@140820.4]
  input  [63:0] io_ins_112, // @[:@140820.4]
  input  [63:0] io_ins_113, // @[:@140820.4]
  input  [63:0] io_ins_114, // @[:@140820.4]
  input  [63:0] io_ins_115, // @[:@140820.4]
  input  [63:0] io_ins_116, // @[:@140820.4]
  input  [63:0] io_ins_117, // @[:@140820.4]
  input  [63:0] io_ins_118, // @[:@140820.4]
  input  [63:0] io_ins_119, // @[:@140820.4]
  input  [63:0] io_ins_120, // @[:@140820.4]
  input  [63:0] io_ins_121, // @[:@140820.4]
  input  [63:0] io_ins_122, // @[:@140820.4]
  input  [63:0] io_ins_123, // @[:@140820.4]
  input  [63:0] io_ins_124, // @[:@140820.4]
  input  [63:0] io_ins_125, // @[:@140820.4]
  input  [63:0] io_ins_126, // @[:@140820.4]
  input  [63:0] io_ins_127, // @[:@140820.4]
  input  [63:0] io_ins_128, // @[:@140820.4]
  input  [63:0] io_ins_129, // @[:@140820.4]
  input  [63:0] io_ins_130, // @[:@140820.4]
  input  [63:0] io_ins_131, // @[:@140820.4]
  input  [63:0] io_ins_132, // @[:@140820.4]
  input  [63:0] io_ins_133, // @[:@140820.4]
  input  [63:0] io_ins_134, // @[:@140820.4]
  input  [63:0] io_ins_135, // @[:@140820.4]
  input  [63:0] io_ins_136, // @[:@140820.4]
  input  [63:0] io_ins_137, // @[:@140820.4]
  input  [63:0] io_ins_138, // @[:@140820.4]
  input  [63:0] io_ins_139, // @[:@140820.4]
  input  [63:0] io_ins_140, // @[:@140820.4]
  input  [63:0] io_ins_141, // @[:@140820.4]
  input  [63:0] io_ins_142, // @[:@140820.4]
  input  [63:0] io_ins_143, // @[:@140820.4]
  input  [63:0] io_ins_144, // @[:@140820.4]
  input  [63:0] io_ins_145, // @[:@140820.4]
  input  [63:0] io_ins_146, // @[:@140820.4]
  input  [63:0] io_ins_147, // @[:@140820.4]
  input  [63:0] io_ins_148, // @[:@140820.4]
  input  [63:0] io_ins_149, // @[:@140820.4]
  input  [63:0] io_ins_150, // @[:@140820.4]
  input  [63:0] io_ins_151, // @[:@140820.4]
  input  [63:0] io_ins_152, // @[:@140820.4]
  input  [63:0] io_ins_153, // @[:@140820.4]
  input  [63:0] io_ins_154, // @[:@140820.4]
  input  [63:0] io_ins_155, // @[:@140820.4]
  input  [63:0] io_ins_156, // @[:@140820.4]
  input  [63:0] io_ins_157, // @[:@140820.4]
  input  [63:0] io_ins_158, // @[:@140820.4]
  input  [63:0] io_ins_159, // @[:@140820.4]
  input  [63:0] io_ins_160, // @[:@140820.4]
  input  [63:0] io_ins_161, // @[:@140820.4]
  input  [63:0] io_ins_162, // @[:@140820.4]
  input  [63:0] io_ins_163, // @[:@140820.4]
  input  [63:0] io_ins_164, // @[:@140820.4]
  input  [63:0] io_ins_165, // @[:@140820.4]
  input  [63:0] io_ins_166, // @[:@140820.4]
  input  [63:0] io_ins_167, // @[:@140820.4]
  input  [63:0] io_ins_168, // @[:@140820.4]
  input  [63:0] io_ins_169, // @[:@140820.4]
  input  [63:0] io_ins_170, // @[:@140820.4]
  input  [63:0] io_ins_171, // @[:@140820.4]
  input  [63:0] io_ins_172, // @[:@140820.4]
  input  [63:0] io_ins_173, // @[:@140820.4]
  input  [63:0] io_ins_174, // @[:@140820.4]
  input  [63:0] io_ins_175, // @[:@140820.4]
  input  [63:0] io_ins_176, // @[:@140820.4]
  input  [63:0] io_ins_177, // @[:@140820.4]
  input  [63:0] io_ins_178, // @[:@140820.4]
  input  [63:0] io_ins_179, // @[:@140820.4]
  input  [63:0] io_ins_180, // @[:@140820.4]
  input  [63:0] io_ins_181, // @[:@140820.4]
  input  [63:0] io_ins_182, // @[:@140820.4]
  input  [63:0] io_ins_183, // @[:@140820.4]
  input  [63:0] io_ins_184, // @[:@140820.4]
  input  [63:0] io_ins_185, // @[:@140820.4]
  input  [63:0] io_ins_186, // @[:@140820.4]
  input  [63:0] io_ins_187, // @[:@140820.4]
  input  [63:0] io_ins_188, // @[:@140820.4]
  input  [63:0] io_ins_189, // @[:@140820.4]
  input  [63:0] io_ins_190, // @[:@140820.4]
  input  [63:0] io_ins_191, // @[:@140820.4]
  input  [63:0] io_ins_192, // @[:@140820.4]
  input  [63:0] io_ins_193, // @[:@140820.4]
  input  [63:0] io_ins_194, // @[:@140820.4]
  input  [63:0] io_ins_195, // @[:@140820.4]
  input  [63:0] io_ins_196, // @[:@140820.4]
  input  [63:0] io_ins_197, // @[:@140820.4]
  input  [63:0] io_ins_198, // @[:@140820.4]
  input  [63:0] io_ins_199, // @[:@140820.4]
  input  [63:0] io_ins_200, // @[:@140820.4]
  input  [63:0] io_ins_201, // @[:@140820.4]
  input  [63:0] io_ins_202, // @[:@140820.4]
  input  [63:0] io_ins_203, // @[:@140820.4]
  input  [63:0] io_ins_204, // @[:@140820.4]
  input  [63:0] io_ins_205, // @[:@140820.4]
  input  [63:0] io_ins_206, // @[:@140820.4]
  input  [63:0] io_ins_207, // @[:@140820.4]
  input  [63:0] io_ins_208, // @[:@140820.4]
  input  [63:0] io_ins_209, // @[:@140820.4]
  input  [63:0] io_ins_210, // @[:@140820.4]
  input  [63:0] io_ins_211, // @[:@140820.4]
  input  [63:0] io_ins_212, // @[:@140820.4]
  input  [63:0] io_ins_213, // @[:@140820.4]
  input  [63:0] io_ins_214, // @[:@140820.4]
  input  [63:0] io_ins_215, // @[:@140820.4]
  input  [63:0] io_ins_216, // @[:@140820.4]
  input  [63:0] io_ins_217, // @[:@140820.4]
  input  [63:0] io_ins_218, // @[:@140820.4]
  input  [63:0] io_ins_219, // @[:@140820.4]
  input  [63:0] io_ins_220, // @[:@140820.4]
  input  [63:0] io_ins_221, // @[:@140820.4]
  input  [63:0] io_ins_222, // @[:@140820.4]
  input  [63:0] io_ins_223, // @[:@140820.4]
  input  [63:0] io_ins_224, // @[:@140820.4]
  input  [63:0] io_ins_225, // @[:@140820.4]
  input  [63:0] io_ins_226, // @[:@140820.4]
  input  [63:0] io_ins_227, // @[:@140820.4]
  input  [63:0] io_ins_228, // @[:@140820.4]
  input  [63:0] io_ins_229, // @[:@140820.4]
  input  [63:0] io_ins_230, // @[:@140820.4]
  input  [63:0] io_ins_231, // @[:@140820.4]
  input  [63:0] io_ins_232, // @[:@140820.4]
  input  [63:0] io_ins_233, // @[:@140820.4]
  input  [63:0] io_ins_234, // @[:@140820.4]
  input  [63:0] io_ins_235, // @[:@140820.4]
  input  [63:0] io_ins_236, // @[:@140820.4]
  input  [63:0] io_ins_237, // @[:@140820.4]
  input  [63:0] io_ins_238, // @[:@140820.4]
  input  [63:0] io_ins_239, // @[:@140820.4]
  input  [63:0] io_ins_240, // @[:@140820.4]
  input  [63:0] io_ins_241, // @[:@140820.4]
  input  [63:0] io_ins_242, // @[:@140820.4]
  input  [63:0] io_ins_243, // @[:@140820.4]
  input  [63:0] io_ins_244, // @[:@140820.4]
  input  [63:0] io_ins_245, // @[:@140820.4]
  input  [63:0] io_ins_246, // @[:@140820.4]
  input  [63:0] io_ins_247, // @[:@140820.4]
  input  [63:0] io_ins_248, // @[:@140820.4]
  input  [63:0] io_ins_249, // @[:@140820.4]
  input  [63:0] io_ins_250, // @[:@140820.4]
  input  [63:0] io_ins_251, // @[:@140820.4]
  input  [63:0] io_ins_252, // @[:@140820.4]
  input  [63:0] io_ins_253, // @[:@140820.4]
  input  [63:0] io_ins_254, // @[:@140820.4]
  input  [63:0] io_ins_255, // @[:@140820.4]
  input  [63:0] io_ins_256, // @[:@140820.4]
  input  [63:0] io_ins_257, // @[:@140820.4]
  input  [63:0] io_ins_258, // @[:@140820.4]
  input  [63:0] io_ins_259, // @[:@140820.4]
  input  [63:0] io_ins_260, // @[:@140820.4]
  input  [63:0] io_ins_261, // @[:@140820.4]
  input  [63:0] io_ins_262, // @[:@140820.4]
  input  [63:0] io_ins_263, // @[:@140820.4]
  input  [63:0] io_ins_264, // @[:@140820.4]
  input  [63:0] io_ins_265, // @[:@140820.4]
  input  [63:0] io_ins_266, // @[:@140820.4]
  input  [63:0] io_ins_267, // @[:@140820.4]
  input  [63:0] io_ins_268, // @[:@140820.4]
  input  [63:0] io_ins_269, // @[:@140820.4]
  input  [63:0] io_ins_270, // @[:@140820.4]
  input  [63:0] io_ins_271, // @[:@140820.4]
  input  [63:0] io_ins_272, // @[:@140820.4]
  input  [63:0] io_ins_273, // @[:@140820.4]
  input  [63:0] io_ins_274, // @[:@140820.4]
  input  [63:0] io_ins_275, // @[:@140820.4]
  input  [63:0] io_ins_276, // @[:@140820.4]
  input  [63:0] io_ins_277, // @[:@140820.4]
  input  [63:0] io_ins_278, // @[:@140820.4]
  input  [63:0] io_ins_279, // @[:@140820.4]
  input  [63:0] io_ins_280, // @[:@140820.4]
  input  [63:0] io_ins_281, // @[:@140820.4]
  input  [63:0] io_ins_282, // @[:@140820.4]
  input  [63:0] io_ins_283, // @[:@140820.4]
  input  [63:0] io_ins_284, // @[:@140820.4]
  input  [63:0] io_ins_285, // @[:@140820.4]
  input  [63:0] io_ins_286, // @[:@140820.4]
  input  [63:0] io_ins_287, // @[:@140820.4]
  input  [63:0] io_ins_288, // @[:@140820.4]
  input  [63:0] io_ins_289, // @[:@140820.4]
  input  [63:0] io_ins_290, // @[:@140820.4]
  input  [63:0] io_ins_291, // @[:@140820.4]
  input  [63:0] io_ins_292, // @[:@140820.4]
  input  [63:0] io_ins_293, // @[:@140820.4]
  input  [63:0] io_ins_294, // @[:@140820.4]
  input  [63:0] io_ins_295, // @[:@140820.4]
  input  [63:0] io_ins_296, // @[:@140820.4]
  input  [63:0] io_ins_297, // @[:@140820.4]
  input  [63:0] io_ins_298, // @[:@140820.4]
  input  [63:0] io_ins_299, // @[:@140820.4]
  input  [63:0] io_ins_300, // @[:@140820.4]
  input  [63:0] io_ins_301, // @[:@140820.4]
  input  [63:0] io_ins_302, // @[:@140820.4]
  input  [63:0] io_ins_303, // @[:@140820.4]
  input  [63:0] io_ins_304, // @[:@140820.4]
  input  [63:0] io_ins_305, // @[:@140820.4]
  input  [63:0] io_ins_306, // @[:@140820.4]
  input  [63:0] io_ins_307, // @[:@140820.4]
  input  [63:0] io_ins_308, // @[:@140820.4]
  input  [63:0] io_ins_309, // @[:@140820.4]
  input  [63:0] io_ins_310, // @[:@140820.4]
  input  [63:0] io_ins_311, // @[:@140820.4]
  input  [63:0] io_ins_312, // @[:@140820.4]
  input  [63:0] io_ins_313, // @[:@140820.4]
  input  [63:0] io_ins_314, // @[:@140820.4]
  input  [63:0] io_ins_315, // @[:@140820.4]
  input  [63:0] io_ins_316, // @[:@140820.4]
  input  [63:0] io_ins_317, // @[:@140820.4]
  input  [63:0] io_ins_318, // @[:@140820.4]
  input  [63:0] io_ins_319, // @[:@140820.4]
  input  [63:0] io_ins_320, // @[:@140820.4]
  input  [63:0] io_ins_321, // @[:@140820.4]
  input  [63:0] io_ins_322, // @[:@140820.4]
  input  [63:0] io_ins_323, // @[:@140820.4]
  input  [63:0] io_ins_324, // @[:@140820.4]
  input  [63:0] io_ins_325, // @[:@140820.4]
  input  [63:0] io_ins_326, // @[:@140820.4]
  input  [63:0] io_ins_327, // @[:@140820.4]
  input  [63:0] io_ins_328, // @[:@140820.4]
  input  [63:0] io_ins_329, // @[:@140820.4]
  input  [63:0] io_ins_330, // @[:@140820.4]
  input  [63:0] io_ins_331, // @[:@140820.4]
  input  [63:0] io_ins_332, // @[:@140820.4]
  input  [63:0] io_ins_333, // @[:@140820.4]
  input  [63:0] io_ins_334, // @[:@140820.4]
  input  [63:0] io_ins_335, // @[:@140820.4]
  input  [63:0] io_ins_336, // @[:@140820.4]
  input  [63:0] io_ins_337, // @[:@140820.4]
  input  [63:0] io_ins_338, // @[:@140820.4]
  input  [63:0] io_ins_339, // @[:@140820.4]
  input  [63:0] io_ins_340, // @[:@140820.4]
  input  [63:0] io_ins_341, // @[:@140820.4]
  input  [63:0] io_ins_342, // @[:@140820.4]
  input  [63:0] io_ins_343, // @[:@140820.4]
  input  [63:0] io_ins_344, // @[:@140820.4]
  input  [63:0] io_ins_345, // @[:@140820.4]
  input  [63:0] io_ins_346, // @[:@140820.4]
  input  [63:0] io_ins_347, // @[:@140820.4]
  input  [63:0] io_ins_348, // @[:@140820.4]
  input  [63:0] io_ins_349, // @[:@140820.4]
  input  [63:0] io_ins_350, // @[:@140820.4]
  input  [63:0] io_ins_351, // @[:@140820.4]
  input  [63:0] io_ins_352, // @[:@140820.4]
  input  [63:0] io_ins_353, // @[:@140820.4]
  input  [63:0] io_ins_354, // @[:@140820.4]
  input  [63:0] io_ins_355, // @[:@140820.4]
  input  [63:0] io_ins_356, // @[:@140820.4]
  input  [63:0] io_ins_357, // @[:@140820.4]
  input  [63:0] io_ins_358, // @[:@140820.4]
  input  [63:0] io_ins_359, // @[:@140820.4]
  input  [63:0] io_ins_360, // @[:@140820.4]
  input  [63:0] io_ins_361, // @[:@140820.4]
  input  [63:0] io_ins_362, // @[:@140820.4]
  input  [63:0] io_ins_363, // @[:@140820.4]
  input  [63:0] io_ins_364, // @[:@140820.4]
  input  [63:0] io_ins_365, // @[:@140820.4]
  input  [63:0] io_ins_366, // @[:@140820.4]
  input  [63:0] io_ins_367, // @[:@140820.4]
  input  [63:0] io_ins_368, // @[:@140820.4]
  input  [63:0] io_ins_369, // @[:@140820.4]
  input  [63:0] io_ins_370, // @[:@140820.4]
  input  [63:0] io_ins_371, // @[:@140820.4]
  input  [63:0] io_ins_372, // @[:@140820.4]
  input  [63:0] io_ins_373, // @[:@140820.4]
  input  [63:0] io_ins_374, // @[:@140820.4]
  input  [63:0] io_ins_375, // @[:@140820.4]
  input  [63:0] io_ins_376, // @[:@140820.4]
  input  [63:0] io_ins_377, // @[:@140820.4]
  input  [63:0] io_ins_378, // @[:@140820.4]
  input  [63:0] io_ins_379, // @[:@140820.4]
  input  [63:0] io_ins_380, // @[:@140820.4]
  input  [63:0] io_ins_381, // @[:@140820.4]
  input  [63:0] io_ins_382, // @[:@140820.4]
  input  [63:0] io_ins_383, // @[:@140820.4]
  input  [63:0] io_ins_384, // @[:@140820.4]
  input  [63:0] io_ins_385, // @[:@140820.4]
  input  [63:0] io_ins_386, // @[:@140820.4]
  input  [63:0] io_ins_387, // @[:@140820.4]
  input  [63:0] io_ins_388, // @[:@140820.4]
  input  [63:0] io_ins_389, // @[:@140820.4]
  input  [63:0] io_ins_390, // @[:@140820.4]
  input  [63:0] io_ins_391, // @[:@140820.4]
  input  [63:0] io_ins_392, // @[:@140820.4]
  input  [63:0] io_ins_393, // @[:@140820.4]
  input  [63:0] io_ins_394, // @[:@140820.4]
  input  [63:0] io_ins_395, // @[:@140820.4]
  input  [63:0] io_ins_396, // @[:@140820.4]
  input  [63:0] io_ins_397, // @[:@140820.4]
  input  [63:0] io_ins_398, // @[:@140820.4]
  input  [63:0] io_ins_399, // @[:@140820.4]
  input  [63:0] io_ins_400, // @[:@140820.4]
  input  [63:0] io_ins_401, // @[:@140820.4]
  input  [63:0] io_ins_402, // @[:@140820.4]
  input  [63:0] io_ins_403, // @[:@140820.4]
  input  [63:0] io_ins_404, // @[:@140820.4]
  input  [63:0] io_ins_405, // @[:@140820.4]
  input  [63:0] io_ins_406, // @[:@140820.4]
  input  [63:0] io_ins_407, // @[:@140820.4]
  input  [63:0] io_ins_408, // @[:@140820.4]
  input  [63:0] io_ins_409, // @[:@140820.4]
  input  [63:0] io_ins_410, // @[:@140820.4]
  input  [63:0] io_ins_411, // @[:@140820.4]
  input  [63:0] io_ins_412, // @[:@140820.4]
  input  [63:0] io_ins_413, // @[:@140820.4]
  input  [63:0] io_ins_414, // @[:@140820.4]
  input  [63:0] io_ins_415, // @[:@140820.4]
  input  [63:0] io_ins_416, // @[:@140820.4]
  input  [63:0] io_ins_417, // @[:@140820.4]
  input  [63:0] io_ins_418, // @[:@140820.4]
  input  [63:0] io_ins_419, // @[:@140820.4]
  input  [63:0] io_ins_420, // @[:@140820.4]
  input  [63:0] io_ins_421, // @[:@140820.4]
  input  [63:0] io_ins_422, // @[:@140820.4]
  input  [63:0] io_ins_423, // @[:@140820.4]
  input  [63:0] io_ins_424, // @[:@140820.4]
  input  [63:0] io_ins_425, // @[:@140820.4]
  input  [63:0] io_ins_426, // @[:@140820.4]
  input  [63:0] io_ins_427, // @[:@140820.4]
  input  [63:0] io_ins_428, // @[:@140820.4]
  input  [63:0] io_ins_429, // @[:@140820.4]
  input  [63:0] io_ins_430, // @[:@140820.4]
  input  [63:0] io_ins_431, // @[:@140820.4]
  input  [63:0] io_ins_432, // @[:@140820.4]
  input  [63:0] io_ins_433, // @[:@140820.4]
  input  [63:0] io_ins_434, // @[:@140820.4]
  input  [63:0] io_ins_435, // @[:@140820.4]
  input  [63:0] io_ins_436, // @[:@140820.4]
  input  [63:0] io_ins_437, // @[:@140820.4]
  input  [63:0] io_ins_438, // @[:@140820.4]
  input  [63:0] io_ins_439, // @[:@140820.4]
  input  [63:0] io_ins_440, // @[:@140820.4]
  input  [63:0] io_ins_441, // @[:@140820.4]
  input  [63:0] io_ins_442, // @[:@140820.4]
  input  [63:0] io_ins_443, // @[:@140820.4]
  input  [63:0] io_ins_444, // @[:@140820.4]
  input  [63:0] io_ins_445, // @[:@140820.4]
  input  [63:0] io_ins_446, // @[:@140820.4]
  input  [63:0] io_ins_447, // @[:@140820.4]
  input  [63:0] io_ins_448, // @[:@140820.4]
  input  [63:0] io_ins_449, // @[:@140820.4]
  input  [63:0] io_ins_450, // @[:@140820.4]
  input  [63:0] io_ins_451, // @[:@140820.4]
  input  [63:0] io_ins_452, // @[:@140820.4]
  input  [63:0] io_ins_453, // @[:@140820.4]
  input  [63:0] io_ins_454, // @[:@140820.4]
  input  [63:0] io_ins_455, // @[:@140820.4]
  input  [63:0] io_ins_456, // @[:@140820.4]
  input  [63:0] io_ins_457, // @[:@140820.4]
  input  [63:0] io_ins_458, // @[:@140820.4]
  input  [63:0] io_ins_459, // @[:@140820.4]
  input  [63:0] io_ins_460, // @[:@140820.4]
  input  [63:0] io_ins_461, // @[:@140820.4]
  input  [63:0] io_ins_462, // @[:@140820.4]
  input  [63:0] io_ins_463, // @[:@140820.4]
  input  [63:0] io_ins_464, // @[:@140820.4]
  input  [63:0] io_ins_465, // @[:@140820.4]
  input  [63:0] io_ins_466, // @[:@140820.4]
  input  [63:0] io_ins_467, // @[:@140820.4]
  input  [63:0] io_ins_468, // @[:@140820.4]
  input  [63:0] io_ins_469, // @[:@140820.4]
  input  [63:0] io_ins_470, // @[:@140820.4]
  input  [63:0] io_ins_471, // @[:@140820.4]
  input  [63:0] io_ins_472, // @[:@140820.4]
  input  [63:0] io_ins_473, // @[:@140820.4]
  input  [63:0] io_ins_474, // @[:@140820.4]
  input  [63:0] io_ins_475, // @[:@140820.4]
  input  [63:0] io_ins_476, // @[:@140820.4]
  input  [63:0] io_ins_477, // @[:@140820.4]
  input  [63:0] io_ins_478, // @[:@140820.4]
  input  [63:0] io_ins_479, // @[:@140820.4]
  input  [63:0] io_ins_480, // @[:@140820.4]
  input  [63:0] io_ins_481, // @[:@140820.4]
  input  [63:0] io_ins_482, // @[:@140820.4]
  input  [63:0] io_ins_483, // @[:@140820.4]
  input  [63:0] io_ins_484, // @[:@140820.4]
  input  [63:0] io_ins_485, // @[:@140820.4]
  input  [63:0] io_ins_486, // @[:@140820.4]
  input  [63:0] io_ins_487, // @[:@140820.4]
  input  [63:0] io_ins_488, // @[:@140820.4]
  input  [63:0] io_ins_489, // @[:@140820.4]
  input  [63:0] io_ins_490, // @[:@140820.4]
  input  [63:0] io_ins_491, // @[:@140820.4]
  input  [63:0] io_ins_492, // @[:@140820.4]
  input  [63:0] io_ins_493, // @[:@140820.4]
  input  [63:0] io_ins_494, // @[:@140820.4]
  input  [63:0] io_ins_495, // @[:@140820.4]
  input  [63:0] io_ins_496, // @[:@140820.4]
  input  [63:0] io_ins_497, // @[:@140820.4]
  input  [63:0] io_ins_498, // @[:@140820.4]
  input  [63:0] io_ins_499, // @[:@140820.4]
  input  [63:0] io_ins_500, // @[:@140820.4]
  input  [63:0] io_ins_501, // @[:@140820.4]
  input  [63:0] io_ins_502, // @[:@140820.4]
  input  [63:0] io_ins_503, // @[:@140820.4]
  input  [63:0] io_ins_504, // @[:@140820.4]
  input  [63:0] io_ins_505, // @[:@140820.4]
  input  [63:0] io_ins_506, // @[:@140820.4]
  input  [63:0] io_ins_507, // @[:@140820.4]
  input  [63:0] io_ins_508, // @[:@140820.4]
  input  [63:0] io_ins_509, // @[:@140820.4]
  input  [63:0] io_ins_510, // @[:@140820.4]
  input  [63:0] io_ins_511, // @[:@140820.4]
  input  [63:0] io_ins_512, // @[:@140820.4]
  input  [63:0] io_ins_513, // @[:@140820.4]
  input  [63:0] io_ins_514, // @[:@140820.4]
  input  [63:0] io_ins_515, // @[:@140820.4]
  input  [63:0] io_ins_516, // @[:@140820.4]
  input  [63:0] io_ins_517, // @[:@140820.4]
  input  [63:0] io_ins_518, // @[:@140820.4]
  input  [63:0] io_ins_519, // @[:@140820.4]
  input  [63:0] io_ins_520, // @[:@140820.4]
  input  [63:0] io_ins_521, // @[:@140820.4]
  input  [63:0] io_ins_522, // @[:@140820.4]
  input  [63:0] io_ins_523, // @[:@140820.4]
  input  [63:0] io_ins_524, // @[:@140820.4]
  input  [63:0] io_ins_525, // @[:@140820.4]
  input  [63:0] io_ins_526, // @[:@140820.4]
  input  [63:0] io_ins_527, // @[:@140820.4]
  input  [63:0] io_ins_528, // @[:@140820.4]
  input  [63:0] io_ins_529, // @[:@140820.4]
  input  [63:0] io_ins_530, // @[:@140820.4]
  input  [63:0] io_ins_531, // @[:@140820.4]
  input  [63:0] io_ins_532, // @[:@140820.4]
  input  [63:0] io_ins_533, // @[:@140820.4]
  input  [63:0] io_ins_534, // @[:@140820.4]
  input  [63:0] io_ins_535, // @[:@140820.4]
  input  [63:0] io_ins_536, // @[:@140820.4]
  input  [63:0] io_ins_537, // @[:@140820.4]
  input  [63:0] io_ins_538, // @[:@140820.4]
  input  [63:0] io_ins_539, // @[:@140820.4]
  input  [63:0] io_ins_540, // @[:@140820.4]
  input  [63:0] io_ins_541, // @[:@140820.4]
  input  [63:0] io_ins_542, // @[:@140820.4]
  input  [63:0] io_ins_543, // @[:@140820.4]
  input  [63:0] io_ins_544, // @[:@140820.4]
  input  [63:0] io_ins_545, // @[:@140820.4]
  input  [63:0] io_ins_546, // @[:@140820.4]
  input  [63:0] io_ins_547, // @[:@140820.4]
  input  [63:0] io_ins_548, // @[:@140820.4]
  input  [63:0] io_ins_549, // @[:@140820.4]
  input  [63:0] io_ins_550, // @[:@140820.4]
  input  [63:0] io_ins_551, // @[:@140820.4]
  input  [63:0] io_ins_552, // @[:@140820.4]
  input  [63:0] io_ins_553, // @[:@140820.4]
  input  [63:0] io_ins_554, // @[:@140820.4]
  input  [63:0] io_ins_555, // @[:@140820.4]
  input  [63:0] io_ins_556, // @[:@140820.4]
  input  [63:0] io_ins_557, // @[:@140820.4]
  input  [63:0] io_ins_558, // @[:@140820.4]
  input  [63:0] io_ins_559, // @[:@140820.4]
  input  [63:0] io_ins_560, // @[:@140820.4]
  input  [63:0] io_ins_561, // @[:@140820.4]
  input  [9:0]  io_sel, // @[:@140820.4]
  output [63:0] io_out // @[:@140820.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_502; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_503; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_504; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_505; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_506; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_507; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_508; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_509; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_510; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_511; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_512; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_513; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_514; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_515; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_516; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_517; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_518; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_519; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_520; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_521; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_522; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_523; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_524; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_525; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_526; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_527; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_528; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_529; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_530; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_531; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_532; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_533; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_534; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_535; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_536; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_537; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_538; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_539; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_540; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_541; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_542; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_543; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_544; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_545; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_546; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_547; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_548; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_549; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_550; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_551; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_552; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_553; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_554; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_555; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_556; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_557; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_558; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_559; // @[MuxN.scala 16:10:@140822.4]
  wire [63:0] _GEN_560; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_1 = 10'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_2 = 10'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_3 = 10'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_4 = 10'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_5 = 10'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_6 = 10'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_7 = 10'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_8 = 10'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_9 = 10'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_10 = 10'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_11 = 10'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_12 = 10'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_13 = 10'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_14 = 10'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_15 = 10'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_16 = 10'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_17 = 10'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_18 = 10'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_19 = 10'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_20 = 10'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_21 = 10'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_22 = 10'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_23 = 10'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_24 = 10'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_25 = 10'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_26 = 10'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_27 = 10'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_28 = 10'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_29 = 10'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_30 = 10'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_31 = 10'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_32 = 10'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_33 = 10'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_34 = 10'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_35 = 10'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_36 = 10'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_37 = 10'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_38 = 10'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_39 = 10'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_40 = 10'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_41 = 10'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_42 = 10'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_43 = 10'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_44 = 10'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_45 = 10'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_46 = 10'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_47 = 10'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_48 = 10'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_49 = 10'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_50 = 10'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_51 = 10'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_52 = 10'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_53 = 10'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_54 = 10'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_55 = 10'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_56 = 10'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_57 = 10'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_58 = 10'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_59 = 10'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_60 = 10'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_61 = 10'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_62 = 10'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_63 = 10'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_64 = 10'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_65 = 10'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_66 = 10'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_67 = 10'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_68 = 10'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_69 = 10'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_70 = 10'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_71 = 10'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_72 = 10'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_73 = 10'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_74 = 10'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_75 = 10'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_76 = 10'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_77 = 10'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_78 = 10'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_79 = 10'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_80 = 10'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_81 = 10'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_82 = 10'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_83 = 10'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_84 = 10'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_85 = 10'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_86 = 10'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_87 = 10'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_88 = 10'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_89 = 10'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_90 = 10'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_91 = 10'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_92 = 10'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_93 = 10'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_94 = 10'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_95 = 10'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_96 = 10'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_97 = 10'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_98 = 10'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_99 = 10'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_100 = 10'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_101 = 10'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_102 = 10'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_103 = 10'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_104 = 10'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_105 = 10'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_106 = 10'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_107 = 10'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_108 = 10'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_109 = 10'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_110 = 10'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_111 = 10'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_112 = 10'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_113 = 10'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_114 = 10'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_115 = 10'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_116 = 10'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_117 = 10'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_118 = 10'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_119 = 10'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_120 = 10'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_121 = 10'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_122 = 10'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_123 = 10'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_124 = 10'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_125 = 10'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_126 = 10'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_127 = 10'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_128 = 10'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_129 = 10'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_130 = 10'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_131 = 10'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_132 = 10'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_133 = 10'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_134 = 10'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_135 = 10'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_136 = 10'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_137 = 10'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_138 = 10'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_139 = 10'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_140 = 10'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_141 = 10'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_142 = 10'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_143 = 10'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_144 = 10'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_145 = 10'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_146 = 10'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_147 = 10'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_148 = 10'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_149 = 10'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_150 = 10'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_151 = 10'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_152 = 10'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_153 = 10'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_154 = 10'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_155 = 10'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_156 = 10'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_157 = 10'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_158 = 10'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_159 = 10'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_160 = 10'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_161 = 10'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_162 = 10'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_163 = 10'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_164 = 10'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_165 = 10'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_166 = 10'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_167 = 10'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_168 = 10'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_169 = 10'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_170 = 10'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_171 = 10'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_172 = 10'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_173 = 10'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_174 = 10'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_175 = 10'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_176 = 10'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_177 = 10'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_178 = 10'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_179 = 10'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_180 = 10'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_181 = 10'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_182 = 10'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_183 = 10'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_184 = 10'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_185 = 10'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_186 = 10'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_187 = 10'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_188 = 10'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_189 = 10'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_190 = 10'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_191 = 10'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_192 = 10'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_193 = 10'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_194 = 10'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_195 = 10'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_196 = 10'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_197 = 10'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_198 = 10'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_199 = 10'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_200 = 10'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_201 = 10'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_202 = 10'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_203 = 10'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_204 = 10'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_205 = 10'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_206 = 10'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_207 = 10'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_208 = 10'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_209 = 10'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_210 = 10'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_211 = 10'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_212 = 10'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_213 = 10'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_214 = 10'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_215 = 10'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_216 = 10'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_217 = 10'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_218 = 10'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_219 = 10'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_220 = 10'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_221 = 10'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_222 = 10'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_223 = 10'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_224 = 10'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_225 = 10'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_226 = 10'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_227 = 10'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_228 = 10'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_229 = 10'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_230 = 10'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_231 = 10'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_232 = 10'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_233 = 10'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_234 = 10'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_235 = 10'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_236 = 10'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_237 = 10'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_238 = 10'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_239 = 10'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_240 = 10'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_241 = 10'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_242 = 10'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_243 = 10'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_244 = 10'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_245 = 10'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_246 = 10'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_247 = 10'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_248 = 10'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_249 = 10'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_250 = 10'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_251 = 10'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_252 = 10'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_253 = 10'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_254 = 10'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_255 = 10'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_256 = 10'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_257 = 10'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_258 = 10'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_259 = 10'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_260 = 10'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_261 = 10'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_262 = 10'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_263 = 10'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_264 = 10'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_265 = 10'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_266 = 10'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_267 = 10'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_268 = 10'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_269 = 10'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_270 = 10'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_271 = 10'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_272 = 10'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_273 = 10'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_274 = 10'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_275 = 10'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_276 = 10'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_277 = 10'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_278 = 10'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_279 = 10'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_280 = 10'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_281 = 10'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_282 = 10'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_283 = 10'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_284 = 10'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_285 = 10'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_286 = 10'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_287 = 10'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_288 = 10'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_289 = 10'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_290 = 10'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_291 = 10'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_292 = 10'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_293 = 10'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_294 = 10'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_295 = 10'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_296 = 10'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_297 = 10'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_298 = 10'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_299 = 10'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_300 = 10'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_301 = 10'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_302 = 10'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_303 = 10'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_304 = 10'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_305 = 10'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_306 = 10'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_307 = 10'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_308 = 10'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_309 = 10'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_310 = 10'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_311 = 10'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_312 = 10'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_313 = 10'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_314 = 10'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_315 = 10'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_316 = 10'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_317 = 10'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_318 = 10'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_319 = 10'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_320 = 10'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_321 = 10'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_322 = 10'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_323 = 10'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_324 = 10'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_325 = 10'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_326 = 10'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_327 = 10'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_328 = 10'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_329 = 10'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_330 = 10'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_331 = 10'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_332 = 10'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_333 = 10'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_334 = 10'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_335 = 10'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_336 = 10'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_337 = 10'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_338 = 10'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_339 = 10'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_340 = 10'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_341 = 10'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_342 = 10'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_343 = 10'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_344 = 10'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_345 = 10'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_346 = 10'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_347 = 10'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_348 = 10'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_349 = 10'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_350 = 10'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_351 = 10'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_352 = 10'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_353 = 10'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_354 = 10'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_355 = 10'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_356 = 10'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_357 = 10'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_358 = 10'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_359 = 10'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_360 = 10'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_361 = 10'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_362 = 10'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_363 = 10'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_364 = 10'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_365 = 10'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_366 = 10'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_367 = 10'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_368 = 10'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_369 = 10'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_370 = 10'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_371 = 10'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_372 = 10'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_373 = 10'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_374 = 10'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_375 = 10'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_376 = 10'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_377 = 10'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_378 = 10'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_379 = 10'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_380 = 10'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_381 = 10'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_382 = 10'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_383 = 10'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_384 = 10'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_385 = 10'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_386 = 10'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_387 = 10'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_388 = 10'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_389 = 10'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_390 = 10'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_391 = 10'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_392 = 10'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_393 = 10'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_394 = 10'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_395 = 10'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_396 = 10'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_397 = 10'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_398 = 10'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_399 = 10'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_400 = 10'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_401 = 10'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_402 = 10'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_403 = 10'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_404 = 10'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_405 = 10'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_406 = 10'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_407 = 10'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_408 = 10'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_409 = 10'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_410 = 10'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_411 = 10'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_412 = 10'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_413 = 10'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_414 = 10'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_415 = 10'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_416 = 10'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_417 = 10'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_418 = 10'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_419 = 10'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_420 = 10'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_421 = 10'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_422 = 10'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_423 = 10'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_424 = 10'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_425 = 10'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_426 = 10'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_427 = 10'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_428 = 10'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_429 = 10'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_430 = 10'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_431 = 10'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_432 = 10'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_433 = 10'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_434 = 10'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_435 = 10'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_436 = 10'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_437 = 10'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_438 = 10'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_439 = 10'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_440 = 10'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_441 = 10'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_442 = 10'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_443 = 10'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_444 = 10'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_445 = 10'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_446 = 10'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_447 = 10'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_448 = 10'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_449 = 10'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_450 = 10'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_451 = 10'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_452 = 10'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_453 = 10'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_454 = 10'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_455 = 10'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_456 = 10'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_457 = 10'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_458 = 10'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_459 = 10'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_460 = 10'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_461 = 10'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_462 = 10'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_463 = 10'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_464 = 10'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_465 = 10'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_466 = 10'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_467 = 10'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_468 = 10'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_469 = 10'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_470 = 10'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_471 = 10'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_472 = 10'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_473 = 10'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_474 = 10'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_475 = 10'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_476 = 10'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_477 = 10'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_478 = 10'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_479 = 10'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_480 = 10'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_481 = 10'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_482 = 10'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_483 = 10'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_484 = 10'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_485 = 10'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_486 = 10'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_487 = 10'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_488 = 10'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_489 = 10'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_490 = 10'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_491 = 10'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_492 = 10'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_493 = 10'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_494 = 10'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_495 = 10'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_496 = 10'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_497 = 10'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_498 = 10'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_499 = 10'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_500 = 10'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_501 = 10'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_502 = 10'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_503 = 10'h1f7 == io_sel ? io_ins_503 : _GEN_502; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_504 = 10'h1f8 == io_sel ? io_ins_504 : _GEN_503; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_505 = 10'h1f9 == io_sel ? io_ins_505 : _GEN_504; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_506 = 10'h1fa == io_sel ? io_ins_506 : _GEN_505; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_507 = 10'h1fb == io_sel ? io_ins_507 : _GEN_506; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_508 = 10'h1fc == io_sel ? io_ins_508 : _GEN_507; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_509 = 10'h1fd == io_sel ? io_ins_509 : _GEN_508; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_510 = 10'h1fe == io_sel ? io_ins_510 : _GEN_509; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_511 = 10'h1ff == io_sel ? io_ins_511 : _GEN_510; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_512 = 10'h200 == io_sel ? io_ins_512 : _GEN_511; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_513 = 10'h201 == io_sel ? io_ins_513 : _GEN_512; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_514 = 10'h202 == io_sel ? io_ins_514 : _GEN_513; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_515 = 10'h203 == io_sel ? io_ins_515 : _GEN_514; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_516 = 10'h204 == io_sel ? io_ins_516 : _GEN_515; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_517 = 10'h205 == io_sel ? io_ins_517 : _GEN_516; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_518 = 10'h206 == io_sel ? io_ins_518 : _GEN_517; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_519 = 10'h207 == io_sel ? io_ins_519 : _GEN_518; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_520 = 10'h208 == io_sel ? io_ins_520 : _GEN_519; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_521 = 10'h209 == io_sel ? io_ins_521 : _GEN_520; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_522 = 10'h20a == io_sel ? io_ins_522 : _GEN_521; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_523 = 10'h20b == io_sel ? io_ins_523 : _GEN_522; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_524 = 10'h20c == io_sel ? io_ins_524 : _GEN_523; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_525 = 10'h20d == io_sel ? io_ins_525 : _GEN_524; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_526 = 10'h20e == io_sel ? io_ins_526 : _GEN_525; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_527 = 10'h20f == io_sel ? io_ins_527 : _GEN_526; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_528 = 10'h210 == io_sel ? io_ins_528 : _GEN_527; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_529 = 10'h211 == io_sel ? io_ins_529 : _GEN_528; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_530 = 10'h212 == io_sel ? io_ins_530 : _GEN_529; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_531 = 10'h213 == io_sel ? io_ins_531 : _GEN_530; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_532 = 10'h214 == io_sel ? io_ins_532 : _GEN_531; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_533 = 10'h215 == io_sel ? io_ins_533 : _GEN_532; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_534 = 10'h216 == io_sel ? io_ins_534 : _GEN_533; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_535 = 10'h217 == io_sel ? io_ins_535 : _GEN_534; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_536 = 10'h218 == io_sel ? io_ins_536 : _GEN_535; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_537 = 10'h219 == io_sel ? io_ins_537 : _GEN_536; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_538 = 10'h21a == io_sel ? io_ins_538 : _GEN_537; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_539 = 10'h21b == io_sel ? io_ins_539 : _GEN_538; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_540 = 10'h21c == io_sel ? io_ins_540 : _GEN_539; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_541 = 10'h21d == io_sel ? io_ins_541 : _GEN_540; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_542 = 10'h21e == io_sel ? io_ins_542 : _GEN_541; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_543 = 10'h21f == io_sel ? io_ins_543 : _GEN_542; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_544 = 10'h220 == io_sel ? io_ins_544 : _GEN_543; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_545 = 10'h221 == io_sel ? io_ins_545 : _GEN_544; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_546 = 10'h222 == io_sel ? io_ins_546 : _GEN_545; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_547 = 10'h223 == io_sel ? io_ins_547 : _GEN_546; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_548 = 10'h224 == io_sel ? io_ins_548 : _GEN_547; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_549 = 10'h225 == io_sel ? io_ins_549 : _GEN_548; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_550 = 10'h226 == io_sel ? io_ins_550 : _GEN_549; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_551 = 10'h227 == io_sel ? io_ins_551 : _GEN_550; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_552 = 10'h228 == io_sel ? io_ins_552 : _GEN_551; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_553 = 10'h229 == io_sel ? io_ins_553 : _GEN_552; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_554 = 10'h22a == io_sel ? io_ins_554 : _GEN_553; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_555 = 10'h22b == io_sel ? io_ins_555 : _GEN_554; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_556 = 10'h22c == io_sel ? io_ins_556 : _GEN_555; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_557 = 10'h22d == io_sel ? io_ins_557 : _GEN_556; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_558 = 10'h22e == io_sel ? io_ins_558 : _GEN_557; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_559 = 10'h22f == io_sel ? io_ins_559 : _GEN_558; // @[MuxN.scala 16:10:@140822.4]
  assign _GEN_560 = 10'h230 == io_sel ? io_ins_560 : _GEN_559; // @[MuxN.scala 16:10:@140822.4]
  assign io_out = 10'h231 == io_sel ? io_ins_561 : _GEN_560; // @[MuxN.scala 16:10:@140822.4]
endmodule
module RegFile( // @[:@140824.2]
  input         clock, // @[:@140825.4]
  input         reset, // @[:@140826.4]
  input  [10:0] io_raddr, // @[:@140827.4]
  input         io_wen, // @[:@140827.4]
  input  [10:0] io_waddr, // @[:@140827.4]
  input  [63:0] io_wdata, // @[:@140827.4]
  output [63:0] io_rdata, // @[:@140827.4]
  input         io_reset, // @[:@140827.4]
  output [63:0] io_argIns_0, // @[:@140827.4]
  output [63:0] io_argIns_1, // @[:@140827.4]
  output [63:0] io_argIns_2, // @[:@140827.4]
  output [63:0] io_argIns_3, // @[:@140827.4]
  input         io_argOuts_0_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_0_bits, // @[:@140827.4]
  input         io_argOuts_1_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_1_bits, // @[:@140827.4]
  input         io_argOuts_2_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_2_bits, // @[:@140827.4]
  input         io_argOuts_3_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_3_bits, // @[:@140827.4]
  input         io_argOuts_4_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_4_bits, // @[:@140827.4]
  input         io_argOuts_5_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_5_bits, // @[:@140827.4]
  input         io_argOuts_6_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_6_bits, // @[:@140827.4]
  input         io_argOuts_7_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_7_bits, // @[:@140827.4]
  input         io_argOuts_8_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_8_bits, // @[:@140827.4]
  input         io_argOuts_9_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_9_bits, // @[:@140827.4]
  input         io_argOuts_10_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_10_bits, // @[:@140827.4]
  input         io_argOuts_11_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_11_bits, // @[:@140827.4]
  input         io_argOuts_12_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_12_bits, // @[:@140827.4]
  input         io_argOuts_13_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_13_bits, // @[:@140827.4]
  input         io_argOuts_14_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_14_bits, // @[:@140827.4]
  input         io_argOuts_15_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_15_bits, // @[:@140827.4]
  input         io_argOuts_16_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_16_bits, // @[:@140827.4]
  input         io_argOuts_17_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_17_bits, // @[:@140827.4]
  input         io_argOuts_18_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_18_bits, // @[:@140827.4]
  input         io_argOuts_19_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_19_bits, // @[:@140827.4]
  input         io_argOuts_20_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_20_bits, // @[:@140827.4]
  input         io_argOuts_21_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_21_bits, // @[:@140827.4]
  input         io_argOuts_22_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_22_bits, // @[:@140827.4]
  input         io_argOuts_23_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_23_bits, // @[:@140827.4]
  input         io_argOuts_24_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_24_bits, // @[:@140827.4]
  input         io_argOuts_25_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_25_bits, // @[:@140827.4]
  input         io_argOuts_26_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_26_bits, // @[:@140827.4]
  input         io_argOuts_27_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_27_bits, // @[:@140827.4]
  input         io_argOuts_28_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_28_bits, // @[:@140827.4]
  input         io_argOuts_29_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_29_bits, // @[:@140827.4]
  input         io_argOuts_30_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_30_bits, // @[:@140827.4]
  input         io_argOuts_31_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_31_bits, // @[:@140827.4]
  input         io_argOuts_32_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_32_bits, // @[:@140827.4]
  input         io_argOuts_33_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_33_bits, // @[:@140827.4]
  input         io_argOuts_34_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_34_bits, // @[:@140827.4]
  input         io_argOuts_35_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_35_bits, // @[:@140827.4]
  input         io_argOuts_36_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_36_bits, // @[:@140827.4]
  input         io_argOuts_37_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_37_bits, // @[:@140827.4]
  input         io_argOuts_38_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_38_bits, // @[:@140827.4]
  input         io_argOuts_39_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_39_bits, // @[:@140827.4]
  input         io_argOuts_40_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_40_bits, // @[:@140827.4]
  input         io_argOuts_41_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_41_bits, // @[:@140827.4]
  input         io_argOuts_42_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_42_bits, // @[:@140827.4]
  input         io_argOuts_43_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_43_bits, // @[:@140827.4]
  input         io_argOuts_44_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_44_bits, // @[:@140827.4]
  input         io_argOuts_45_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_45_bits, // @[:@140827.4]
  input         io_argOuts_46_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_46_bits, // @[:@140827.4]
  input         io_argOuts_47_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_47_bits, // @[:@140827.4]
  input         io_argOuts_48_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_48_bits, // @[:@140827.4]
  input         io_argOuts_49_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_49_bits, // @[:@140827.4]
  input         io_argOuts_50_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_50_bits, // @[:@140827.4]
  input         io_argOuts_51_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_51_bits, // @[:@140827.4]
  input         io_argOuts_52_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_52_bits, // @[:@140827.4]
  input         io_argOuts_53_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_53_bits, // @[:@140827.4]
  input         io_argOuts_54_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_54_bits, // @[:@140827.4]
  input         io_argOuts_55_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_55_bits, // @[:@140827.4]
  input         io_argOuts_56_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_56_bits, // @[:@140827.4]
  input         io_argOuts_57_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_57_bits, // @[:@140827.4]
  input         io_argOuts_58_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_58_bits, // @[:@140827.4]
  input         io_argOuts_59_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_59_bits, // @[:@140827.4]
  input         io_argOuts_60_valid, // @[:@140827.4]
  input  [63:0] io_argOuts_60_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_61_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_62_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_63_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_64_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_65_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_66_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_67_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_68_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_69_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_70_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_71_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_72_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_73_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_74_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_75_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_76_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_77_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_78_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_79_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_80_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_81_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_82_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_83_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_84_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_85_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_86_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_87_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_88_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_89_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_90_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_91_bits, // @[:@140827.4]
  input  [63:0] io_argOuts_102_bits, // @[:@140827.4]
  output [63:0] io_argEchos_1, // @[:@140827.4]
  output [63:0] io_argEchos_2, // @[:@140827.4]
  output [63:0] io_argEchos_3, // @[:@140827.4]
  output [63:0] io_argEchos_4, // @[:@140827.4]
  output [63:0] io_argEchos_5, // @[:@140827.4]
  output [63:0] io_argEchos_6, // @[:@140827.4]
  output [63:0] io_argEchos_7, // @[:@140827.4]
  output [63:0] io_argEchos_8, // @[:@140827.4]
  output [63:0] io_argEchos_9, // @[:@140827.4]
  output [63:0] io_argEchos_10, // @[:@140827.4]
  output [63:0] io_argEchos_11, // @[:@140827.4]
  output [63:0] io_argEchos_12, // @[:@140827.4]
  output [63:0] io_argEchos_13, // @[:@140827.4]
  output [63:0] io_argEchos_14, // @[:@140827.4]
  output [63:0] io_argEchos_15, // @[:@140827.4]
  output [63:0] io_argEchos_16, // @[:@140827.4]
  output [63:0] io_argEchos_17, // @[:@140827.4]
  output [63:0] io_argEchos_18, // @[:@140827.4]
  output [63:0] io_argEchos_19, // @[:@140827.4]
  output [63:0] io_argEchos_20, // @[:@140827.4]
  output [63:0] io_argEchos_21, // @[:@140827.4]
  output [63:0] io_argEchos_22, // @[:@140827.4]
  output [63:0] io_argEchos_23, // @[:@140827.4]
  output [63:0] io_argEchos_24, // @[:@140827.4]
  output [63:0] io_argEchos_25, // @[:@140827.4]
  output [63:0] io_argEchos_26, // @[:@140827.4]
  output [63:0] io_argEchos_27, // @[:@140827.4]
  output [63:0] io_argEchos_28, // @[:@140827.4]
  output [63:0] io_argEchos_29, // @[:@140827.4]
  output [63:0] io_argEchos_30, // @[:@140827.4]
  output [63:0] io_argEchos_31, // @[:@140827.4]
  output [63:0] io_argEchos_32, // @[:@140827.4]
  output [63:0] io_argEchos_33, // @[:@140827.4]
  output [63:0] io_argEchos_34, // @[:@140827.4]
  output [63:0] io_argEchos_35, // @[:@140827.4]
  output [63:0] io_argEchos_36, // @[:@140827.4]
  output [63:0] io_argEchos_37, // @[:@140827.4]
  output [63:0] io_argEchos_38, // @[:@140827.4]
  output [63:0] io_argEchos_39, // @[:@140827.4]
  output [63:0] io_argEchos_40, // @[:@140827.4]
  output [63:0] io_argEchos_41, // @[:@140827.4]
  output [63:0] io_argEchos_42, // @[:@140827.4]
  output [63:0] io_argEchos_43, // @[:@140827.4]
  output [63:0] io_argEchos_44, // @[:@140827.4]
  output [63:0] io_argEchos_45, // @[:@140827.4]
  output [63:0] io_argEchos_46, // @[:@140827.4]
  output [63:0] io_argEchos_47, // @[:@140827.4]
  output [63:0] io_argEchos_48, // @[:@140827.4]
  output [63:0] io_argEchos_49, // @[:@140827.4]
  output [63:0] io_argEchos_50, // @[:@140827.4]
  output [63:0] io_argEchos_51, // @[:@140827.4]
  output [63:0] io_argEchos_52, // @[:@140827.4]
  output [63:0] io_argEchos_53, // @[:@140827.4]
  output [63:0] io_argEchos_54, // @[:@140827.4]
  output [63:0] io_argEchos_55, // @[:@140827.4]
  output [63:0] io_argEchos_56, // @[:@140827.4]
  output [63:0] io_argEchos_57, // @[:@140827.4]
  output [63:0] io_argEchos_58, // @[:@140827.4]
  output [63:0] io_argEchos_59, // @[:@140827.4]
  output [63:0] io_argEchos_60 // @[:@140827.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@143073.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@143073.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@143073.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@143073.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@143073.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@143073.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@143085.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@143085.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@143085.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@143085.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@143085.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@143085.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@143104.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@143104.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@143104.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@143104.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@143104.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@143104.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@143116.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@143116.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@143116.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@143116.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@143116.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@143116.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@143128.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@143128.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@143128.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@143128.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@143128.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@143128.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@143142.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@143142.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@143142.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@143142.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@143142.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@143142.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@143156.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@143156.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@143156.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@143156.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@143156.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@143156.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@143170.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@143170.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@143170.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@143170.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@143170.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@143170.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@143184.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@143184.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@143184.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@143184.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@143184.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@143184.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@143198.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@143198.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@143198.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@143198.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@143198.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@143198.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@143212.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@143212.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@143212.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@143212.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@143212.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@143212.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@143226.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@143226.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@143226.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@143226.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@143226.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@143226.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@143240.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@143240.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@143240.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@143240.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@143240.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@143240.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@143254.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@143254.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@143254.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@143254.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@143254.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@143254.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@143268.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@143268.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@143268.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@143268.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@143268.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@143268.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@143282.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@143282.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@143282.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@143282.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@143282.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@143282.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@143296.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@143296.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@143296.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@143296.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@143296.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@143296.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@143310.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@143310.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@143310.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@143310.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@143310.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@143310.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@143324.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@143324.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@143324.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@143324.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@143324.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@143324.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@143338.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@143338.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@143338.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@143338.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@143338.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@143338.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@143352.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@143352.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@143352.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@143352.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@143352.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@143352.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@143366.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@143366.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@143366.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@143366.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@143366.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@143366.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@143380.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@143380.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@143380.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@143380.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@143380.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@143380.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@143394.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@143394.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@143394.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@143394.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@143394.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@143394.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@143408.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@143408.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@143408.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@143408.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@143408.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@143408.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@143422.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@143422.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@143422.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@143422.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@143422.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@143422.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@143436.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@143436.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@143436.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@143436.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@143436.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@143436.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@143450.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@143450.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@143450.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@143450.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@143450.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@143450.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@143464.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@143464.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@143464.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@143464.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@143464.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@143464.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@143478.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@143478.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@143478.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@143478.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@143478.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@143478.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@143492.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@143492.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@143492.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@143492.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@143492.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@143492.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@143506.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@143506.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@143506.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@143506.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@143506.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@143506.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@143520.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@143520.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@143520.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@143520.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@143520.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@143520.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@143534.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@143534.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@143534.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@143534.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@143534.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@143534.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@143548.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@143548.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@143548.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@143548.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@143548.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@143548.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@143562.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@143562.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@143562.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@143562.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@143562.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@143562.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@143576.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@143576.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@143576.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@143576.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@143576.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@143576.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@143590.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@143590.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@143590.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@143590.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@143590.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@143590.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@143604.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@143604.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@143604.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@143604.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@143604.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@143604.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@143618.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@143618.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@143618.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@143618.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@143618.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@143618.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@143632.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@143632.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@143632.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@143632.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@143632.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@143632.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@143646.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@143646.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@143646.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@143646.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@143646.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@143646.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@143660.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@143660.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@143660.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@143660.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@143660.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@143660.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@143674.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@143674.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@143674.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@143674.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@143674.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@143674.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@143688.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@143688.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@143688.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@143688.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@143688.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@143688.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@143702.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@143702.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@143702.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@143702.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@143702.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@143702.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@143716.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@143716.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@143716.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@143716.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@143716.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@143716.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@143730.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@143730.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@143730.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@143730.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@143730.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@143730.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@143744.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@143744.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@143744.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@143744.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@143744.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@143744.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@143758.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@143758.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@143758.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@143758.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@143758.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@143758.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@143772.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@143772.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@143772.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@143772.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@143772.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@143772.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@143786.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@143786.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@143786.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@143786.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@143786.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@143786.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@143800.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@143800.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@143800.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@143800.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@143800.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@143800.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@143814.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@143814.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@143814.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@143814.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@143814.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@143814.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@143828.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@143828.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@143828.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@143828.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@143828.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@143828.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@143842.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@143842.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@143842.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@143842.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@143842.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@143842.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@143856.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@143856.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@143856.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@143856.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@143856.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@143856.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@143870.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@143870.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@143870.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@143870.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@143870.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@143870.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@143884.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@143884.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@143884.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@143884.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@143884.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@143884.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@143898.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@143898.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@143898.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@143898.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@143898.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@143898.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@143912.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@143912.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@143912.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@143912.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@143912.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@143912.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@143926.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@143926.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@143926.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@143926.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@143926.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@143926.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@143940.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@143940.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@143940.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@143940.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@143940.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@143940.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@143954.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@143954.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@143954.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@143954.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@143954.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@143954.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@143968.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@143968.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@143968.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@143968.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@143968.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@143968.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@143982.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@143982.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@143982.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@143982.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@143982.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@143982.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@143996.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@143996.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@143996.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@143996.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@143996.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@143996.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@144010.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@144010.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@144010.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@144010.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@144010.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@144010.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@144024.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@144024.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@144024.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@144024.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@144024.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@144024.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@144038.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@144038.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@144038.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@144038.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@144038.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@144038.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@144052.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@144052.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@144052.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@144052.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@144052.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@144052.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@144066.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@144066.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@144066.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@144066.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@144066.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@144066.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@144080.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@144080.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@144080.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@144080.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@144080.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@144080.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@144094.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@144094.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@144094.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@144094.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@144094.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@144094.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@144108.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@144108.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@144108.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@144108.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@144108.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@144108.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@144122.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@144122.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@144122.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@144122.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@144122.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@144122.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@144136.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@144136.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@144136.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@144136.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@144136.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@144136.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@144150.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@144150.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@144150.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@144150.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@144150.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@144150.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@144164.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@144164.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@144164.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@144164.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@144164.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@144164.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@144178.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@144178.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@144178.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@144178.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@144178.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@144178.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@144192.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@144192.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@144192.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@144192.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@144192.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@144192.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@144206.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@144206.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@144206.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@144206.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@144206.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@144206.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@144220.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@144220.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@144220.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@144220.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@144220.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@144220.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@144234.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@144234.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@144234.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@144234.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@144234.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@144234.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@144248.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@144248.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@144248.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@144248.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@144248.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@144248.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@144262.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@144262.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@144262.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@144262.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@144262.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@144262.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@144276.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@144276.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@144276.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@144276.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@144276.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@144276.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@144290.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@144290.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@144290.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@144290.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@144290.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@144290.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@144304.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@144304.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@144304.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@144304.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@144304.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@144304.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@144318.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@144318.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@144318.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@144318.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@144318.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@144318.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@144332.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@144332.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@144332.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@144332.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@144332.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@144332.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@144346.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@144346.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@144346.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@144346.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@144346.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@144346.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@144360.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@144360.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@144360.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@144360.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@144360.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@144360.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@144374.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@144374.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@144374.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@144374.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@144374.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@144374.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@144388.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@144388.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@144388.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@144388.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@144388.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@144388.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@144402.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@144402.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@144402.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@144402.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@144402.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@144402.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@144416.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@144416.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@144416.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@144416.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@144416.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@144416.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@144430.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@144430.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@144430.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@144430.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@144430.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@144430.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@144444.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@144444.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@144444.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@144444.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@144444.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@144444.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@144458.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@144458.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@144458.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@144458.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@144458.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@144458.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@144472.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@144472.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@144472.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@144472.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@144472.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@144472.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@144486.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@144486.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@144486.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@144486.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@144486.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@144486.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@144500.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@144500.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@144500.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@144500.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@144500.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@144500.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@144514.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@144514.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@144514.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@144514.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@144514.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@144514.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@144528.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@144528.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@144528.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@144528.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@144528.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@144528.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@144542.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@144542.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@144542.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@144542.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@144542.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@144542.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@144556.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@144556.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@144556.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@144556.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@144556.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@144556.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@144570.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@144570.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@144570.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@144570.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@144570.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@144570.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@144584.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@144584.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@144584.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@144584.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@144584.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@144584.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@144598.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@144598.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@144598.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@144598.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@144598.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@144598.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@144612.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@144612.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@144612.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@144612.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@144612.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@144612.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@144626.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@144626.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@144626.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@144626.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@144626.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@144626.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@144640.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@144640.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@144640.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@144640.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@144640.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@144640.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@144654.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@144654.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@144654.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@144654.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@144654.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@144654.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@144668.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@144668.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@144668.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@144668.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@144668.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@144668.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@144682.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@144682.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@144682.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@144682.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@144682.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@144682.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@144696.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@144696.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@144696.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@144696.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@144696.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@144696.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@144710.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@144710.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@144710.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@144710.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@144710.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@144710.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@144724.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@144724.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@144724.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@144724.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@144724.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@144724.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@144738.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@144738.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@144738.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@144738.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@144738.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@144738.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@144752.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@144752.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@144752.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@144752.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@144752.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@144752.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@144766.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@144766.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@144766.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@144766.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@144766.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@144766.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@144780.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@144780.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@144780.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@144780.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@144780.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@144780.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@144794.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@144794.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@144794.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@144794.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@144794.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@144794.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@144808.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@144808.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@144808.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@144808.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@144808.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@144808.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@144822.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@144822.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@144822.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@144822.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@144822.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@144822.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@144836.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@144836.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@144836.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@144836.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@144836.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@144836.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@144850.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@144850.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@144850.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@144850.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@144850.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@144850.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@144864.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@144864.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@144864.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@144864.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@144864.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@144864.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@144878.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@144878.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@144878.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@144878.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@144878.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@144878.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@144892.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@144892.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@144892.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@144892.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@144892.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@144892.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@144906.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@144906.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@144906.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@144906.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@144906.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@144906.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@144920.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@144920.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@144920.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@144920.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@144920.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@144920.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@144934.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@144934.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@144934.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@144934.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@144934.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@144934.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@144948.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@144948.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@144948.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@144948.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@144948.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@144948.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@144962.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@144962.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@144962.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@144962.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@144962.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@144962.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@144976.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@144976.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@144976.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@144976.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@144976.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@144976.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@144990.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@144990.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@144990.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@144990.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@144990.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@144990.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@145004.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@145004.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@145004.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@145004.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@145004.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@145004.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@145018.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@145018.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@145018.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@145018.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@145018.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@145018.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@145032.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@145032.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@145032.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@145032.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@145032.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@145032.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@145046.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@145046.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@145046.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@145046.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@145046.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@145046.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@145060.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@145060.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@145060.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@145060.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@145060.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@145060.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@145074.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@145074.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@145074.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@145074.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@145074.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@145074.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@145088.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@145088.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@145088.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@145088.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@145088.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@145088.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@145102.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@145102.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@145102.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@145102.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@145102.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@145102.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@145116.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@145116.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@145116.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@145116.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@145116.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@145116.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@145130.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@145130.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@145130.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@145130.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@145130.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@145130.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@145144.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@145144.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@145144.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@145144.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@145144.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@145144.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@145158.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@145158.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@145158.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@145158.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@145158.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@145158.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@145172.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@145172.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@145172.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@145172.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@145172.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@145172.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@145186.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@145186.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@145186.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@145186.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@145186.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@145186.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@145200.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@145200.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@145200.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@145200.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@145200.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@145200.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@145214.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@145214.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@145214.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@145214.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@145214.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@145214.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@145228.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@145228.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@145228.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@145228.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@145228.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@145228.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@145242.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@145242.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@145242.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@145242.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@145242.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@145242.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@145256.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@145256.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@145256.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@145256.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@145256.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@145256.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@145270.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@145270.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@145270.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@145270.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@145270.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@145270.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@145284.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@145284.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@145284.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@145284.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@145284.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@145284.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@145298.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@145298.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@145298.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@145298.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@145298.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@145298.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@145312.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@145312.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@145312.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@145312.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@145312.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@145312.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@145326.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@145326.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@145326.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@145326.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@145326.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@145326.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@145340.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@145340.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@145340.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@145340.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@145340.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@145340.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@145354.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@145354.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@145354.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@145354.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@145354.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@145354.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@145368.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@145368.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@145368.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@145368.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@145368.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@145368.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@145382.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@145382.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@145382.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@145382.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@145382.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@145382.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@145396.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@145396.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@145396.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@145396.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@145396.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@145396.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@145410.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@145410.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@145410.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@145410.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@145410.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@145410.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@145424.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@145424.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@145424.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@145424.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@145424.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@145424.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@145438.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@145438.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@145438.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@145438.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@145438.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@145438.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@145452.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@145452.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@145452.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@145452.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@145452.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@145452.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@145466.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@145466.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@145466.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@145466.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@145466.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@145466.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@145480.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@145480.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@145480.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@145480.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@145480.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@145480.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@145494.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@145494.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@145494.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@145494.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@145494.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@145494.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@145508.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@145508.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@145508.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@145508.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@145508.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@145508.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@145522.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@145522.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@145522.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@145522.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@145522.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@145522.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@145536.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@145536.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@145536.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@145536.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@145536.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@145536.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@145550.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@145550.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@145550.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@145550.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@145550.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@145550.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@145564.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@145564.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@145564.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@145564.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@145564.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@145564.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@145578.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@145578.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@145578.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@145578.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@145578.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@145578.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@145592.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@145592.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@145592.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@145592.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@145592.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@145592.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@145606.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@145606.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@145606.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@145606.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@145606.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@145606.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@145620.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@145620.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@145620.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@145620.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@145620.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@145620.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@145634.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@145634.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@145634.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@145634.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@145634.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@145634.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@145648.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@145648.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@145648.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@145648.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@145648.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@145648.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@145662.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@145662.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@145662.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@145662.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@145662.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@145662.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@145676.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@145676.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@145676.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@145676.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@145676.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@145676.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@145690.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@145690.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@145690.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@145690.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@145690.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@145690.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@145704.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@145704.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@145704.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@145704.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@145704.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@145704.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@145718.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@145718.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@145718.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@145718.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@145718.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@145718.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@145732.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@145732.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@145732.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@145732.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@145732.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@145732.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@145746.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@145746.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@145746.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@145746.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@145746.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@145746.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@145760.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@145760.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@145760.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@145760.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@145760.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@145760.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@145774.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@145774.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@145774.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@145774.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@145774.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@145774.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@145788.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@145788.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@145788.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@145788.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@145788.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@145788.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@145802.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@145802.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@145802.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@145802.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@145802.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@145802.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@145816.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@145816.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@145816.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@145816.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@145816.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@145816.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@145830.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@145830.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@145830.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@145830.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@145830.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@145830.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@145844.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@145844.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@145844.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@145844.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@145844.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@145844.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@145858.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@145858.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@145858.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@145858.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@145858.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@145858.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@145872.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@145872.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@145872.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@145872.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@145872.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@145872.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@145886.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@145886.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@145886.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@145886.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@145886.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@145886.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@145900.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@145900.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@145900.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@145900.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@145900.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@145900.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@145914.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@145914.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@145914.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@145914.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@145914.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@145914.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@145928.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@145928.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@145928.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@145928.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@145928.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@145928.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@145942.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@145942.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@145942.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@145942.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@145942.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@145942.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@145956.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@145956.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@145956.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@145956.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@145956.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@145956.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@145970.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@145970.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@145970.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@145970.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@145970.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@145970.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@145984.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@145984.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@145984.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@145984.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@145984.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@145984.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@145998.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@145998.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@145998.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@145998.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@145998.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@145998.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@146012.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@146012.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@146012.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@146012.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@146012.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@146012.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@146026.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@146026.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@146026.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@146026.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@146026.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@146026.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@146040.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@146040.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@146040.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@146040.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@146040.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@146040.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@146054.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@146054.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@146054.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@146054.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@146054.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@146054.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@146068.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@146068.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@146068.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@146068.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@146068.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@146068.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@146082.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@146082.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@146082.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@146082.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@146082.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@146082.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@146096.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@146096.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@146096.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@146096.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@146096.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@146096.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@146110.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@146110.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@146110.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@146110.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@146110.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@146110.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@146124.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@146124.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@146124.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@146124.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@146124.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@146124.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@146138.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@146138.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@146138.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@146138.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@146138.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@146138.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@146152.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@146152.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@146152.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@146152.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@146152.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@146152.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@146166.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@146166.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@146166.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@146166.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@146166.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@146166.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@146180.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@146180.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@146180.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@146180.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@146180.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@146180.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@146194.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@146194.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@146194.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@146194.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@146194.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@146194.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@146208.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@146208.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@146208.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@146208.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@146208.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@146208.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@146222.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@146222.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@146222.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@146222.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@146222.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@146222.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@146236.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@146236.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@146236.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@146236.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@146236.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@146236.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@146250.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@146250.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@146250.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@146250.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@146250.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@146250.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@146264.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@146264.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@146264.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@146264.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@146264.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@146264.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@146278.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@146278.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@146278.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@146278.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@146278.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@146278.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@146292.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@146292.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@146292.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@146292.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@146292.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@146292.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@146306.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@146306.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@146306.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@146306.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@146306.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@146306.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@146320.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@146320.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@146320.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@146320.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@146320.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@146320.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@146334.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@146334.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@146334.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@146334.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@146334.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@146334.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@146348.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@146348.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@146348.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@146348.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@146348.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@146348.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@146362.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@146362.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@146362.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@146362.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@146362.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@146362.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@146376.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@146376.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@146376.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@146376.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@146376.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@146376.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@146390.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@146390.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@146390.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@146390.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@146390.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@146390.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@146404.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@146404.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@146404.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@146404.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@146404.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@146404.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@146418.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@146418.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@146418.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@146418.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@146418.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@146418.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@146432.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@146432.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@146432.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@146432.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@146432.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@146432.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@146446.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@146446.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@146446.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@146446.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@146446.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@146446.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@146460.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@146460.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@146460.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@146460.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@146460.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@146460.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@146474.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@146474.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@146474.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@146474.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@146474.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@146474.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@146488.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@146488.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@146488.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@146488.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@146488.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@146488.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@146502.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@146502.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@146502.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@146502.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@146502.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@146502.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@146516.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@146516.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@146516.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@146516.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@146516.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@146516.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@146530.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@146530.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@146530.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@146530.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@146530.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@146530.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@146544.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@146544.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@146544.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@146544.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@146544.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@146544.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@146558.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@146558.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@146558.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@146558.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@146558.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@146558.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@146572.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@146572.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@146572.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@146572.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@146572.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@146572.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@146586.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@146586.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@146586.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@146586.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@146586.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@146586.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@146600.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@146600.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@146600.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@146600.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@146600.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@146600.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@146614.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@146614.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@146614.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@146614.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@146614.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@146614.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@146628.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@146628.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@146628.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@146628.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@146628.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@146628.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@146642.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@146642.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@146642.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@146642.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@146642.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@146642.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@146656.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@146656.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@146656.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@146656.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@146656.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@146656.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@146670.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@146670.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@146670.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@146670.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@146670.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@146670.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@146684.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@146684.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@146684.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@146684.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@146684.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@146684.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@146698.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@146698.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@146698.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@146698.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@146698.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@146698.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@146712.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@146712.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@146712.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@146712.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@146712.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@146712.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@146726.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@146726.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@146726.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@146726.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@146726.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@146726.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@146740.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@146740.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@146740.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@146740.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@146740.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@146740.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@146754.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@146754.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@146754.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@146754.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@146754.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@146754.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@146768.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@146768.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@146768.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@146768.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@146768.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@146768.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@146782.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@146782.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@146782.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@146782.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@146782.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@146782.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@146796.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@146796.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@146796.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@146796.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@146796.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@146796.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@146810.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@146810.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@146810.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@146810.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@146810.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@146810.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@146824.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@146824.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@146824.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@146824.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@146824.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@146824.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@146838.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@146838.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@146838.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@146838.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@146838.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@146838.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@146852.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@146852.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@146852.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@146852.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@146852.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@146852.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@146866.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@146866.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@146866.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@146866.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@146866.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@146866.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@146880.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@146880.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@146880.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@146880.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@146880.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@146880.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@146894.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@146894.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@146894.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@146894.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@146894.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@146894.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@146908.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@146908.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@146908.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@146908.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@146908.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@146908.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@146922.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@146922.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@146922.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@146922.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@146922.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@146922.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@146936.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@146936.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@146936.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@146936.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@146936.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@146936.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@146950.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@146950.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@146950.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@146950.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@146950.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@146950.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@146964.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@146964.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@146964.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@146964.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@146964.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@146964.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@146978.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@146978.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@146978.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@146978.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@146978.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@146978.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@146992.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@146992.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@146992.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@146992.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@146992.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@146992.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@147006.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@147006.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@147006.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@147006.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@147006.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@147006.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@147020.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@147020.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@147020.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@147020.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@147020.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@147020.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@147034.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@147034.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@147034.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@147034.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@147034.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@147034.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@147048.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@147048.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@147048.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@147048.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@147048.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@147048.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@147062.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@147062.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@147062.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@147062.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@147062.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@147062.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@147076.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@147076.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@147076.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@147076.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@147076.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@147076.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@147090.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@147090.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@147090.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@147090.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@147090.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@147090.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@147104.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@147104.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@147104.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@147104.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@147104.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@147104.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@147118.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@147118.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@147118.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@147118.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@147118.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@147118.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@147132.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@147132.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@147132.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@147132.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@147132.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@147132.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@147146.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@147146.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@147146.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@147146.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@147146.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@147146.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@147160.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@147160.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@147160.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@147160.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@147160.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@147160.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@147174.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@147174.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@147174.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@147174.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@147174.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@147174.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@147188.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@147188.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@147188.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@147188.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@147188.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@147188.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@147202.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@147202.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@147202.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@147202.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@147202.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@147202.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@147216.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@147216.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@147216.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@147216.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@147216.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@147216.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@147230.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@147230.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@147230.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@147230.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@147230.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@147230.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@147244.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@147244.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@147244.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@147244.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@147244.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@147244.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@147258.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@147258.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@147258.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@147258.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@147258.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@147258.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@147272.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@147272.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@147272.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@147272.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@147272.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@147272.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@147286.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@147286.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@147286.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@147286.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@147286.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@147286.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@147300.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@147300.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@147300.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@147300.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@147300.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@147300.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@147314.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@147314.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@147314.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@147314.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@147314.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@147314.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@147328.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@147328.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@147328.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@147328.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@147328.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@147328.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@147342.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@147342.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@147342.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@147342.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@147342.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@147342.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@147356.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@147356.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@147356.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@147356.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@147356.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@147356.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@147370.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@147370.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@147370.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@147370.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@147370.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@147370.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@147384.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@147384.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@147384.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@147384.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@147384.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@147384.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@147398.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@147398.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@147398.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@147398.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@147398.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@147398.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@147412.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@147412.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@147412.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@147412.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@147412.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@147412.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@147426.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@147426.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@147426.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@147426.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@147426.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@147426.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@147440.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@147440.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@147440.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@147440.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@147440.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@147440.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@147454.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@147454.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@147454.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@147454.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@147454.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@147454.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@147468.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@147468.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@147468.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@147468.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@147468.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@147468.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@147482.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@147482.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@147482.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@147482.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@147482.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@147482.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@147496.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@147496.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@147496.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@147496.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@147496.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@147496.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@147510.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@147510.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@147510.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@147510.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@147510.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@147510.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@147524.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@147524.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@147524.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@147524.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@147524.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@147524.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@147538.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@147538.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@147538.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@147538.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@147538.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@147538.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@147552.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@147552.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@147552.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@147552.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@147552.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@147552.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@147566.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@147566.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@147566.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@147566.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@147566.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@147566.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@147580.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@147580.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@147580.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@147580.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@147580.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@147580.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@147594.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@147594.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@147594.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@147594.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@147594.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@147594.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@147608.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@147608.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@147608.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@147608.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@147608.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@147608.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@147622.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@147622.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@147622.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@147622.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@147622.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@147622.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@147636.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@147636.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@147636.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@147636.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@147636.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@147636.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@147650.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@147650.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@147650.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@147650.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@147650.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@147650.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@147664.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@147664.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@147664.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@147664.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@147664.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@147664.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@147678.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@147678.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@147678.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@147678.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@147678.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@147678.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@147692.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@147692.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@147692.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@147692.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@147692.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@147692.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@147706.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@147706.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@147706.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@147706.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@147706.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@147706.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@147720.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@147720.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@147720.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@147720.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@147720.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@147720.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@147734.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@147734.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@147734.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@147734.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@147734.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@147734.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@147748.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@147748.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@147748.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@147748.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@147748.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@147748.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@147762.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@147762.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@147762.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@147762.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@147762.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@147762.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@147776.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@147776.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@147776.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@147776.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@147776.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@147776.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@147790.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@147790.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@147790.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@147790.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@147790.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@147790.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@147804.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@147804.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@147804.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@147804.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@147804.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@147804.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@147818.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@147818.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@147818.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@147818.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@147818.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@147818.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@147832.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@147832.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@147832.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@147832.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@147832.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@147832.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@147846.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@147846.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@147846.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@147846.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@147846.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@147846.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@147860.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@147860.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@147860.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@147860.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@147860.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@147860.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@147874.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@147874.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@147874.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@147874.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@147874.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@147874.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@147888.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@147888.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@147888.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@147888.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@147888.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@147888.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@147902.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@147902.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@147902.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@147902.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@147902.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@147902.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@147916.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@147916.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@147916.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@147916.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@147916.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@147916.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@147930.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@147930.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@147930.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@147930.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@147930.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@147930.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@147944.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@147944.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@147944.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@147944.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@147944.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@147944.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@147958.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@147958.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@147958.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@147958.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@147958.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@147958.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@147972.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@147972.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@147972.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@147972.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@147972.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@147972.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@147986.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@147986.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@147986.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@147986.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@147986.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@147986.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@148000.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@148000.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@148000.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@148000.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@148000.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@148000.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@148014.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@148014.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@148014.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@148014.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@148014.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@148014.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@148028.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@148028.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@148028.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@148028.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@148028.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@148028.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@148042.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@148042.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@148042.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@148042.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@148042.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@148042.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@148056.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@148056.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@148056.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@148056.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@148056.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@148056.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@148070.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@148070.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@148070.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@148070.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@148070.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@148070.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@148084.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@148084.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@148084.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@148084.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@148084.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@148084.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@148098.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@148098.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@148098.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@148098.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@148098.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@148098.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@148112.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@148112.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@148112.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@148112.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@148112.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@148112.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@148126.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@148126.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@148126.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@148126.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@148126.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@148126.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@148140.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@148140.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@148140.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@148140.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@148140.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@148140.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@148154.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@148154.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@148154.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@148154.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@148154.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@148154.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@148168.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@148168.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@148168.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@148168.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@148168.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@148168.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@148182.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@148182.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@148182.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@148182.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@148182.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@148182.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@148196.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@148196.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@148196.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@148196.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@148196.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@148196.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@148210.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@148210.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@148210.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@148210.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@148210.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@148210.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@148224.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@148224.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@148224.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@148224.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@148224.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@148224.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@148238.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@148238.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@148238.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@148238.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@148238.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@148238.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@148252.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@148252.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@148252.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@148252.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@148252.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@148252.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@148266.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@148266.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@148266.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@148266.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@148266.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@148266.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@148280.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@148280.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@148280.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@148280.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@148280.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@148280.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@148294.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@148294.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@148294.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@148294.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@148294.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@148294.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@148308.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@148308.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@148308.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@148308.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@148308.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@148308.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@148322.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@148322.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@148322.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@148322.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@148322.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@148322.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@148336.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@148336.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@148336.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@148336.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@148336.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@148336.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@148350.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@148350.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@148350.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@148350.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@148350.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@148350.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@148364.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@148364.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@148364.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@148364.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@148364.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@148364.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@148378.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@148378.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@148378.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@148378.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@148378.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@148378.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@148392.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@148392.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@148392.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@148392.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@148392.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@148392.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@148406.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@148406.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@148406.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@148406.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@148406.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@148406.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@148420.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@148420.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@148420.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@148420.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@148420.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@148420.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@148434.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@148434.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@148434.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@148434.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@148434.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@148434.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@148448.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@148448.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@148448.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@148448.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@148448.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@148448.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@148462.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@148462.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@148462.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@148462.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@148462.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@148462.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@148476.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@148476.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@148476.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@148476.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@148476.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@148476.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@148490.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@148490.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@148490.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@148490.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@148490.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@148490.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@148504.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@148504.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@148504.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@148504.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@148504.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@148504.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@148518.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@148518.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@148518.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@148518.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@148518.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@148518.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@148532.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@148532.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@148532.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@148532.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@148532.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@148532.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@148546.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@148546.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@148546.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@148546.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@148546.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@148546.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@148560.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@148560.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@148560.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@148560.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@148560.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@148560.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@148574.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@148574.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@148574.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@148574.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@148574.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@148574.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@148588.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@148588.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@148588.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@148588.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@148588.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@148588.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@148602.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@148602.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@148602.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@148602.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@148602.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@148602.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@148616.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@148616.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@148616.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@148616.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@148616.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@148616.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@148630.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@148630.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@148630.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@148630.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@148630.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@148630.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@148644.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@148644.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@148644.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@148644.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@148644.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@148644.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@148658.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@148658.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@148658.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@148658.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@148658.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@148658.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@148672.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@148672.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@148672.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@148672.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@148672.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@148672.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@148686.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@148686.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@148686.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@148686.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@148686.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@148686.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@148700.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@148700.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@148700.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@148700.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@148700.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@148700.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@148714.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@148714.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@148714.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@148714.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@148714.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@148714.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@148728.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@148728.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@148728.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@148728.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@148728.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@148728.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@148742.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@148742.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@148742.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@148742.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@148742.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@148742.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@148756.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@148756.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@148756.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@148756.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@148756.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@148756.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@148770.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@148770.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@148770.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@148770.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@148770.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@148770.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@148784.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@148784.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@148784.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@148784.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@148784.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@148784.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@148798.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@148798.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@148798.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@148798.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@148798.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@148798.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@148812.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@148812.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@148812.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@148812.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@148812.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@148812.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@148826.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@148826.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@148826.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@148826.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@148826.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@148826.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@148840.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@148840.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@148840.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@148840.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@148840.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@148840.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@148854.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@148854.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@148854.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@148854.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@148854.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@148854.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@148868.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@148868.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@148868.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@148868.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@148868.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@148868.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@148882.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@148882.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@148882.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@148882.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@148882.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@148882.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@148896.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@148896.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@148896.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@148896.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@148896.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@148896.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@148910.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@148910.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@148910.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@148910.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@148910.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@148910.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@148924.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@148924.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@148924.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@148924.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@148924.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@148924.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@148938.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@148938.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@148938.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@148938.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@148938.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@148938.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@148952.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@148952.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@148952.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@148952.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@148952.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@148952.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@148966.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@148966.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@148966.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@148966.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@148966.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@148966.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@148980.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@148980.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@148980.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@148980.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@148980.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@148980.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@148994.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@148994.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@148994.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@148994.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@148994.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@148994.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@149008.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@149008.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@149008.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@149008.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@149008.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@149008.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@149022.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@149022.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@149022.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@149022.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@149022.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@149022.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@149036.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@149036.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@149036.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@149036.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@149036.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@149036.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@149050.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@149050.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@149050.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@149050.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@149050.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@149050.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@149064.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@149064.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@149064.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@149064.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@149064.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@149064.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@149078.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@149078.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@149078.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@149078.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@149078.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@149078.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@149092.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@149092.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@149092.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@149092.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@149092.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@149092.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@149106.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@149106.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@149106.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@149106.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@149106.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@149106.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@149120.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@149120.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@149120.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@149120.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@149120.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@149120.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@149134.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@149134.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@149134.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@149134.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@149134.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@149134.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@149148.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@149148.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@149148.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@149148.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@149148.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@149148.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@149162.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@149162.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@149162.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@149162.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@149162.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@149162.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@149176.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@149176.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@149176.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@149176.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@149176.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@149176.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@149190.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@149190.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@149190.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@149190.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@149190.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@149190.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@149204.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@149204.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@149204.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@149204.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@149204.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@149204.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@149218.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@149218.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@149218.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@149218.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@149218.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@149218.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@149232.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@149232.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@149232.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@149232.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@149232.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@149232.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@149246.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@149246.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@149246.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@149246.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@149246.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@149246.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@149260.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@149260.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@149260.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@149260.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@149260.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@149260.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@149274.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@149274.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@149274.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@149274.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@149274.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@149274.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@149288.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@149288.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@149288.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@149288.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@149288.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@149288.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@149302.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@149302.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@149302.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@149302.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@149302.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@149302.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@149316.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@149316.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@149316.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@149316.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@149316.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@149316.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@149330.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@149330.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@149330.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@149330.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@149330.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@149330.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@149344.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@149344.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@149344.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@149344.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@149344.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@149344.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@149358.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@149358.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@149358.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@149358.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@149358.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@149358.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@149372.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@149372.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@149372.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@149372.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@149372.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@149372.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@149386.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@149386.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@149386.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@149386.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@149386.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@149386.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@149400.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@149400.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@149400.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@149400.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@149400.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@149400.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@149414.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@149414.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@149414.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@149414.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@149414.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@149414.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@149428.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@149428.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@149428.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@149428.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@149428.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@149428.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@149442.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@149442.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@149442.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@149442.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@149442.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@149442.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@149456.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@149456.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@149456.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@149456.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@149456.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@149456.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@149470.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@149470.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@149470.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@149470.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@149470.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@149470.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@149484.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@149484.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@149484.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@149484.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@149484.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@149484.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@149498.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@149498.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@149498.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@149498.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@149498.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@149498.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@149512.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@149512.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@149512.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@149512.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@149512.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@149512.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@149526.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@149526.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@149526.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@149526.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@149526.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@149526.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@149540.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@149540.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@149540.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@149540.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@149540.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@149540.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@149554.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@149554.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@149554.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@149554.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@149554.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@149554.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@149568.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@149568.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@149568.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@149568.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@149568.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@149568.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@149582.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@149582.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@149582.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@149582.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@149582.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@149582.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@149596.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@149596.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@149596.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@149596.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@149596.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@149596.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@149610.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@149610.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@149610.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@149610.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@149610.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@149610.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@149624.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@149624.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@149624.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@149624.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@149624.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@149624.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@149638.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@149638.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@149638.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@149638.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@149638.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@149638.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@149652.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@149652.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@149652.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@149652.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@149652.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@149652.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@149666.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@149666.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@149666.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@149666.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@149666.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@149666.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@149680.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@149680.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@149680.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@149680.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@149680.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@149680.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@149694.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@149694.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@149694.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@149694.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@149694.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@149694.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@149708.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@149708.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@149708.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@149708.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@149708.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@149708.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@149722.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@149722.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@149722.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@149722.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@149722.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@149722.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@149736.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@149736.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@149736.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@149736.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@149736.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@149736.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@149750.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@149750.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@149750.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@149750.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@149750.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@149750.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@149764.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@149764.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@149764.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@149764.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@149764.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@149764.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@149778.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@149778.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@149778.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@149778.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@149778.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@149778.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@149792.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@149792.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@149792.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@149792.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@149792.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@149792.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@149806.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@149806.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@149806.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@149806.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@149806.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@149806.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@149820.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@149820.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@149820.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@149820.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@149820.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@149820.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@149834.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@149834.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@149834.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@149834.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@149834.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@149834.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@149848.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@149848.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@149848.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@149848.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@149848.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@149848.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@149862.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@149862.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@149862.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@149862.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@149862.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@149862.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@149876.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@149876.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@149876.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@149876.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@149876.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@149876.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@149890.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@149890.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@149890.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@149890.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@149890.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@149890.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@149904.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@149904.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@149904.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@149904.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@149904.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@149904.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@149918.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@149918.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@149918.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@149918.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@149918.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@149918.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@149932.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@149932.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@149932.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@149932.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@149932.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@149932.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@149946.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@149946.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@149946.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@149946.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@149946.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@149946.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@149960.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@149960.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@149960.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@149960.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@149960.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@149960.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@149974.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@149974.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@149974.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@149974.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@149974.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@149974.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@149988.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@149988.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@149988.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@149988.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@149988.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@149988.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@150002.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@150002.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@150002.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@150002.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@150002.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@150002.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@150016.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@150016.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@150016.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@150016.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@150016.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@150016.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@150030.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@150030.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@150030.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@150030.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@150030.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@150030.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@150044.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@150044.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@150044.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@150044.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@150044.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@150044.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@150058.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@150058.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@150058.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@150058.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@150058.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@150058.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@150072.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@150072.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@150072.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@150072.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@150072.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@150072.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@150086.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@150086.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@150086.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@150086.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@150086.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@150086.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@150100.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@150100.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@150100.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@150100.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@150100.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@150100.4]
  wire  regs_503_clock; // @[RegFile.scala 66:20:@150114.4]
  wire  regs_503_reset; // @[RegFile.scala 66:20:@150114.4]
  wire [63:0] regs_503_io_in; // @[RegFile.scala 66:20:@150114.4]
  wire  regs_503_io_reset; // @[RegFile.scala 66:20:@150114.4]
  wire [63:0] regs_503_io_out; // @[RegFile.scala 66:20:@150114.4]
  wire  regs_503_io_enable; // @[RegFile.scala 66:20:@150114.4]
  wire  regs_504_clock; // @[RegFile.scala 66:20:@150128.4]
  wire  regs_504_reset; // @[RegFile.scala 66:20:@150128.4]
  wire [63:0] regs_504_io_in; // @[RegFile.scala 66:20:@150128.4]
  wire  regs_504_io_reset; // @[RegFile.scala 66:20:@150128.4]
  wire [63:0] regs_504_io_out; // @[RegFile.scala 66:20:@150128.4]
  wire  regs_504_io_enable; // @[RegFile.scala 66:20:@150128.4]
  wire  regs_505_clock; // @[RegFile.scala 66:20:@150142.4]
  wire  regs_505_reset; // @[RegFile.scala 66:20:@150142.4]
  wire [63:0] regs_505_io_in; // @[RegFile.scala 66:20:@150142.4]
  wire  regs_505_io_reset; // @[RegFile.scala 66:20:@150142.4]
  wire [63:0] regs_505_io_out; // @[RegFile.scala 66:20:@150142.4]
  wire  regs_505_io_enable; // @[RegFile.scala 66:20:@150142.4]
  wire  regs_506_clock; // @[RegFile.scala 66:20:@150156.4]
  wire  regs_506_reset; // @[RegFile.scala 66:20:@150156.4]
  wire [63:0] regs_506_io_in; // @[RegFile.scala 66:20:@150156.4]
  wire  regs_506_io_reset; // @[RegFile.scala 66:20:@150156.4]
  wire [63:0] regs_506_io_out; // @[RegFile.scala 66:20:@150156.4]
  wire  regs_506_io_enable; // @[RegFile.scala 66:20:@150156.4]
  wire  regs_507_clock; // @[RegFile.scala 66:20:@150170.4]
  wire  regs_507_reset; // @[RegFile.scala 66:20:@150170.4]
  wire [63:0] regs_507_io_in; // @[RegFile.scala 66:20:@150170.4]
  wire  regs_507_io_reset; // @[RegFile.scala 66:20:@150170.4]
  wire [63:0] regs_507_io_out; // @[RegFile.scala 66:20:@150170.4]
  wire  regs_507_io_enable; // @[RegFile.scala 66:20:@150170.4]
  wire  regs_508_clock; // @[RegFile.scala 66:20:@150184.4]
  wire  regs_508_reset; // @[RegFile.scala 66:20:@150184.4]
  wire [63:0] regs_508_io_in; // @[RegFile.scala 66:20:@150184.4]
  wire  regs_508_io_reset; // @[RegFile.scala 66:20:@150184.4]
  wire [63:0] regs_508_io_out; // @[RegFile.scala 66:20:@150184.4]
  wire  regs_508_io_enable; // @[RegFile.scala 66:20:@150184.4]
  wire  regs_509_clock; // @[RegFile.scala 66:20:@150198.4]
  wire  regs_509_reset; // @[RegFile.scala 66:20:@150198.4]
  wire [63:0] regs_509_io_in; // @[RegFile.scala 66:20:@150198.4]
  wire  regs_509_io_reset; // @[RegFile.scala 66:20:@150198.4]
  wire [63:0] regs_509_io_out; // @[RegFile.scala 66:20:@150198.4]
  wire  regs_509_io_enable; // @[RegFile.scala 66:20:@150198.4]
  wire  regs_510_clock; // @[RegFile.scala 66:20:@150212.4]
  wire  regs_510_reset; // @[RegFile.scala 66:20:@150212.4]
  wire [63:0] regs_510_io_in; // @[RegFile.scala 66:20:@150212.4]
  wire  regs_510_io_reset; // @[RegFile.scala 66:20:@150212.4]
  wire [63:0] regs_510_io_out; // @[RegFile.scala 66:20:@150212.4]
  wire  regs_510_io_enable; // @[RegFile.scala 66:20:@150212.4]
  wire  regs_511_clock; // @[RegFile.scala 66:20:@150226.4]
  wire  regs_511_reset; // @[RegFile.scala 66:20:@150226.4]
  wire [63:0] regs_511_io_in; // @[RegFile.scala 66:20:@150226.4]
  wire  regs_511_io_reset; // @[RegFile.scala 66:20:@150226.4]
  wire [63:0] regs_511_io_out; // @[RegFile.scala 66:20:@150226.4]
  wire  regs_511_io_enable; // @[RegFile.scala 66:20:@150226.4]
  wire  regs_512_clock; // @[RegFile.scala 66:20:@150240.4]
  wire  regs_512_reset; // @[RegFile.scala 66:20:@150240.4]
  wire [63:0] regs_512_io_in; // @[RegFile.scala 66:20:@150240.4]
  wire  regs_512_io_reset; // @[RegFile.scala 66:20:@150240.4]
  wire [63:0] regs_512_io_out; // @[RegFile.scala 66:20:@150240.4]
  wire  regs_512_io_enable; // @[RegFile.scala 66:20:@150240.4]
  wire  regs_513_clock; // @[RegFile.scala 66:20:@150254.4]
  wire  regs_513_reset; // @[RegFile.scala 66:20:@150254.4]
  wire [63:0] regs_513_io_in; // @[RegFile.scala 66:20:@150254.4]
  wire  regs_513_io_reset; // @[RegFile.scala 66:20:@150254.4]
  wire [63:0] regs_513_io_out; // @[RegFile.scala 66:20:@150254.4]
  wire  regs_513_io_enable; // @[RegFile.scala 66:20:@150254.4]
  wire  regs_514_clock; // @[RegFile.scala 66:20:@150268.4]
  wire  regs_514_reset; // @[RegFile.scala 66:20:@150268.4]
  wire [63:0] regs_514_io_in; // @[RegFile.scala 66:20:@150268.4]
  wire  regs_514_io_reset; // @[RegFile.scala 66:20:@150268.4]
  wire [63:0] regs_514_io_out; // @[RegFile.scala 66:20:@150268.4]
  wire  regs_514_io_enable; // @[RegFile.scala 66:20:@150268.4]
  wire  regs_515_clock; // @[RegFile.scala 66:20:@150282.4]
  wire  regs_515_reset; // @[RegFile.scala 66:20:@150282.4]
  wire [63:0] regs_515_io_in; // @[RegFile.scala 66:20:@150282.4]
  wire  regs_515_io_reset; // @[RegFile.scala 66:20:@150282.4]
  wire [63:0] regs_515_io_out; // @[RegFile.scala 66:20:@150282.4]
  wire  regs_515_io_enable; // @[RegFile.scala 66:20:@150282.4]
  wire  regs_516_clock; // @[RegFile.scala 66:20:@150296.4]
  wire  regs_516_reset; // @[RegFile.scala 66:20:@150296.4]
  wire [63:0] regs_516_io_in; // @[RegFile.scala 66:20:@150296.4]
  wire  regs_516_io_reset; // @[RegFile.scala 66:20:@150296.4]
  wire [63:0] regs_516_io_out; // @[RegFile.scala 66:20:@150296.4]
  wire  regs_516_io_enable; // @[RegFile.scala 66:20:@150296.4]
  wire  regs_517_clock; // @[RegFile.scala 66:20:@150310.4]
  wire  regs_517_reset; // @[RegFile.scala 66:20:@150310.4]
  wire [63:0] regs_517_io_in; // @[RegFile.scala 66:20:@150310.4]
  wire  regs_517_io_reset; // @[RegFile.scala 66:20:@150310.4]
  wire [63:0] regs_517_io_out; // @[RegFile.scala 66:20:@150310.4]
  wire  regs_517_io_enable; // @[RegFile.scala 66:20:@150310.4]
  wire  regs_518_clock; // @[RegFile.scala 66:20:@150324.4]
  wire  regs_518_reset; // @[RegFile.scala 66:20:@150324.4]
  wire [63:0] regs_518_io_in; // @[RegFile.scala 66:20:@150324.4]
  wire  regs_518_io_reset; // @[RegFile.scala 66:20:@150324.4]
  wire [63:0] regs_518_io_out; // @[RegFile.scala 66:20:@150324.4]
  wire  regs_518_io_enable; // @[RegFile.scala 66:20:@150324.4]
  wire  regs_519_clock; // @[RegFile.scala 66:20:@150338.4]
  wire  regs_519_reset; // @[RegFile.scala 66:20:@150338.4]
  wire [63:0] regs_519_io_in; // @[RegFile.scala 66:20:@150338.4]
  wire  regs_519_io_reset; // @[RegFile.scala 66:20:@150338.4]
  wire [63:0] regs_519_io_out; // @[RegFile.scala 66:20:@150338.4]
  wire  regs_519_io_enable; // @[RegFile.scala 66:20:@150338.4]
  wire  regs_520_clock; // @[RegFile.scala 66:20:@150352.4]
  wire  regs_520_reset; // @[RegFile.scala 66:20:@150352.4]
  wire [63:0] regs_520_io_in; // @[RegFile.scala 66:20:@150352.4]
  wire  regs_520_io_reset; // @[RegFile.scala 66:20:@150352.4]
  wire [63:0] regs_520_io_out; // @[RegFile.scala 66:20:@150352.4]
  wire  regs_520_io_enable; // @[RegFile.scala 66:20:@150352.4]
  wire  regs_521_clock; // @[RegFile.scala 66:20:@150366.4]
  wire  regs_521_reset; // @[RegFile.scala 66:20:@150366.4]
  wire [63:0] regs_521_io_in; // @[RegFile.scala 66:20:@150366.4]
  wire  regs_521_io_reset; // @[RegFile.scala 66:20:@150366.4]
  wire [63:0] regs_521_io_out; // @[RegFile.scala 66:20:@150366.4]
  wire  regs_521_io_enable; // @[RegFile.scala 66:20:@150366.4]
  wire  regs_522_clock; // @[RegFile.scala 66:20:@150380.4]
  wire  regs_522_reset; // @[RegFile.scala 66:20:@150380.4]
  wire [63:0] regs_522_io_in; // @[RegFile.scala 66:20:@150380.4]
  wire  regs_522_io_reset; // @[RegFile.scala 66:20:@150380.4]
  wire [63:0] regs_522_io_out; // @[RegFile.scala 66:20:@150380.4]
  wire  regs_522_io_enable; // @[RegFile.scala 66:20:@150380.4]
  wire  regs_523_clock; // @[RegFile.scala 66:20:@150394.4]
  wire  regs_523_reset; // @[RegFile.scala 66:20:@150394.4]
  wire [63:0] regs_523_io_in; // @[RegFile.scala 66:20:@150394.4]
  wire  regs_523_io_reset; // @[RegFile.scala 66:20:@150394.4]
  wire [63:0] regs_523_io_out; // @[RegFile.scala 66:20:@150394.4]
  wire  regs_523_io_enable; // @[RegFile.scala 66:20:@150394.4]
  wire  regs_524_clock; // @[RegFile.scala 66:20:@150408.4]
  wire  regs_524_reset; // @[RegFile.scala 66:20:@150408.4]
  wire [63:0] regs_524_io_in; // @[RegFile.scala 66:20:@150408.4]
  wire  regs_524_io_reset; // @[RegFile.scala 66:20:@150408.4]
  wire [63:0] regs_524_io_out; // @[RegFile.scala 66:20:@150408.4]
  wire  regs_524_io_enable; // @[RegFile.scala 66:20:@150408.4]
  wire  regs_525_clock; // @[RegFile.scala 66:20:@150422.4]
  wire  regs_525_reset; // @[RegFile.scala 66:20:@150422.4]
  wire [63:0] regs_525_io_in; // @[RegFile.scala 66:20:@150422.4]
  wire  regs_525_io_reset; // @[RegFile.scala 66:20:@150422.4]
  wire [63:0] regs_525_io_out; // @[RegFile.scala 66:20:@150422.4]
  wire  regs_525_io_enable; // @[RegFile.scala 66:20:@150422.4]
  wire  regs_526_clock; // @[RegFile.scala 66:20:@150436.4]
  wire  regs_526_reset; // @[RegFile.scala 66:20:@150436.4]
  wire [63:0] regs_526_io_in; // @[RegFile.scala 66:20:@150436.4]
  wire  regs_526_io_reset; // @[RegFile.scala 66:20:@150436.4]
  wire [63:0] regs_526_io_out; // @[RegFile.scala 66:20:@150436.4]
  wire  regs_526_io_enable; // @[RegFile.scala 66:20:@150436.4]
  wire  regs_527_clock; // @[RegFile.scala 66:20:@150450.4]
  wire  regs_527_reset; // @[RegFile.scala 66:20:@150450.4]
  wire [63:0] regs_527_io_in; // @[RegFile.scala 66:20:@150450.4]
  wire  regs_527_io_reset; // @[RegFile.scala 66:20:@150450.4]
  wire [63:0] regs_527_io_out; // @[RegFile.scala 66:20:@150450.4]
  wire  regs_527_io_enable; // @[RegFile.scala 66:20:@150450.4]
  wire  regs_528_clock; // @[RegFile.scala 66:20:@150464.4]
  wire  regs_528_reset; // @[RegFile.scala 66:20:@150464.4]
  wire [63:0] regs_528_io_in; // @[RegFile.scala 66:20:@150464.4]
  wire  regs_528_io_reset; // @[RegFile.scala 66:20:@150464.4]
  wire [63:0] regs_528_io_out; // @[RegFile.scala 66:20:@150464.4]
  wire  regs_528_io_enable; // @[RegFile.scala 66:20:@150464.4]
  wire  regs_529_clock; // @[RegFile.scala 66:20:@150478.4]
  wire  regs_529_reset; // @[RegFile.scala 66:20:@150478.4]
  wire [63:0] regs_529_io_in; // @[RegFile.scala 66:20:@150478.4]
  wire  regs_529_io_reset; // @[RegFile.scala 66:20:@150478.4]
  wire [63:0] regs_529_io_out; // @[RegFile.scala 66:20:@150478.4]
  wire  regs_529_io_enable; // @[RegFile.scala 66:20:@150478.4]
  wire  regs_530_clock; // @[RegFile.scala 66:20:@150492.4]
  wire  regs_530_reset; // @[RegFile.scala 66:20:@150492.4]
  wire [63:0] regs_530_io_in; // @[RegFile.scala 66:20:@150492.4]
  wire  regs_530_io_reset; // @[RegFile.scala 66:20:@150492.4]
  wire [63:0] regs_530_io_out; // @[RegFile.scala 66:20:@150492.4]
  wire  regs_530_io_enable; // @[RegFile.scala 66:20:@150492.4]
  wire  regs_531_clock; // @[RegFile.scala 66:20:@150506.4]
  wire  regs_531_reset; // @[RegFile.scala 66:20:@150506.4]
  wire [63:0] regs_531_io_in; // @[RegFile.scala 66:20:@150506.4]
  wire  regs_531_io_reset; // @[RegFile.scala 66:20:@150506.4]
  wire [63:0] regs_531_io_out; // @[RegFile.scala 66:20:@150506.4]
  wire  regs_531_io_enable; // @[RegFile.scala 66:20:@150506.4]
  wire  regs_532_clock; // @[RegFile.scala 66:20:@150520.4]
  wire  regs_532_reset; // @[RegFile.scala 66:20:@150520.4]
  wire [63:0] regs_532_io_in; // @[RegFile.scala 66:20:@150520.4]
  wire  regs_532_io_reset; // @[RegFile.scala 66:20:@150520.4]
  wire [63:0] regs_532_io_out; // @[RegFile.scala 66:20:@150520.4]
  wire  regs_532_io_enable; // @[RegFile.scala 66:20:@150520.4]
  wire  regs_533_clock; // @[RegFile.scala 66:20:@150534.4]
  wire  regs_533_reset; // @[RegFile.scala 66:20:@150534.4]
  wire [63:0] regs_533_io_in; // @[RegFile.scala 66:20:@150534.4]
  wire  regs_533_io_reset; // @[RegFile.scala 66:20:@150534.4]
  wire [63:0] regs_533_io_out; // @[RegFile.scala 66:20:@150534.4]
  wire  regs_533_io_enable; // @[RegFile.scala 66:20:@150534.4]
  wire  regs_534_clock; // @[RegFile.scala 66:20:@150548.4]
  wire  regs_534_reset; // @[RegFile.scala 66:20:@150548.4]
  wire [63:0] regs_534_io_in; // @[RegFile.scala 66:20:@150548.4]
  wire  regs_534_io_reset; // @[RegFile.scala 66:20:@150548.4]
  wire [63:0] regs_534_io_out; // @[RegFile.scala 66:20:@150548.4]
  wire  regs_534_io_enable; // @[RegFile.scala 66:20:@150548.4]
  wire  regs_535_clock; // @[RegFile.scala 66:20:@150562.4]
  wire  regs_535_reset; // @[RegFile.scala 66:20:@150562.4]
  wire [63:0] regs_535_io_in; // @[RegFile.scala 66:20:@150562.4]
  wire  regs_535_io_reset; // @[RegFile.scala 66:20:@150562.4]
  wire [63:0] regs_535_io_out; // @[RegFile.scala 66:20:@150562.4]
  wire  regs_535_io_enable; // @[RegFile.scala 66:20:@150562.4]
  wire  regs_536_clock; // @[RegFile.scala 66:20:@150576.4]
  wire  regs_536_reset; // @[RegFile.scala 66:20:@150576.4]
  wire [63:0] regs_536_io_in; // @[RegFile.scala 66:20:@150576.4]
  wire  regs_536_io_reset; // @[RegFile.scala 66:20:@150576.4]
  wire [63:0] regs_536_io_out; // @[RegFile.scala 66:20:@150576.4]
  wire  regs_536_io_enable; // @[RegFile.scala 66:20:@150576.4]
  wire  regs_537_clock; // @[RegFile.scala 66:20:@150590.4]
  wire  regs_537_reset; // @[RegFile.scala 66:20:@150590.4]
  wire [63:0] regs_537_io_in; // @[RegFile.scala 66:20:@150590.4]
  wire  regs_537_io_reset; // @[RegFile.scala 66:20:@150590.4]
  wire [63:0] regs_537_io_out; // @[RegFile.scala 66:20:@150590.4]
  wire  regs_537_io_enable; // @[RegFile.scala 66:20:@150590.4]
  wire  regs_538_clock; // @[RegFile.scala 66:20:@150604.4]
  wire  regs_538_reset; // @[RegFile.scala 66:20:@150604.4]
  wire [63:0] regs_538_io_in; // @[RegFile.scala 66:20:@150604.4]
  wire  regs_538_io_reset; // @[RegFile.scala 66:20:@150604.4]
  wire [63:0] regs_538_io_out; // @[RegFile.scala 66:20:@150604.4]
  wire  regs_538_io_enable; // @[RegFile.scala 66:20:@150604.4]
  wire  regs_539_clock; // @[RegFile.scala 66:20:@150618.4]
  wire  regs_539_reset; // @[RegFile.scala 66:20:@150618.4]
  wire [63:0] regs_539_io_in; // @[RegFile.scala 66:20:@150618.4]
  wire  regs_539_io_reset; // @[RegFile.scala 66:20:@150618.4]
  wire [63:0] regs_539_io_out; // @[RegFile.scala 66:20:@150618.4]
  wire  regs_539_io_enable; // @[RegFile.scala 66:20:@150618.4]
  wire  regs_540_clock; // @[RegFile.scala 66:20:@150632.4]
  wire  regs_540_reset; // @[RegFile.scala 66:20:@150632.4]
  wire [63:0] regs_540_io_in; // @[RegFile.scala 66:20:@150632.4]
  wire  regs_540_io_reset; // @[RegFile.scala 66:20:@150632.4]
  wire [63:0] regs_540_io_out; // @[RegFile.scala 66:20:@150632.4]
  wire  regs_540_io_enable; // @[RegFile.scala 66:20:@150632.4]
  wire  regs_541_clock; // @[RegFile.scala 66:20:@150646.4]
  wire  regs_541_reset; // @[RegFile.scala 66:20:@150646.4]
  wire [63:0] regs_541_io_in; // @[RegFile.scala 66:20:@150646.4]
  wire  regs_541_io_reset; // @[RegFile.scala 66:20:@150646.4]
  wire [63:0] regs_541_io_out; // @[RegFile.scala 66:20:@150646.4]
  wire  regs_541_io_enable; // @[RegFile.scala 66:20:@150646.4]
  wire  regs_542_clock; // @[RegFile.scala 66:20:@150660.4]
  wire  regs_542_reset; // @[RegFile.scala 66:20:@150660.4]
  wire [63:0] regs_542_io_in; // @[RegFile.scala 66:20:@150660.4]
  wire  regs_542_io_reset; // @[RegFile.scala 66:20:@150660.4]
  wire [63:0] regs_542_io_out; // @[RegFile.scala 66:20:@150660.4]
  wire  regs_542_io_enable; // @[RegFile.scala 66:20:@150660.4]
  wire  regs_543_clock; // @[RegFile.scala 66:20:@150674.4]
  wire  regs_543_reset; // @[RegFile.scala 66:20:@150674.4]
  wire [63:0] regs_543_io_in; // @[RegFile.scala 66:20:@150674.4]
  wire  regs_543_io_reset; // @[RegFile.scala 66:20:@150674.4]
  wire [63:0] regs_543_io_out; // @[RegFile.scala 66:20:@150674.4]
  wire  regs_543_io_enable; // @[RegFile.scala 66:20:@150674.4]
  wire  regs_544_clock; // @[RegFile.scala 66:20:@150688.4]
  wire  regs_544_reset; // @[RegFile.scala 66:20:@150688.4]
  wire [63:0] regs_544_io_in; // @[RegFile.scala 66:20:@150688.4]
  wire  regs_544_io_reset; // @[RegFile.scala 66:20:@150688.4]
  wire [63:0] regs_544_io_out; // @[RegFile.scala 66:20:@150688.4]
  wire  regs_544_io_enable; // @[RegFile.scala 66:20:@150688.4]
  wire  regs_545_clock; // @[RegFile.scala 66:20:@150702.4]
  wire  regs_545_reset; // @[RegFile.scala 66:20:@150702.4]
  wire [63:0] regs_545_io_in; // @[RegFile.scala 66:20:@150702.4]
  wire  regs_545_io_reset; // @[RegFile.scala 66:20:@150702.4]
  wire [63:0] regs_545_io_out; // @[RegFile.scala 66:20:@150702.4]
  wire  regs_545_io_enable; // @[RegFile.scala 66:20:@150702.4]
  wire  regs_546_clock; // @[RegFile.scala 66:20:@150716.4]
  wire  regs_546_reset; // @[RegFile.scala 66:20:@150716.4]
  wire [63:0] regs_546_io_in; // @[RegFile.scala 66:20:@150716.4]
  wire  regs_546_io_reset; // @[RegFile.scala 66:20:@150716.4]
  wire [63:0] regs_546_io_out; // @[RegFile.scala 66:20:@150716.4]
  wire  regs_546_io_enable; // @[RegFile.scala 66:20:@150716.4]
  wire  regs_547_clock; // @[RegFile.scala 66:20:@150730.4]
  wire  regs_547_reset; // @[RegFile.scala 66:20:@150730.4]
  wire [63:0] regs_547_io_in; // @[RegFile.scala 66:20:@150730.4]
  wire  regs_547_io_reset; // @[RegFile.scala 66:20:@150730.4]
  wire [63:0] regs_547_io_out; // @[RegFile.scala 66:20:@150730.4]
  wire  regs_547_io_enable; // @[RegFile.scala 66:20:@150730.4]
  wire  regs_548_clock; // @[RegFile.scala 66:20:@150744.4]
  wire  regs_548_reset; // @[RegFile.scala 66:20:@150744.4]
  wire [63:0] regs_548_io_in; // @[RegFile.scala 66:20:@150744.4]
  wire  regs_548_io_reset; // @[RegFile.scala 66:20:@150744.4]
  wire [63:0] regs_548_io_out; // @[RegFile.scala 66:20:@150744.4]
  wire  regs_548_io_enable; // @[RegFile.scala 66:20:@150744.4]
  wire  regs_549_clock; // @[RegFile.scala 66:20:@150758.4]
  wire  regs_549_reset; // @[RegFile.scala 66:20:@150758.4]
  wire [63:0] regs_549_io_in; // @[RegFile.scala 66:20:@150758.4]
  wire  regs_549_io_reset; // @[RegFile.scala 66:20:@150758.4]
  wire [63:0] regs_549_io_out; // @[RegFile.scala 66:20:@150758.4]
  wire  regs_549_io_enable; // @[RegFile.scala 66:20:@150758.4]
  wire  regs_550_clock; // @[RegFile.scala 66:20:@150772.4]
  wire  regs_550_reset; // @[RegFile.scala 66:20:@150772.4]
  wire [63:0] regs_550_io_in; // @[RegFile.scala 66:20:@150772.4]
  wire  regs_550_io_reset; // @[RegFile.scala 66:20:@150772.4]
  wire [63:0] regs_550_io_out; // @[RegFile.scala 66:20:@150772.4]
  wire  regs_550_io_enable; // @[RegFile.scala 66:20:@150772.4]
  wire  regs_551_clock; // @[RegFile.scala 66:20:@150786.4]
  wire  regs_551_reset; // @[RegFile.scala 66:20:@150786.4]
  wire [63:0] regs_551_io_in; // @[RegFile.scala 66:20:@150786.4]
  wire  regs_551_io_reset; // @[RegFile.scala 66:20:@150786.4]
  wire [63:0] regs_551_io_out; // @[RegFile.scala 66:20:@150786.4]
  wire  regs_551_io_enable; // @[RegFile.scala 66:20:@150786.4]
  wire  regs_552_clock; // @[RegFile.scala 66:20:@150800.4]
  wire  regs_552_reset; // @[RegFile.scala 66:20:@150800.4]
  wire [63:0] regs_552_io_in; // @[RegFile.scala 66:20:@150800.4]
  wire  regs_552_io_reset; // @[RegFile.scala 66:20:@150800.4]
  wire [63:0] regs_552_io_out; // @[RegFile.scala 66:20:@150800.4]
  wire  regs_552_io_enable; // @[RegFile.scala 66:20:@150800.4]
  wire  regs_553_clock; // @[RegFile.scala 66:20:@150814.4]
  wire  regs_553_reset; // @[RegFile.scala 66:20:@150814.4]
  wire [63:0] regs_553_io_in; // @[RegFile.scala 66:20:@150814.4]
  wire  regs_553_io_reset; // @[RegFile.scala 66:20:@150814.4]
  wire [63:0] regs_553_io_out; // @[RegFile.scala 66:20:@150814.4]
  wire  regs_553_io_enable; // @[RegFile.scala 66:20:@150814.4]
  wire  regs_554_clock; // @[RegFile.scala 66:20:@150828.4]
  wire  regs_554_reset; // @[RegFile.scala 66:20:@150828.4]
  wire [63:0] regs_554_io_in; // @[RegFile.scala 66:20:@150828.4]
  wire  regs_554_io_reset; // @[RegFile.scala 66:20:@150828.4]
  wire [63:0] regs_554_io_out; // @[RegFile.scala 66:20:@150828.4]
  wire  regs_554_io_enable; // @[RegFile.scala 66:20:@150828.4]
  wire  regs_555_clock; // @[RegFile.scala 66:20:@150842.4]
  wire  regs_555_reset; // @[RegFile.scala 66:20:@150842.4]
  wire [63:0] regs_555_io_in; // @[RegFile.scala 66:20:@150842.4]
  wire  regs_555_io_reset; // @[RegFile.scala 66:20:@150842.4]
  wire [63:0] regs_555_io_out; // @[RegFile.scala 66:20:@150842.4]
  wire  regs_555_io_enable; // @[RegFile.scala 66:20:@150842.4]
  wire  regs_556_clock; // @[RegFile.scala 66:20:@150856.4]
  wire  regs_556_reset; // @[RegFile.scala 66:20:@150856.4]
  wire [63:0] regs_556_io_in; // @[RegFile.scala 66:20:@150856.4]
  wire  regs_556_io_reset; // @[RegFile.scala 66:20:@150856.4]
  wire [63:0] regs_556_io_out; // @[RegFile.scala 66:20:@150856.4]
  wire  regs_556_io_enable; // @[RegFile.scala 66:20:@150856.4]
  wire  regs_557_clock; // @[RegFile.scala 66:20:@150870.4]
  wire  regs_557_reset; // @[RegFile.scala 66:20:@150870.4]
  wire [63:0] regs_557_io_in; // @[RegFile.scala 66:20:@150870.4]
  wire  regs_557_io_reset; // @[RegFile.scala 66:20:@150870.4]
  wire [63:0] regs_557_io_out; // @[RegFile.scala 66:20:@150870.4]
  wire  regs_557_io_enable; // @[RegFile.scala 66:20:@150870.4]
  wire  regs_558_clock; // @[RegFile.scala 66:20:@150884.4]
  wire  regs_558_reset; // @[RegFile.scala 66:20:@150884.4]
  wire [63:0] regs_558_io_in; // @[RegFile.scala 66:20:@150884.4]
  wire  regs_558_io_reset; // @[RegFile.scala 66:20:@150884.4]
  wire [63:0] regs_558_io_out; // @[RegFile.scala 66:20:@150884.4]
  wire  regs_558_io_enable; // @[RegFile.scala 66:20:@150884.4]
  wire  regs_559_clock; // @[RegFile.scala 66:20:@150898.4]
  wire  regs_559_reset; // @[RegFile.scala 66:20:@150898.4]
  wire [63:0] regs_559_io_in; // @[RegFile.scala 66:20:@150898.4]
  wire  regs_559_io_reset; // @[RegFile.scala 66:20:@150898.4]
  wire [63:0] regs_559_io_out; // @[RegFile.scala 66:20:@150898.4]
  wire  regs_559_io_enable; // @[RegFile.scala 66:20:@150898.4]
  wire  regs_560_clock; // @[RegFile.scala 66:20:@150912.4]
  wire  regs_560_reset; // @[RegFile.scala 66:20:@150912.4]
  wire [63:0] regs_560_io_in; // @[RegFile.scala 66:20:@150912.4]
  wire  regs_560_io_reset; // @[RegFile.scala 66:20:@150912.4]
  wire [63:0] regs_560_io_out; // @[RegFile.scala 66:20:@150912.4]
  wire  regs_560_io_enable; // @[RegFile.scala 66:20:@150912.4]
  wire  regs_561_clock; // @[RegFile.scala 66:20:@150926.4]
  wire  regs_561_reset; // @[RegFile.scala 66:20:@150926.4]
  wire [63:0] regs_561_io_in; // @[RegFile.scala 66:20:@150926.4]
  wire  regs_561_io_reset; // @[RegFile.scala 66:20:@150926.4]
  wire [63:0] regs_561_io_out; // @[RegFile.scala 66:20:@150926.4]
  wire  regs_561_io_enable; // @[RegFile.scala 66:20:@150926.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_503; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_504; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_505; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_506; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_507; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_508; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_509; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_510; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_511; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_512; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_513; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_514; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_515; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_516; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_517; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_518; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_519; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_520; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_521; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_522; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_523; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_524; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_525; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_526; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_527; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_528; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_529; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_530; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_531; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_532; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_533; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_534; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_535; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_536; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_537; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_538; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_539; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_540; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_541; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_542; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_543; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_544; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_545; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_546; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_547; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_548; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_549; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_550; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_551; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_552; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_553; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_554; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_555; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_556; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_557; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_558; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_559; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_560; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_ins_561; // @[RegFile.scala 95:21:@150940.4]
  wire [9:0] rport_io_sel; // @[RegFile.scala 95:21:@150940.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@150940.4]
  wire  _T_3432; // @[RegFile.scala 80:42:@143076.4]
  wire  _T_3438; // @[RegFile.scala 68:46:@143088.4]
  wire  _T_3439; // @[RegFile.scala 68:34:@143089.4]
  wire  _T_3452; // @[RegFile.scala 80:42:@143107.4]
  wire  _T_3458; // @[RegFile.scala 80:42:@143119.4]
  wire  _T_3464; // @[RegFile.scala 74:80:@143131.4]
  wire  _T_3465; // @[RegFile.scala 74:68:@143132.4]
  wire  _T_3471; // @[RegFile.scala 74:80:@143145.4]
  wire  _T_3472; // @[RegFile.scala 74:68:@143146.4]
  wire  _T_3478; // @[RegFile.scala 74:80:@143159.4]
  wire  _T_3479; // @[RegFile.scala 74:68:@143160.4]
  wire  _T_3485; // @[RegFile.scala 74:80:@143173.4]
  wire  _T_3486; // @[RegFile.scala 74:68:@143174.4]
  wire  _T_3492; // @[RegFile.scala 74:80:@143187.4]
  wire  _T_3493; // @[RegFile.scala 74:68:@143188.4]
  wire  _T_3499; // @[RegFile.scala 74:80:@143201.4]
  wire  _T_3500; // @[RegFile.scala 74:68:@143202.4]
  wire  _T_3506; // @[RegFile.scala 74:80:@143215.4]
  wire  _T_3507; // @[RegFile.scala 74:68:@143216.4]
  wire  _T_3513; // @[RegFile.scala 74:80:@143229.4]
  wire  _T_3514; // @[RegFile.scala 74:68:@143230.4]
  wire  _T_3520; // @[RegFile.scala 74:80:@143243.4]
  wire  _T_3521; // @[RegFile.scala 74:68:@143244.4]
  wire  _T_3527; // @[RegFile.scala 74:80:@143257.4]
  wire  _T_3528; // @[RegFile.scala 74:68:@143258.4]
  wire  _T_3534; // @[RegFile.scala 74:80:@143271.4]
  wire  _T_3535; // @[RegFile.scala 74:68:@143272.4]
  wire  _T_3541; // @[RegFile.scala 74:80:@143285.4]
  wire  _T_3542; // @[RegFile.scala 74:68:@143286.4]
  wire  _T_3548; // @[RegFile.scala 74:80:@143299.4]
  wire  _T_3549; // @[RegFile.scala 74:68:@143300.4]
  wire  _T_3555; // @[RegFile.scala 74:80:@143313.4]
  wire  _T_3556; // @[RegFile.scala 74:68:@143314.4]
  wire  _T_3562; // @[RegFile.scala 74:80:@143327.4]
  wire  _T_3563; // @[RegFile.scala 74:68:@143328.4]
  wire  _T_3569; // @[RegFile.scala 74:80:@143341.4]
  wire  _T_3570; // @[RegFile.scala 74:68:@143342.4]
  wire  _T_3576; // @[RegFile.scala 74:80:@143355.4]
  wire  _T_3577; // @[RegFile.scala 74:68:@143356.4]
  wire  _T_3583; // @[RegFile.scala 74:80:@143369.4]
  wire  _T_3584; // @[RegFile.scala 74:68:@143370.4]
  wire  _T_3590; // @[RegFile.scala 74:80:@143383.4]
  wire  _T_3591; // @[RegFile.scala 74:68:@143384.4]
  wire  _T_3597; // @[RegFile.scala 74:80:@143397.4]
  wire  _T_3598; // @[RegFile.scala 74:68:@143398.4]
  wire  _T_3604; // @[RegFile.scala 74:80:@143411.4]
  wire  _T_3605; // @[RegFile.scala 74:68:@143412.4]
  wire  _T_3611; // @[RegFile.scala 74:80:@143425.4]
  wire  _T_3612; // @[RegFile.scala 74:68:@143426.4]
  wire  _T_3618; // @[RegFile.scala 74:80:@143439.4]
  wire  _T_3619; // @[RegFile.scala 74:68:@143440.4]
  wire  _T_3625; // @[RegFile.scala 74:80:@143453.4]
  wire  _T_3626; // @[RegFile.scala 74:68:@143454.4]
  wire  _T_3632; // @[RegFile.scala 74:80:@143467.4]
  wire  _T_3633; // @[RegFile.scala 74:68:@143468.4]
  wire  _T_3639; // @[RegFile.scala 74:80:@143481.4]
  wire  _T_3640; // @[RegFile.scala 74:68:@143482.4]
  wire  _T_3646; // @[RegFile.scala 74:80:@143495.4]
  wire  _T_3647; // @[RegFile.scala 74:68:@143496.4]
  wire  _T_3653; // @[RegFile.scala 74:80:@143509.4]
  wire  _T_3654; // @[RegFile.scala 74:68:@143510.4]
  wire  _T_3660; // @[RegFile.scala 74:80:@143523.4]
  wire  _T_3661; // @[RegFile.scala 74:68:@143524.4]
  wire  _T_3667; // @[RegFile.scala 74:80:@143537.4]
  wire  _T_3668; // @[RegFile.scala 74:68:@143538.4]
  wire  _T_3674; // @[RegFile.scala 74:80:@143551.4]
  wire  _T_3675; // @[RegFile.scala 74:68:@143552.4]
  wire  _T_3681; // @[RegFile.scala 74:80:@143565.4]
  wire  _T_3682; // @[RegFile.scala 74:68:@143566.4]
  wire  _T_3688; // @[RegFile.scala 74:80:@143579.4]
  wire  _T_3689; // @[RegFile.scala 74:68:@143580.4]
  wire  _T_3695; // @[RegFile.scala 74:80:@143593.4]
  wire  _T_3696; // @[RegFile.scala 74:68:@143594.4]
  wire  _T_3702; // @[RegFile.scala 74:80:@143607.4]
  wire  _T_3703; // @[RegFile.scala 74:68:@143608.4]
  wire  _T_3709; // @[RegFile.scala 74:80:@143621.4]
  wire  _T_3710; // @[RegFile.scala 74:68:@143622.4]
  wire  _T_3716; // @[RegFile.scala 74:80:@143635.4]
  wire  _T_3717; // @[RegFile.scala 74:68:@143636.4]
  wire  _T_3723; // @[RegFile.scala 74:80:@143649.4]
  wire  _T_3724; // @[RegFile.scala 74:68:@143650.4]
  wire  _T_3730; // @[RegFile.scala 74:80:@143663.4]
  wire  _T_3731; // @[RegFile.scala 74:68:@143664.4]
  wire  _T_3737; // @[RegFile.scala 74:80:@143677.4]
  wire  _T_3738; // @[RegFile.scala 74:68:@143678.4]
  wire  _T_3744; // @[RegFile.scala 74:80:@143691.4]
  wire  _T_3745; // @[RegFile.scala 74:68:@143692.4]
  wire  _T_3751; // @[RegFile.scala 74:80:@143705.4]
  wire  _T_3752; // @[RegFile.scala 74:68:@143706.4]
  wire  _T_3758; // @[RegFile.scala 74:80:@143719.4]
  wire  _T_3759; // @[RegFile.scala 74:68:@143720.4]
  wire  _T_3765; // @[RegFile.scala 74:80:@143733.4]
  wire  _T_3766; // @[RegFile.scala 74:68:@143734.4]
  wire  _T_3772; // @[RegFile.scala 74:80:@143747.4]
  wire  _T_3773; // @[RegFile.scala 74:68:@143748.4]
  wire  _T_3779; // @[RegFile.scala 74:80:@143761.4]
  wire  _T_3780; // @[RegFile.scala 74:68:@143762.4]
  wire  _T_3786; // @[RegFile.scala 74:80:@143775.4]
  wire  _T_3787; // @[RegFile.scala 74:68:@143776.4]
  wire  _T_3793; // @[RegFile.scala 74:80:@143789.4]
  wire  _T_3794; // @[RegFile.scala 74:68:@143790.4]
  wire  _T_3800; // @[RegFile.scala 74:80:@143803.4]
  wire  _T_3801; // @[RegFile.scala 74:68:@143804.4]
  wire  _T_3807; // @[RegFile.scala 74:80:@143817.4]
  wire  _T_3808; // @[RegFile.scala 74:68:@143818.4]
  wire  _T_3814; // @[RegFile.scala 74:80:@143831.4]
  wire  _T_3815; // @[RegFile.scala 74:68:@143832.4]
  wire  _T_3821; // @[RegFile.scala 74:80:@143845.4]
  wire  _T_3822; // @[RegFile.scala 74:68:@143846.4]
  wire  _T_3828; // @[RegFile.scala 74:80:@143859.4]
  wire  _T_3829; // @[RegFile.scala 74:68:@143860.4]
  wire  _T_3835; // @[RegFile.scala 74:80:@143873.4]
  wire  _T_3836; // @[RegFile.scala 74:68:@143874.4]
  wire  _T_3842; // @[RegFile.scala 74:80:@143887.4]
  wire  _T_3843; // @[RegFile.scala 74:68:@143888.4]
  wire  _T_3849; // @[RegFile.scala 74:80:@143901.4]
  wire  _T_3850; // @[RegFile.scala 74:68:@143902.4]
  wire  _T_3856; // @[RegFile.scala 74:80:@143915.4]
  wire  _T_3857; // @[RegFile.scala 74:68:@143916.4]
  wire  _T_3863; // @[RegFile.scala 74:80:@143929.4]
  wire  _T_3864; // @[RegFile.scala 74:68:@143930.4]
  wire  _T_3870; // @[RegFile.scala 74:80:@143943.4]
  wire  _T_3871; // @[RegFile.scala 74:68:@143944.4]
  wire  _T_3877; // @[RegFile.scala 74:80:@143957.4]
  wire  _T_3878; // @[RegFile.scala 74:68:@143958.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@143073.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@143085.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@143104.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@143116.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@143128.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@143142.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@143156.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@143170.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@143184.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@143198.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@143212.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@143226.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@143240.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@143254.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@143268.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@143282.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@143296.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@143310.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@143324.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@143338.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@143352.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@143366.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@143380.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@143394.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@143408.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@143422.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@143436.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@143450.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@143464.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@143478.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@143492.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@143506.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@143520.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@143534.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@143548.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@143562.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@143576.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@143590.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@143604.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@143618.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@143632.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@143646.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@143660.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@143674.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@143688.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@143702.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@143716.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@143730.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@143744.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@143758.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@143772.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@143786.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@143800.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@143814.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@143828.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@143842.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@143856.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@143870.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@143884.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@143898.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@143912.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@143926.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@143940.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@143954.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@143968.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@143982.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@143996.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@144010.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@144024.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@144038.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@144052.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@144066.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@144080.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@144094.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@144108.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@144122.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@144136.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@144150.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@144164.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@144178.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@144192.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@144206.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@144220.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@144234.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@144248.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@144262.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@144276.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@144290.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@144304.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@144318.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@144332.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@144346.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@144360.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@144374.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@144388.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@144402.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@144416.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@144430.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@144444.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@144458.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@144472.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@144486.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@144500.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@144514.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@144528.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@144542.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@144556.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@144570.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@144584.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@144598.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@144612.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@144626.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@144640.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@144654.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@144668.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@144682.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@144696.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@144710.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@144724.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@144738.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@144752.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@144766.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@144780.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@144794.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@144808.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@144822.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@144836.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@144850.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@144864.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@144878.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@144892.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@144906.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@144920.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@144934.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@144948.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@144962.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@144976.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@144990.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@145004.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@145018.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@145032.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@145046.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@145060.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@145074.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@145088.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@145102.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@145116.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@145130.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@145144.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@145158.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@145172.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@145186.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@145200.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@145214.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@145228.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@145242.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@145256.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@145270.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@145284.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@145298.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@145312.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@145326.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@145340.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@145354.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@145368.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@145382.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@145396.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@145410.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@145424.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@145438.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@145452.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@145466.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@145480.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@145494.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@145508.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@145522.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@145536.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@145550.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@145564.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@145578.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@145592.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@145606.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@145620.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@145634.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@145648.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@145662.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@145676.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@145690.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@145704.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@145718.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@145732.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@145746.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@145760.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@145774.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@145788.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@145802.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@145816.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@145830.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@145844.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@145858.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@145872.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@145886.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@145900.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@145914.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@145928.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@145942.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@145956.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@145970.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@145984.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@145998.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@146012.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@146026.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@146040.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@146054.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@146068.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@146082.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@146096.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@146110.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@146124.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@146138.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@146152.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@146166.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@146180.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@146194.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@146208.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@146222.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@146236.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@146250.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@146264.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@146278.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@146292.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@146306.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@146320.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@146334.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@146348.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@146362.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@146376.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@146390.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@146404.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@146418.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@146432.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@146446.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@146460.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@146474.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@146488.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@146502.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@146516.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@146530.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@146544.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@146558.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@146572.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@146586.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@146600.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@146614.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@146628.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@146642.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@146656.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@146670.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@146684.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@146698.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@146712.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@146726.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@146740.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@146754.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@146768.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@146782.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@146796.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@146810.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@146824.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@146838.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@146852.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@146866.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@146880.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@146894.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@146908.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@146922.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@146936.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@146950.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@146964.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@146978.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@146992.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@147006.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@147020.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@147034.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@147048.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@147062.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@147076.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@147090.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@147104.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@147118.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@147132.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@147146.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@147160.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@147174.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@147188.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@147202.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@147216.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@147230.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@147244.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@147258.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@147272.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@147286.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@147300.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@147314.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@147328.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@147342.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@147356.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@147370.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@147384.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@147398.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@147412.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@147426.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@147440.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@147454.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@147468.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@147482.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@147496.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@147510.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@147524.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@147538.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@147552.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@147566.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@147580.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@147594.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@147608.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@147622.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@147636.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@147650.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@147664.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@147678.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@147692.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@147706.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@147720.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@147734.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@147748.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@147762.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@147776.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@147790.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@147804.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@147818.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@147832.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@147846.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@147860.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@147874.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@147888.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@147902.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@147916.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@147930.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@147944.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@147958.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@147972.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@147986.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@148000.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@148014.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@148028.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@148042.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@148056.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@148070.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@148084.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@148098.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@148112.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@148126.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@148140.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@148154.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@148168.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@148182.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@148196.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@148210.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@148224.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@148238.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@148252.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@148266.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@148280.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@148294.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@148308.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@148322.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@148336.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@148350.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@148364.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@148378.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@148392.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@148406.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@148420.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@148434.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@148448.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@148462.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@148476.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@148490.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@148504.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@148518.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@148532.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@148546.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@148560.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@148574.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@148588.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@148602.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@148616.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@148630.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@148644.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@148658.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@148672.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@148686.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@148700.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@148714.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@148728.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@148742.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@148756.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@148770.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@148784.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@148798.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@148812.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@148826.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@148840.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@148854.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@148868.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@148882.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@148896.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@148910.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@148924.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@148938.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@148952.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@148966.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@148980.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@148994.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@149008.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@149022.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@149036.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@149050.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@149064.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@149078.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@149092.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@149106.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@149120.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@149134.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@149148.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@149162.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@149176.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@149190.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@149204.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@149218.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@149232.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@149246.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@149260.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@149274.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@149288.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@149302.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@149316.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@149330.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@149344.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@149358.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@149372.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@149386.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@149400.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@149414.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@149428.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@149442.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@149456.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@149470.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@149484.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@149498.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@149512.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@149526.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@149540.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@149554.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@149568.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@149582.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@149596.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@149610.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@149624.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@149638.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@149652.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@149666.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@149680.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@149694.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@149708.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@149722.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@149736.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@149750.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@149764.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@149778.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@149792.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@149806.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@149820.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@149834.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@149848.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@149862.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@149876.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@149890.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@149904.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@149918.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@149932.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@149946.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@149960.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@149974.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@149988.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@150002.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@150016.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@150030.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@150044.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@150058.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@150072.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@150086.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@150100.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  FringeFF regs_503 ( // @[RegFile.scala 66:20:@150114.4]
    .clock(regs_503_clock),
    .reset(regs_503_reset),
    .io_in(regs_503_io_in),
    .io_reset(regs_503_io_reset),
    .io_out(regs_503_io_out),
    .io_enable(regs_503_io_enable)
  );
  FringeFF regs_504 ( // @[RegFile.scala 66:20:@150128.4]
    .clock(regs_504_clock),
    .reset(regs_504_reset),
    .io_in(regs_504_io_in),
    .io_reset(regs_504_io_reset),
    .io_out(regs_504_io_out),
    .io_enable(regs_504_io_enable)
  );
  FringeFF regs_505 ( // @[RegFile.scala 66:20:@150142.4]
    .clock(regs_505_clock),
    .reset(regs_505_reset),
    .io_in(regs_505_io_in),
    .io_reset(regs_505_io_reset),
    .io_out(regs_505_io_out),
    .io_enable(regs_505_io_enable)
  );
  FringeFF regs_506 ( // @[RegFile.scala 66:20:@150156.4]
    .clock(regs_506_clock),
    .reset(regs_506_reset),
    .io_in(regs_506_io_in),
    .io_reset(regs_506_io_reset),
    .io_out(regs_506_io_out),
    .io_enable(regs_506_io_enable)
  );
  FringeFF regs_507 ( // @[RegFile.scala 66:20:@150170.4]
    .clock(regs_507_clock),
    .reset(regs_507_reset),
    .io_in(regs_507_io_in),
    .io_reset(regs_507_io_reset),
    .io_out(regs_507_io_out),
    .io_enable(regs_507_io_enable)
  );
  FringeFF regs_508 ( // @[RegFile.scala 66:20:@150184.4]
    .clock(regs_508_clock),
    .reset(regs_508_reset),
    .io_in(regs_508_io_in),
    .io_reset(regs_508_io_reset),
    .io_out(regs_508_io_out),
    .io_enable(regs_508_io_enable)
  );
  FringeFF regs_509 ( // @[RegFile.scala 66:20:@150198.4]
    .clock(regs_509_clock),
    .reset(regs_509_reset),
    .io_in(regs_509_io_in),
    .io_reset(regs_509_io_reset),
    .io_out(regs_509_io_out),
    .io_enable(regs_509_io_enable)
  );
  FringeFF regs_510 ( // @[RegFile.scala 66:20:@150212.4]
    .clock(regs_510_clock),
    .reset(regs_510_reset),
    .io_in(regs_510_io_in),
    .io_reset(regs_510_io_reset),
    .io_out(regs_510_io_out),
    .io_enable(regs_510_io_enable)
  );
  FringeFF regs_511 ( // @[RegFile.scala 66:20:@150226.4]
    .clock(regs_511_clock),
    .reset(regs_511_reset),
    .io_in(regs_511_io_in),
    .io_reset(regs_511_io_reset),
    .io_out(regs_511_io_out),
    .io_enable(regs_511_io_enable)
  );
  FringeFF regs_512 ( // @[RegFile.scala 66:20:@150240.4]
    .clock(regs_512_clock),
    .reset(regs_512_reset),
    .io_in(regs_512_io_in),
    .io_reset(regs_512_io_reset),
    .io_out(regs_512_io_out),
    .io_enable(regs_512_io_enable)
  );
  FringeFF regs_513 ( // @[RegFile.scala 66:20:@150254.4]
    .clock(regs_513_clock),
    .reset(regs_513_reset),
    .io_in(regs_513_io_in),
    .io_reset(regs_513_io_reset),
    .io_out(regs_513_io_out),
    .io_enable(regs_513_io_enable)
  );
  FringeFF regs_514 ( // @[RegFile.scala 66:20:@150268.4]
    .clock(regs_514_clock),
    .reset(regs_514_reset),
    .io_in(regs_514_io_in),
    .io_reset(regs_514_io_reset),
    .io_out(regs_514_io_out),
    .io_enable(regs_514_io_enable)
  );
  FringeFF regs_515 ( // @[RegFile.scala 66:20:@150282.4]
    .clock(regs_515_clock),
    .reset(regs_515_reset),
    .io_in(regs_515_io_in),
    .io_reset(regs_515_io_reset),
    .io_out(regs_515_io_out),
    .io_enable(regs_515_io_enable)
  );
  FringeFF regs_516 ( // @[RegFile.scala 66:20:@150296.4]
    .clock(regs_516_clock),
    .reset(regs_516_reset),
    .io_in(regs_516_io_in),
    .io_reset(regs_516_io_reset),
    .io_out(regs_516_io_out),
    .io_enable(regs_516_io_enable)
  );
  FringeFF regs_517 ( // @[RegFile.scala 66:20:@150310.4]
    .clock(regs_517_clock),
    .reset(regs_517_reset),
    .io_in(regs_517_io_in),
    .io_reset(regs_517_io_reset),
    .io_out(regs_517_io_out),
    .io_enable(regs_517_io_enable)
  );
  FringeFF regs_518 ( // @[RegFile.scala 66:20:@150324.4]
    .clock(regs_518_clock),
    .reset(regs_518_reset),
    .io_in(regs_518_io_in),
    .io_reset(regs_518_io_reset),
    .io_out(regs_518_io_out),
    .io_enable(regs_518_io_enable)
  );
  FringeFF regs_519 ( // @[RegFile.scala 66:20:@150338.4]
    .clock(regs_519_clock),
    .reset(regs_519_reset),
    .io_in(regs_519_io_in),
    .io_reset(regs_519_io_reset),
    .io_out(regs_519_io_out),
    .io_enable(regs_519_io_enable)
  );
  FringeFF regs_520 ( // @[RegFile.scala 66:20:@150352.4]
    .clock(regs_520_clock),
    .reset(regs_520_reset),
    .io_in(regs_520_io_in),
    .io_reset(regs_520_io_reset),
    .io_out(regs_520_io_out),
    .io_enable(regs_520_io_enable)
  );
  FringeFF regs_521 ( // @[RegFile.scala 66:20:@150366.4]
    .clock(regs_521_clock),
    .reset(regs_521_reset),
    .io_in(regs_521_io_in),
    .io_reset(regs_521_io_reset),
    .io_out(regs_521_io_out),
    .io_enable(regs_521_io_enable)
  );
  FringeFF regs_522 ( // @[RegFile.scala 66:20:@150380.4]
    .clock(regs_522_clock),
    .reset(regs_522_reset),
    .io_in(regs_522_io_in),
    .io_reset(regs_522_io_reset),
    .io_out(regs_522_io_out),
    .io_enable(regs_522_io_enable)
  );
  FringeFF regs_523 ( // @[RegFile.scala 66:20:@150394.4]
    .clock(regs_523_clock),
    .reset(regs_523_reset),
    .io_in(regs_523_io_in),
    .io_reset(regs_523_io_reset),
    .io_out(regs_523_io_out),
    .io_enable(regs_523_io_enable)
  );
  FringeFF regs_524 ( // @[RegFile.scala 66:20:@150408.4]
    .clock(regs_524_clock),
    .reset(regs_524_reset),
    .io_in(regs_524_io_in),
    .io_reset(regs_524_io_reset),
    .io_out(regs_524_io_out),
    .io_enable(regs_524_io_enable)
  );
  FringeFF regs_525 ( // @[RegFile.scala 66:20:@150422.4]
    .clock(regs_525_clock),
    .reset(regs_525_reset),
    .io_in(regs_525_io_in),
    .io_reset(regs_525_io_reset),
    .io_out(regs_525_io_out),
    .io_enable(regs_525_io_enable)
  );
  FringeFF regs_526 ( // @[RegFile.scala 66:20:@150436.4]
    .clock(regs_526_clock),
    .reset(regs_526_reset),
    .io_in(regs_526_io_in),
    .io_reset(regs_526_io_reset),
    .io_out(regs_526_io_out),
    .io_enable(regs_526_io_enable)
  );
  FringeFF regs_527 ( // @[RegFile.scala 66:20:@150450.4]
    .clock(regs_527_clock),
    .reset(regs_527_reset),
    .io_in(regs_527_io_in),
    .io_reset(regs_527_io_reset),
    .io_out(regs_527_io_out),
    .io_enable(regs_527_io_enable)
  );
  FringeFF regs_528 ( // @[RegFile.scala 66:20:@150464.4]
    .clock(regs_528_clock),
    .reset(regs_528_reset),
    .io_in(regs_528_io_in),
    .io_reset(regs_528_io_reset),
    .io_out(regs_528_io_out),
    .io_enable(regs_528_io_enable)
  );
  FringeFF regs_529 ( // @[RegFile.scala 66:20:@150478.4]
    .clock(regs_529_clock),
    .reset(regs_529_reset),
    .io_in(regs_529_io_in),
    .io_reset(regs_529_io_reset),
    .io_out(regs_529_io_out),
    .io_enable(regs_529_io_enable)
  );
  FringeFF regs_530 ( // @[RegFile.scala 66:20:@150492.4]
    .clock(regs_530_clock),
    .reset(regs_530_reset),
    .io_in(regs_530_io_in),
    .io_reset(regs_530_io_reset),
    .io_out(regs_530_io_out),
    .io_enable(regs_530_io_enable)
  );
  FringeFF regs_531 ( // @[RegFile.scala 66:20:@150506.4]
    .clock(regs_531_clock),
    .reset(regs_531_reset),
    .io_in(regs_531_io_in),
    .io_reset(regs_531_io_reset),
    .io_out(regs_531_io_out),
    .io_enable(regs_531_io_enable)
  );
  FringeFF regs_532 ( // @[RegFile.scala 66:20:@150520.4]
    .clock(regs_532_clock),
    .reset(regs_532_reset),
    .io_in(regs_532_io_in),
    .io_reset(regs_532_io_reset),
    .io_out(regs_532_io_out),
    .io_enable(regs_532_io_enable)
  );
  FringeFF regs_533 ( // @[RegFile.scala 66:20:@150534.4]
    .clock(regs_533_clock),
    .reset(regs_533_reset),
    .io_in(regs_533_io_in),
    .io_reset(regs_533_io_reset),
    .io_out(regs_533_io_out),
    .io_enable(regs_533_io_enable)
  );
  FringeFF regs_534 ( // @[RegFile.scala 66:20:@150548.4]
    .clock(regs_534_clock),
    .reset(regs_534_reset),
    .io_in(regs_534_io_in),
    .io_reset(regs_534_io_reset),
    .io_out(regs_534_io_out),
    .io_enable(regs_534_io_enable)
  );
  FringeFF regs_535 ( // @[RegFile.scala 66:20:@150562.4]
    .clock(regs_535_clock),
    .reset(regs_535_reset),
    .io_in(regs_535_io_in),
    .io_reset(regs_535_io_reset),
    .io_out(regs_535_io_out),
    .io_enable(regs_535_io_enable)
  );
  FringeFF regs_536 ( // @[RegFile.scala 66:20:@150576.4]
    .clock(regs_536_clock),
    .reset(regs_536_reset),
    .io_in(regs_536_io_in),
    .io_reset(regs_536_io_reset),
    .io_out(regs_536_io_out),
    .io_enable(regs_536_io_enable)
  );
  FringeFF regs_537 ( // @[RegFile.scala 66:20:@150590.4]
    .clock(regs_537_clock),
    .reset(regs_537_reset),
    .io_in(regs_537_io_in),
    .io_reset(regs_537_io_reset),
    .io_out(regs_537_io_out),
    .io_enable(regs_537_io_enable)
  );
  FringeFF regs_538 ( // @[RegFile.scala 66:20:@150604.4]
    .clock(regs_538_clock),
    .reset(regs_538_reset),
    .io_in(regs_538_io_in),
    .io_reset(regs_538_io_reset),
    .io_out(regs_538_io_out),
    .io_enable(regs_538_io_enable)
  );
  FringeFF regs_539 ( // @[RegFile.scala 66:20:@150618.4]
    .clock(regs_539_clock),
    .reset(regs_539_reset),
    .io_in(regs_539_io_in),
    .io_reset(regs_539_io_reset),
    .io_out(regs_539_io_out),
    .io_enable(regs_539_io_enable)
  );
  FringeFF regs_540 ( // @[RegFile.scala 66:20:@150632.4]
    .clock(regs_540_clock),
    .reset(regs_540_reset),
    .io_in(regs_540_io_in),
    .io_reset(regs_540_io_reset),
    .io_out(regs_540_io_out),
    .io_enable(regs_540_io_enable)
  );
  FringeFF regs_541 ( // @[RegFile.scala 66:20:@150646.4]
    .clock(regs_541_clock),
    .reset(regs_541_reset),
    .io_in(regs_541_io_in),
    .io_reset(regs_541_io_reset),
    .io_out(regs_541_io_out),
    .io_enable(regs_541_io_enable)
  );
  FringeFF regs_542 ( // @[RegFile.scala 66:20:@150660.4]
    .clock(regs_542_clock),
    .reset(regs_542_reset),
    .io_in(regs_542_io_in),
    .io_reset(regs_542_io_reset),
    .io_out(regs_542_io_out),
    .io_enable(regs_542_io_enable)
  );
  FringeFF regs_543 ( // @[RegFile.scala 66:20:@150674.4]
    .clock(regs_543_clock),
    .reset(regs_543_reset),
    .io_in(regs_543_io_in),
    .io_reset(regs_543_io_reset),
    .io_out(regs_543_io_out),
    .io_enable(regs_543_io_enable)
  );
  FringeFF regs_544 ( // @[RegFile.scala 66:20:@150688.4]
    .clock(regs_544_clock),
    .reset(regs_544_reset),
    .io_in(regs_544_io_in),
    .io_reset(regs_544_io_reset),
    .io_out(regs_544_io_out),
    .io_enable(regs_544_io_enable)
  );
  FringeFF regs_545 ( // @[RegFile.scala 66:20:@150702.4]
    .clock(regs_545_clock),
    .reset(regs_545_reset),
    .io_in(regs_545_io_in),
    .io_reset(regs_545_io_reset),
    .io_out(regs_545_io_out),
    .io_enable(regs_545_io_enable)
  );
  FringeFF regs_546 ( // @[RegFile.scala 66:20:@150716.4]
    .clock(regs_546_clock),
    .reset(regs_546_reset),
    .io_in(regs_546_io_in),
    .io_reset(regs_546_io_reset),
    .io_out(regs_546_io_out),
    .io_enable(regs_546_io_enable)
  );
  FringeFF regs_547 ( // @[RegFile.scala 66:20:@150730.4]
    .clock(regs_547_clock),
    .reset(regs_547_reset),
    .io_in(regs_547_io_in),
    .io_reset(regs_547_io_reset),
    .io_out(regs_547_io_out),
    .io_enable(regs_547_io_enable)
  );
  FringeFF regs_548 ( // @[RegFile.scala 66:20:@150744.4]
    .clock(regs_548_clock),
    .reset(regs_548_reset),
    .io_in(regs_548_io_in),
    .io_reset(regs_548_io_reset),
    .io_out(regs_548_io_out),
    .io_enable(regs_548_io_enable)
  );
  FringeFF regs_549 ( // @[RegFile.scala 66:20:@150758.4]
    .clock(regs_549_clock),
    .reset(regs_549_reset),
    .io_in(regs_549_io_in),
    .io_reset(regs_549_io_reset),
    .io_out(regs_549_io_out),
    .io_enable(regs_549_io_enable)
  );
  FringeFF regs_550 ( // @[RegFile.scala 66:20:@150772.4]
    .clock(regs_550_clock),
    .reset(regs_550_reset),
    .io_in(regs_550_io_in),
    .io_reset(regs_550_io_reset),
    .io_out(regs_550_io_out),
    .io_enable(regs_550_io_enable)
  );
  FringeFF regs_551 ( // @[RegFile.scala 66:20:@150786.4]
    .clock(regs_551_clock),
    .reset(regs_551_reset),
    .io_in(regs_551_io_in),
    .io_reset(regs_551_io_reset),
    .io_out(regs_551_io_out),
    .io_enable(regs_551_io_enable)
  );
  FringeFF regs_552 ( // @[RegFile.scala 66:20:@150800.4]
    .clock(regs_552_clock),
    .reset(regs_552_reset),
    .io_in(regs_552_io_in),
    .io_reset(regs_552_io_reset),
    .io_out(regs_552_io_out),
    .io_enable(regs_552_io_enable)
  );
  FringeFF regs_553 ( // @[RegFile.scala 66:20:@150814.4]
    .clock(regs_553_clock),
    .reset(regs_553_reset),
    .io_in(regs_553_io_in),
    .io_reset(regs_553_io_reset),
    .io_out(regs_553_io_out),
    .io_enable(regs_553_io_enable)
  );
  FringeFF regs_554 ( // @[RegFile.scala 66:20:@150828.4]
    .clock(regs_554_clock),
    .reset(regs_554_reset),
    .io_in(regs_554_io_in),
    .io_reset(regs_554_io_reset),
    .io_out(regs_554_io_out),
    .io_enable(regs_554_io_enable)
  );
  FringeFF regs_555 ( // @[RegFile.scala 66:20:@150842.4]
    .clock(regs_555_clock),
    .reset(regs_555_reset),
    .io_in(regs_555_io_in),
    .io_reset(regs_555_io_reset),
    .io_out(regs_555_io_out),
    .io_enable(regs_555_io_enable)
  );
  FringeFF regs_556 ( // @[RegFile.scala 66:20:@150856.4]
    .clock(regs_556_clock),
    .reset(regs_556_reset),
    .io_in(regs_556_io_in),
    .io_reset(regs_556_io_reset),
    .io_out(regs_556_io_out),
    .io_enable(regs_556_io_enable)
  );
  FringeFF regs_557 ( // @[RegFile.scala 66:20:@150870.4]
    .clock(regs_557_clock),
    .reset(regs_557_reset),
    .io_in(regs_557_io_in),
    .io_reset(regs_557_io_reset),
    .io_out(regs_557_io_out),
    .io_enable(regs_557_io_enable)
  );
  FringeFF regs_558 ( // @[RegFile.scala 66:20:@150884.4]
    .clock(regs_558_clock),
    .reset(regs_558_reset),
    .io_in(regs_558_io_in),
    .io_reset(regs_558_io_reset),
    .io_out(regs_558_io_out),
    .io_enable(regs_558_io_enable)
  );
  FringeFF regs_559 ( // @[RegFile.scala 66:20:@150898.4]
    .clock(regs_559_clock),
    .reset(regs_559_reset),
    .io_in(regs_559_io_in),
    .io_reset(regs_559_io_reset),
    .io_out(regs_559_io_out),
    .io_enable(regs_559_io_enable)
  );
  FringeFF regs_560 ( // @[RegFile.scala 66:20:@150912.4]
    .clock(regs_560_clock),
    .reset(regs_560_reset),
    .io_in(regs_560_io_in),
    .io_reset(regs_560_io_reset),
    .io_out(regs_560_io_out),
    .io_enable(regs_560_io_enable)
  );
  FringeFF regs_561 ( // @[RegFile.scala 66:20:@150926.4]
    .clock(regs_561_clock),
    .reset(regs_561_reset),
    .io_in(regs_561_io_in),
    .io_reset(regs_561_io_reset),
    .io_out(regs_561_io_out),
    .io_enable(regs_561_io_enable)
  );
  MuxN_2 rport ( // @[RegFile.scala 95:21:@150940.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_ins_503(rport_io_ins_503),
    .io_ins_504(rport_io_ins_504),
    .io_ins_505(rport_io_ins_505),
    .io_ins_506(rport_io_ins_506),
    .io_ins_507(rport_io_ins_507),
    .io_ins_508(rport_io_ins_508),
    .io_ins_509(rport_io_ins_509),
    .io_ins_510(rport_io_ins_510),
    .io_ins_511(rport_io_ins_511),
    .io_ins_512(rport_io_ins_512),
    .io_ins_513(rport_io_ins_513),
    .io_ins_514(rport_io_ins_514),
    .io_ins_515(rport_io_ins_515),
    .io_ins_516(rport_io_ins_516),
    .io_ins_517(rport_io_ins_517),
    .io_ins_518(rport_io_ins_518),
    .io_ins_519(rport_io_ins_519),
    .io_ins_520(rport_io_ins_520),
    .io_ins_521(rport_io_ins_521),
    .io_ins_522(rport_io_ins_522),
    .io_ins_523(rport_io_ins_523),
    .io_ins_524(rport_io_ins_524),
    .io_ins_525(rport_io_ins_525),
    .io_ins_526(rport_io_ins_526),
    .io_ins_527(rport_io_ins_527),
    .io_ins_528(rport_io_ins_528),
    .io_ins_529(rport_io_ins_529),
    .io_ins_530(rport_io_ins_530),
    .io_ins_531(rport_io_ins_531),
    .io_ins_532(rport_io_ins_532),
    .io_ins_533(rport_io_ins_533),
    .io_ins_534(rport_io_ins_534),
    .io_ins_535(rport_io_ins_535),
    .io_ins_536(rport_io_ins_536),
    .io_ins_537(rport_io_ins_537),
    .io_ins_538(rport_io_ins_538),
    .io_ins_539(rport_io_ins_539),
    .io_ins_540(rport_io_ins_540),
    .io_ins_541(rport_io_ins_541),
    .io_ins_542(rport_io_ins_542),
    .io_ins_543(rport_io_ins_543),
    .io_ins_544(rport_io_ins_544),
    .io_ins_545(rport_io_ins_545),
    .io_ins_546(rport_io_ins_546),
    .io_ins_547(rport_io_ins_547),
    .io_ins_548(rport_io_ins_548),
    .io_ins_549(rport_io_ins_549),
    .io_ins_550(rport_io_ins_550),
    .io_ins_551(rport_io_ins_551),
    .io_ins_552(rport_io_ins_552),
    .io_ins_553(rport_io_ins_553),
    .io_ins_554(rport_io_ins_554),
    .io_ins_555(rport_io_ins_555),
    .io_ins_556(rport_io_ins_556),
    .io_ins_557(rport_io_ins_557),
    .io_ins_558(rport_io_ins_558),
    .io_ins_559(rport_io_ins_559),
    .io_ins_560(rport_io_ins_560),
    .io_ins_561(rport_io_ins_561),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3432 = io_waddr == 11'h0; // @[RegFile.scala 80:42:@143076.4]
  assign _T_3438 = io_waddr == 11'h1; // @[RegFile.scala 68:46:@143088.4]
  assign _T_3439 = io_wen & _T_3438; // @[RegFile.scala 68:34:@143089.4]
  assign _T_3452 = io_waddr == 11'h2; // @[RegFile.scala 80:42:@143107.4]
  assign _T_3458 = io_waddr == 11'h3; // @[RegFile.scala 80:42:@143119.4]
  assign _T_3464 = io_waddr == 11'h4; // @[RegFile.scala 74:80:@143131.4]
  assign _T_3465 = io_wen & _T_3464; // @[RegFile.scala 74:68:@143132.4]
  assign _T_3471 = io_waddr == 11'h5; // @[RegFile.scala 74:80:@143145.4]
  assign _T_3472 = io_wen & _T_3471; // @[RegFile.scala 74:68:@143146.4]
  assign _T_3478 = io_waddr == 11'h6; // @[RegFile.scala 74:80:@143159.4]
  assign _T_3479 = io_wen & _T_3478; // @[RegFile.scala 74:68:@143160.4]
  assign _T_3485 = io_waddr == 11'h7; // @[RegFile.scala 74:80:@143173.4]
  assign _T_3486 = io_wen & _T_3485; // @[RegFile.scala 74:68:@143174.4]
  assign _T_3492 = io_waddr == 11'h8; // @[RegFile.scala 74:80:@143187.4]
  assign _T_3493 = io_wen & _T_3492; // @[RegFile.scala 74:68:@143188.4]
  assign _T_3499 = io_waddr == 11'h9; // @[RegFile.scala 74:80:@143201.4]
  assign _T_3500 = io_wen & _T_3499; // @[RegFile.scala 74:68:@143202.4]
  assign _T_3506 = io_waddr == 11'ha; // @[RegFile.scala 74:80:@143215.4]
  assign _T_3507 = io_wen & _T_3506; // @[RegFile.scala 74:68:@143216.4]
  assign _T_3513 = io_waddr == 11'hb; // @[RegFile.scala 74:80:@143229.4]
  assign _T_3514 = io_wen & _T_3513; // @[RegFile.scala 74:68:@143230.4]
  assign _T_3520 = io_waddr == 11'hc; // @[RegFile.scala 74:80:@143243.4]
  assign _T_3521 = io_wen & _T_3520; // @[RegFile.scala 74:68:@143244.4]
  assign _T_3527 = io_waddr == 11'hd; // @[RegFile.scala 74:80:@143257.4]
  assign _T_3528 = io_wen & _T_3527; // @[RegFile.scala 74:68:@143258.4]
  assign _T_3534 = io_waddr == 11'he; // @[RegFile.scala 74:80:@143271.4]
  assign _T_3535 = io_wen & _T_3534; // @[RegFile.scala 74:68:@143272.4]
  assign _T_3541 = io_waddr == 11'hf; // @[RegFile.scala 74:80:@143285.4]
  assign _T_3542 = io_wen & _T_3541; // @[RegFile.scala 74:68:@143286.4]
  assign _T_3548 = io_waddr == 11'h10; // @[RegFile.scala 74:80:@143299.4]
  assign _T_3549 = io_wen & _T_3548; // @[RegFile.scala 74:68:@143300.4]
  assign _T_3555 = io_waddr == 11'h11; // @[RegFile.scala 74:80:@143313.4]
  assign _T_3556 = io_wen & _T_3555; // @[RegFile.scala 74:68:@143314.4]
  assign _T_3562 = io_waddr == 11'h12; // @[RegFile.scala 74:80:@143327.4]
  assign _T_3563 = io_wen & _T_3562; // @[RegFile.scala 74:68:@143328.4]
  assign _T_3569 = io_waddr == 11'h13; // @[RegFile.scala 74:80:@143341.4]
  assign _T_3570 = io_wen & _T_3569; // @[RegFile.scala 74:68:@143342.4]
  assign _T_3576 = io_waddr == 11'h14; // @[RegFile.scala 74:80:@143355.4]
  assign _T_3577 = io_wen & _T_3576; // @[RegFile.scala 74:68:@143356.4]
  assign _T_3583 = io_waddr == 11'h15; // @[RegFile.scala 74:80:@143369.4]
  assign _T_3584 = io_wen & _T_3583; // @[RegFile.scala 74:68:@143370.4]
  assign _T_3590 = io_waddr == 11'h16; // @[RegFile.scala 74:80:@143383.4]
  assign _T_3591 = io_wen & _T_3590; // @[RegFile.scala 74:68:@143384.4]
  assign _T_3597 = io_waddr == 11'h17; // @[RegFile.scala 74:80:@143397.4]
  assign _T_3598 = io_wen & _T_3597; // @[RegFile.scala 74:68:@143398.4]
  assign _T_3604 = io_waddr == 11'h18; // @[RegFile.scala 74:80:@143411.4]
  assign _T_3605 = io_wen & _T_3604; // @[RegFile.scala 74:68:@143412.4]
  assign _T_3611 = io_waddr == 11'h19; // @[RegFile.scala 74:80:@143425.4]
  assign _T_3612 = io_wen & _T_3611; // @[RegFile.scala 74:68:@143426.4]
  assign _T_3618 = io_waddr == 11'h1a; // @[RegFile.scala 74:80:@143439.4]
  assign _T_3619 = io_wen & _T_3618; // @[RegFile.scala 74:68:@143440.4]
  assign _T_3625 = io_waddr == 11'h1b; // @[RegFile.scala 74:80:@143453.4]
  assign _T_3626 = io_wen & _T_3625; // @[RegFile.scala 74:68:@143454.4]
  assign _T_3632 = io_waddr == 11'h1c; // @[RegFile.scala 74:80:@143467.4]
  assign _T_3633 = io_wen & _T_3632; // @[RegFile.scala 74:68:@143468.4]
  assign _T_3639 = io_waddr == 11'h1d; // @[RegFile.scala 74:80:@143481.4]
  assign _T_3640 = io_wen & _T_3639; // @[RegFile.scala 74:68:@143482.4]
  assign _T_3646 = io_waddr == 11'h1e; // @[RegFile.scala 74:80:@143495.4]
  assign _T_3647 = io_wen & _T_3646; // @[RegFile.scala 74:68:@143496.4]
  assign _T_3653 = io_waddr == 11'h1f; // @[RegFile.scala 74:80:@143509.4]
  assign _T_3654 = io_wen & _T_3653; // @[RegFile.scala 74:68:@143510.4]
  assign _T_3660 = io_waddr == 11'h20; // @[RegFile.scala 74:80:@143523.4]
  assign _T_3661 = io_wen & _T_3660; // @[RegFile.scala 74:68:@143524.4]
  assign _T_3667 = io_waddr == 11'h21; // @[RegFile.scala 74:80:@143537.4]
  assign _T_3668 = io_wen & _T_3667; // @[RegFile.scala 74:68:@143538.4]
  assign _T_3674 = io_waddr == 11'h22; // @[RegFile.scala 74:80:@143551.4]
  assign _T_3675 = io_wen & _T_3674; // @[RegFile.scala 74:68:@143552.4]
  assign _T_3681 = io_waddr == 11'h23; // @[RegFile.scala 74:80:@143565.4]
  assign _T_3682 = io_wen & _T_3681; // @[RegFile.scala 74:68:@143566.4]
  assign _T_3688 = io_waddr == 11'h24; // @[RegFile.scala 74:80:@143579.4]
  assign _T_3689 = io_wen & _T_3688; // @[RegFile.scala 74:68:@143580.4]
  assign _T_3695 = io_waddr == 11'h25; // @[RegFile.scala 74:80:@143593.4]
  assign _T_3696 = io_wen & _T_3695; // @[RegFile.scala 74:68:@143594.4]
  assign _T_3702 = io_waddr == 11'h26; // @[RegFile.scala 74:80:@143607.4]
  assign _T_3703 = io_wen & _T_3702; // @[RegFile.scala 74:68:@143608.4]
  assign _T_3709 = io_waddr == 11'h27; // @[RegFile.scala 74:80:@143621.4]
  assign _T_3710 = io_wen & _T_3709; // @[RegFile.scala 74:68:@143622.4]
  assign _T_3716 = io_waddr == 11'h28; // @[RegFile.scala 74:80:@143635.4]
  assign _T_3717 = io_wen & _T_3716; // @[RegFile.scala 74:68:@143636.4]
  assign _T_3723 = io_waddr == 11'h29; // @[RegFile.scala 74:80:@143649.4]
  assign _T_3724 = io_wen & _T_3723; // @[RegFile.scala 74:68:@143650.4]
  assign _T_3730 = io_waddr == 11'h2a; // @[RegFile.scala 74:80:@143663.4]
  assign _T_3731 = io_wen & _T_3730; // @[RegFile.scala 74:68:@143664.4]
  assign _T_3737 = io_waddr == 11'h2b; // @[RegFile.scala 74:80:@143677.4]
  assign _T_3738 = io_wen & _T_3737; // @[RegFile.scala 74:68:@143678.4]
  assign _T_3744 = io_waddr == 11'h2c; // @[RegFile.scala 74:80:@143691.4]
  assign _T_3745 = io_wen & _T_3744; // @[RegFile.scala 74:68:@143692.4]
  assign _T_3751 = io_waddr == 11'h2d; // @[RegFile.scala 74:80:@143705.4]
  assign _T_3752 = io_wen & _T_3751; // @[RegFile.scala 74:68:@143706.4]
  assign _T_3758 = io_waddr == 11'h2e; // @[RegFile.scala 74:80:@143719.4]
  assign _T_3759 = io_wen & _T_3758; // @[RegFile.scala 74:68:@143720.4]
  assign _T_3765 = io_waddr == 11'h2f; // @[RegFile.scala 74:80:@143733.4]
  assign _T_3766 = io_wen & _T_3765; // @[RegFile.scala 74:68:@143734.4]
  assign _T_3772 = io_waddr == 11'h30; // @[RegFile.scala 74:80:@143747.4]
  assign _T_3773 = io_wen & _T_3772; // @[RegFile.scala 74:68:@143748.4]
  assign _T_3779 = io_waddr == 11'h31; // @[RegFile.scala 74:80:@143761.4]
  assign _T_3780 = io_wen & _T_3779; // @[RegFile.scala 74:68:@143762.4]
  assign _T_3786 = io_waddr == 11'h32; // @[RegFile.scala 74:80:@143775.4]
  assign _T_3787 = io_wen & _T_3786; // @[RegFile.scala 74:68:@143776.4]
  assign _T_3793 = io_waddr == 11'h33; // @[RegFile.scala 74:80:@143789.4]
  assign _T_3794 = io_wen & _T_3793; // @[RegFile.scala 74:68:@143790.4]
  assign _T_3800 = io_waddr == 11'h34; // @[RegFile.scala 74:80:@143803.4]
  assign _T_3801 = io_wen & _T_3800; // @[RegFile.scala 74:68:@143804.4]
  assign _T_3807 = io_waddr == 11'h35; // @[RegFile.scala 74:80:@143817.4]
  assign _T_3808 = io_wen & _T_3807; // @[RegFile.scala 74:68:@143818.4]
  assign _T_3814 = io_waddr == 11'h36; // @[RegFile.scala 74:80:@143831.4]
  assign _T_3815 = io_wen & _T_3814; // @[RegFile.scala 74:68:@143832.4]
  assign _T_3821 = io_waddr == 11'h37; // @[RegFile.scala 74:80:@143845.4]
  assign _T_3822 = io_wen & _T_3821; // @[RegFile.scala 74:68:@143846.4]
  assign _T_3828 = io_waddr == 11'h38; // @[RegFile.scala 74:80:@143859.4]
  assign _T_3829 = io_wen & _T_3828; // @[RegFile.scala 74:68:@143860.4]
  assign _T_3835 = io_waddr == 11'h39; // @[RegFile.scala 74:80:@143873.4]
  assign _T_3836 = io_wen & _T_3835; // @[RegFile.scala 74:68:@143874.4]
  assign _T_3842 = io_waddr == 11'h3a; // @[RegFile.scala 74:80:@143887.4]
  assign _T_3843 = io_wen & _T_3842; // @[RegFile.scala 74:68:@143888.4]
  assign _T_3849 = io_waddr == 11'h3b; // @[RegFile.scala 74:80:@143901.4]
  assign _T_3850 = io_wen & _T_3849; // @[RegFile.scala 74:68:@143902.4]
  assign _T_3856 = io_waddr == 11'h3c; // @[RegFile.scala 74:80:@143915.4]
  assign _T_3857 = io_wen & _T_3856; // @[RegFile.scala 74:68:@143916.4]
  assign _T_3863 = io_waddr == 11'h3d; // @[RegFile.scala 74:80:@143929.4]
  assign _T_3864 = io_wen & _T_3863; // @[RegFile.scala 74:68:@143930.4]
  assign _T_3870 = io_waddr == 11'h3e; // @[RegFile.scala 74:80:@143943.4]
  assign _T_3871 = io_wen & _T_3870; // @[RegFile.scala 74:68:@143944.4]
  assign _T_3877 = io_waddr == 11'h3f; // @[RegFile.scala 74:80:@143957.4]
  assign _T_3878 = io_wen & _T_3877; // @[RegFile.scala 74:68:@143958.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@152069.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@152075.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@152076.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@152077.4]
  assign io_argIns_3 = regs_3_io_out; // @[RegFile.scala 111:13:@152078.4]
  assign io_argEchos_1 = regs_4_io_out; // @[RegFile.scala 77:37:@143138.4]
  assign io_argEchos_2 = regs_5_io_out; // @[RegFile.scala 77:37:@143152.4]
  assign io_argEchos_3 = regs_6_io_out; // @[RegFile.scala 77:37:@143166.4]
  assign io_argEchos_4 = regs_7_io_out; // @[RegFile.scala 77:37:@143180.4]
  assign io_argEchos_5 = regs_8_io_out; // @[RegFile.scala 77:37:@143194.4]
  assign io_argEchos_6 = regs_9_io_out; // @[RegFile.scala 77:37:@143208.4]
  assign io_argEchos_7 = regs_10_io_out; // @[RegFile.scala 77:37:@143222.4]
  assign io_argEchos_8 = regs_11_io_out; // @[RegFile.scala 77:37:@143236.4]
  assign io_argEchos_9 = regs_12_io_out; // @[RegFile.scala 77:37:@143250.4]
  assign io_argEchos_10 = regs_13_io_out; // @[RegFile.scala 77:37:@143264.4]
  assign io_argEchos_11 = regs_14_io_out; // @[RegFile.scala 77:37:@143278.4]
  assign io_argEchos_12 = regs_15_io_out; // @[RegFile.scala 77:37:@143292.4]
  assign io_argEchos_13 = regs_16_io_out; // @[RegFile.scala 77:37:@143306.4]
  assign io_argEchos_14 = regs_17_io_out; // @[RegFile.scala 77:37:@143320.4]
  assign io_argEchos_15 = regs_18_io_out; // @[RegFile.scala 77:37:@143334.4]
  assign io_argEchos_16 = regs_19_io_out; // @[RegFile.scala 77:37:@143348.4]
  assign io_argEchos_17 = regs_20_io_out; // @[RegFile.scala 77:37:@143362.4]
  assign io_argEchos_18 = regs_21_io_out; // @[RegFile.scala 77:37:@143376.4]
  assign io_argEchos_19 = regs_22_io_out; // @[RegFile.scala 77:37:@143390.4]
  assign io_argEchos_20 = regs_23_io_out; // @[RegFile.scala 77:37:@143404.4]
  assign io_argEchos_21 = regs_24_io_out; // @[RegFile.scala 77:37:@143418.4]
  assign io_argEchos_22 = regs_25_io_out; // @[RegFile.scala 77:37:@143432.4]
  assign io_argEchos_23 = regs_26_io_out; // @[RegFile.scala 77:37:@143446.4]
  assign io_argEchos_24 = regs_27_io_out; // @[RegFile.scala 77:37:@143460.4]
  assign io_argEchos_25 = regs_28_io_out; // @[RegFile.scala 77:37:@143474.4]
  assign io_argEchos_26 = regs_29_io_out; // @[RegFile.scala 77:37:@143488.4]
  assign io_argEchos_27 = regs_30_io_out; // @[RegFile.scala 77:37:@143502.4]
  assign io_argEchos_28 = regs_31_io_out; // @[RegFile.scala 77:37:@143516.4]
  assign io_argEchos_29 = regs_32_io_out; // @[RegFile.scala 77:37:@143530.4]
  assign io_argEchos_30 = regs_33_io_out; // @[RegFile.scala 77:37:@143544.4]
  assign io_argEchos_31 = regs_34_io_out; // @[RegFile.scala 77:37:@143558.4]
  assign io_argEchos_32 = regs_35_io_out; // @[RegFile.scala 77:37:@143572.4]
  assign io_argEchos_33 = regs_36_io_out; // @[RegFile.scala 77:37:@143586.4]
  assign io_argEchos_34 = regs_37_io_out; // @[RegFile.scala 77:37:@143600.4]
  assign io_argEchos_35 = regs_38_io_out; // @[RegFile.scala 77:37:@143614.4]
  assign io_argEchos_36 = regs_39_io_out; // @[RegFile.scala 77:37:@143628.4]
  assign io_argEchos_37 = regs_40_io_out; // @[RegFile.scala 77:37:@143642.4]
  assign io_argEchos_38 = regs_41_io_out; // @[RegFile.scala 77:37:@143656.4]
  assign io_argEchos_39 = regs_42_io_out; // @[RegFile.scala 77:37:@143670.4]
  assign io_argEchos_40 = regs_43_io_out; // @[RegFile.scala 77:37:@143684.4]
  assign io_argEchos_41 = regs_44_io_out; // @[RegFile.scala 77:37:@143698.4]
  assign io_argEchos_42 = regs_45_io_out; // @[RegFile.scala 77:37:@143712.4]
  assign io_argEchos_43 = regs_46_io_out; // @[RegFile.scala 77:37:@143726.4]
  assign io_argEchos_44 = regs_47_io_out; // @[RegFile.scala 77:37:@143740.4]
  assign io_argEchos_45 = regs_48_io_out; // @[RegFile.scala 77:37:@143754.4]
  assign io_argEchos_46 = regs_49_io_out; // @[RegFile.scala 77:37:@143768.4]
  assign io_argEchos_47 = regs_50_io_out; // @[RegFile.scala 77:37:@143782.4]
  assign io_argEchos_48 = regs_51_io_out; // @[RegFile.scala 77:37:@143796.4]
  assign io_argEchos_49 = regs_52_io_out; // @[RegFile.scala 77:37:@143810.4]
  assign io_argEchos_50 = regs_53_io_out; // @[RegFile.scala 77:37:@143824.4]
  assign io_argEchos_51 = regs_54_io_out; // @[RegFile.scala 77:37:@143838.4]
  assign io_argEchos_52 = regs_55_io_out; // @[RegFile.scala 77:37:@143852.4]
  assign io_argEchos_53 = regs_56_io_out; // @[RegFile.scala 77:37:@143866.4]
  assign io_argEchos_54 = regs_57_io_out; // @[RegFile.scala 77:37:@143880.4]
  assign io_argEchos_55 = regs_58_io_out; // @[RegFile.scala 77:37:@143894.4]
  assign io_argEchos_56 = regs_59_io_out; // @[RegFile.scala 77:37:@143908.4]
  assign io_argEchos_57 = regs_60_io_out; // @[RegFile.scala 77:37:@143922.4]
  assign io_argEchos_58 = regs_61_io_out; // @[RegFile.scala 77:37:@143936.4]
  assign io_argEchos_59 = regs_62_io_out; // @[RegFile.scala 77:37:@143950.4]
  assign io_argEchos_60 = regs_63_io_out; // @[RegFile.scala 77:37:@143964.4]
  assign regs_0_clock = clock; // @[:@143074.4]
  assign regs_0_reset = reset; // @[:@143075.4 RegFile.scala 82:16:@143081.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@143079.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@143083.4]
  assign regs_0_io_enable = io_wen & _T_3432; // @[RegFile.scala 80:20:@143078.4]
  assign regs_1_clock = clock; // @[:@143086.4]
  assign regs_1_reset = reset; // @[:@143087.4 RegFile.scala 70:16:@143099.4]
  assign regs_1_io_in = _T_3439 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@143097.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@143102.4]
  assign regs_1_io_enable = _T_3439 ? _T_3439 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@143093.4]
  assign regs_2_clock = clock; // @[:@143105.4]
  assign regs_2_reset = reset; // @[:@143106.4 RegFile.scala 82:16:@143112.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@143110.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@143114.4]
  assign regs_2_io_enable = io_wen & _T_3452; // @[RegFile.scala 80:20:@143109.4]
  assign regs_3_clock = clock; // @[:@143117.4]
  assign regs_3_reset = reset; // @[:@143118.4 RegFile.scala 82:16:@143124.4]
  assign regs_3_io_in = io_wdata; // @[RegFile.scala 81:16:@143122.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 83:19:@143126.4]
  assign regs_3_io_enable = io_wen & _T_3458; // @[RegFile.scala 80:20:@143121.4]
  assign regs_4_clock = clock; // @[:@143129.4]
  assign regs_4_reset = io_reset; // @[:@143130.4 RegFile.scala 76:16:@143137.4]
  assign regs_4_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@143136.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@143140.4]
  assign regs_4_io_enable = io_argOuts_1_valid | _T_3465; // @[RegFile.scala 74:20:@143134.4]
  assign regs_5_clock = clock; // @[:@143143.4]
  assign regs_5_reset = io_reset; // @[:@143144.4 RegFile.scala 76:16:@143151.4]
  assign regs_5_io_in = io_argOuts_2_valid ? io_argOuts_2_bits : io_wdata; // @[RegFile.scala 75:16:@143150.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@143154.4]
  assign regs_5_io_enable = io_argOuts_2_valid | _T_3472; // @[RegFile.scala 74:20:@143148.4]
  assign regs_6_clock = clock; // @[:@143157.4]
  assign regs_6_reset = io_reset; // @[:@143158.4 RegFile.scala 76:16:@143165.4]
  assign regs_6_io_in = io_argOuts_3_valid ? io_argOuts_3_bits : io_wdata; // @[RegFile.scala 75:16:@143164.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@143168.4]
  assign regs_6_io_enable = io_argOuts_3_valid | _T_3479; // @[RegFile.scala 74:20:@143162.4]
  assign regs_7_clock = clock; // @[:@143171.4]
  assign regs_7_reset = io_reset; // @[:@143172.4 RegFile.scala 76:16:@143179.4]
  assign regs_7_io_in = io_argOuts_4_valid ? io_argOuts_4_bits : io_wdata; // @[RegFile.scala 75:16:@143178.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@143182.4]
  assign regs_7_io_enable = io_argOuts_4_valid | _T_3486; // @[RegFile.scala 74:20:@143176.4]
  assign regs_8_clock = clock; // @[:@143185.4]
  assign regs_8_reset = io_reset; // @[:@143186.4 RegFile.scala 76:16:@143193.4]
  assign regs_8_io_in = io_argOuts_5_valid ? io_argOuts_5_bits : io_wdata; // @[RegFile.scala 75:16:@143192.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@143196.4]
  assign regs_8_io_enable = io_argOuts_5_valid | _T_3493; // @[RegFile.scala 74:20:@143190.4]
  assign regs_9_clock = clock; // @[:@143199.4]
  assign regs_9_reset = io_reset; // @[:@143200.4 RegFile.scala 76:16:@143207.4]
  assign regs_9_io_in = io_argOuts_6_valid ? io_argOuts_6_bits : io_wdata; // @[RegFile.scala 75:16:@143206.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@143210.4]
  assign regs_9_io_enable = io_argOuts_6_valid | _T_3500; // @[RegFile.scala 74:20:@143204.4]
  assign regs_10_clock = clock; // @[:@143213.4]
  assign regs_10_reset = io_reset; // @[:@143214.4 RegFile.scala 76:16:@143221.4]
  assign regs_10_io_in = io_argOuts_7_valid ? io_argOuts_7_bits : io_wdata; // @[RegFile.scala 75:16:@143220.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@143224.4]
  assign regs_10_io_enable = io_argOuts_7_valid | _T_3507; // @[RegFile.scala 74:20:@143218.4]
  assign regs_11_clock = clock; // @[:@143227.4]
  assign regs_11_reset = io_reset; // @[:@143228.4 RegFile.scala 76:16:@143235.4]
  assign regs_11_io_in = io_argOuts_8_valid ? io_argOuts_8_bits : io_wdata; // @[RegFile.scala 75:16:@143234.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@143238.4]
  assign regs_11_io_enable = io_argOuts_8_valid | _T_3514; // @[RegFile.scala 74:20:@143232.4]
  assign regs_12_clock = clock; // @[:@143241.4]
  assign regs_12_reset = io_reset; // @[:@143242.4 RegFile.scala 76:16:@143249.4]
  assign regs_12_io_in = io_argOuts_9_valid ? io_argOuts_9_bits : io_wdata; // @[RegFile.scala 75:16:@143248.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@143252.4]
  assign regs_12_io_enable = io_argOuts_9_valid | _T_3521; // @[RegFile.scala 74:20:@143246.4]
  assign regs_13_clock = clock; // @[:@143255.4]
  assign regs_13_reset = io_reset; // @[:@143256.4 RegFile.scala 76:16:@143263.4]
  assign regs_13_io_in = io_argOuts_10_valid ? io_argOuts_10_bits : io_wdata; // @[RegFile.scala 75:16:@143262.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@143266.4]
  assign regs_13_io_enable = io_argOuts_10_valid | _T_3528; // @[RegFile.scala 74:20:@143260.4]
  assign regs_14_clock = clock; // @[:@143269.4]
  assign regs_14_reset = io_reset; // @[:@143270.4 RegFile.scala 76:16:@143277.4]
  assign regs_14_io_in = io_argOuts_11_valid ? io_argOuts_11_bits : io_wdata; // @[RegFile.scala 75:16:@143276.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@143280.4]
  assign regs_14_io_enable = io_argOuts_11_valid | _T_3535; // @[RegFile.scala 74:20:@143274.4]
  assign regs_15_clock = clock; // @[:@143283.4]
  assign regs_15_reset = io_reset; // @[:@143284.4 RegFile.scala 76:16:@143291.4]
  assign regs_15_io_in = io_argOuts_12_valid ? io_argOuts_12_bits : io_wdata; // @[RegFile.scala 75:16:@143290.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@143294.4]
  assign regs_15_io_enable = io_argOuts_12_valid | _T_3542; // @[RegFile.scala 74:20:@143288.4]
  assign regs_16_clock = clock; // @[:@143297.4]
  assign regs_16_reset = io_reset; // @[:@143298.4 RegFile.scala 76:16:@143305.4]
  assign regs_16_io_in = io_argOuts_13_valid ? io_argOuts_13_bits : io_wdata; // @[RegFile.scala 75:16:@143304.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@143308.4]
  assign regs_16_io_enable = io_argOuts_13_valid | _T_3549; // @[RegFile.scala 74:20:@143302.4]
  assign regs_17_clock = clock; // @[:@143311.4]
  assign regs_17_reset = io_reset; // @[:@143312.4 RegFile.scala 76:16:@143319.4]
  assign regs_17_io_in = io_argOuts_14_valid ? io_argOuts_14_bits : io_wdata; // @[RegFile.scala 75:16:@143318.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@143322.4]
  assign regs_17_io_enable = io_argOuts_14_valid | _T_3556; // @[RegFile.scala 74:20:@143316.4]
  assign regs_18_clock = clock; // @[:@143325.4]
  assign regs_18_reset = io_reset; // @[:@143326.4 RegFile.scala 76:16:@143333.4]
  assign regs_18_io_in = io_argOuts_15_valid ? io_argOuts_15_bits : io_wdata; // @[RegFile.scala 75:16:@143332.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@143336.4]
  assign regs_18_io_enable = io_argOuts_15_valid | _T_3563; // @[RegFile.scala 74:20:@143330.4]
  assign regs_19_clock = clock; // @[:@143339.4]
  assign regs_19_reset = io_reset; // @[:@143340.4 RegFile.scala 76:16:@143347.4]
  assign regs_19_io_in = io_argOuts_16_valid ? io_argOuts_16_bits : io_wdata; // @[RegFile.scala 75:16:@143346.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@143350.4]
  assign regs_19_io_enable = io_argOuts_16_valid | _T_3570; // @[RegFile.scala 74:20:@143344.4]
  assign regs_20_clock = clock; // @[:@143353.4]
  assign regs_20_reset = io_reset; // @[:@143354.4 RegFile.scala 76:16:@143361.4]
  assign regs_20_io_in = io_argOuts_17_valid ? io_argOuts_17_bits : io_wdata; // @[RegFile.scala 75:16:@143360.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@143364.4]
  assign regs_20_io_enable = io_argOuts_17_valid | _T_3577; // @[RegFile.scala 74:20:@143358.4]
  assign regs_21_clock = clock; // @[:@143367.4]
  assign regs_21_reset = io_reset; // @[:@143368.4 RegFile.scala 76:16:@143375.4]
  assign regs_21_io_in = io_argOuts_18_valid ? io_argOuts_18_bits : io_wdata; // @[RegFile.scala 75:16:@143374.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@143378.4]
  assign regs_21_io_enable = io_argOuts_18_valid | _T_3584; // @[RegFile.scala 74:20:@143372.4]
  assign regs_22_clock = clock; // @[:@143381.4]
  assign regs_22_reset = io_reset; // @[:@143382.4 RegFile.scala 76:16:@143389.4]
  assign regs_22_io_in = io_argOuts_19_valid ? io_argOuts_19_bits : io_wdata; // @[RegFile.scala 75:16:@143388.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@143392.4]
  assign regs_22_io_enable = io_argOuts_19_valid | _T_3591; // @[RegFile.scala 74:20:@143386.4]
  assign regs_23_clock = clock; // @[:@143395.4]
  assign regs_23_reset = io_reset; // @[:@143396.4 RegFile.scala 76:16:@143403.4]
  assign regs_23_io_in = io_argOuts_20_valid ? io_argOuts_20_bits : io_wdata; // @[RegFile.scala 75:16:@143402.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@143406.4]
  assign regs_23_io_enable = io_argOuts_20_valid | _T_3598; // @[RegFile.scala 74:20:@143400.4]
  assign regs_24_clock = clock; // @[:@143409.4]
  assign regs_24_reset = io_reset; // @[:@143410.4 RegFile.scala 76:16:@143417.4]
  assign regs_24_io_in = io_argOuts_21_valid ? io_argOuts_21_bits : io_wdata; // @[RegFile.scala 75:16:@143416.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@143420.4]
  assign regs_24_io_enable = io_argOuts_21_valid | _T_3605; // @[RegFile.scala 74:20:@143414.4]
  assign regs_25_clock = clock; // @[:@143423.4]
  assign regs_25_reset = io_reset; // @[:@143424.4 RegFile.scala 76:16:@143431.4]
  assign regs_25_io_in = io_argOuts_22_valid ? io_argOuts_22_bits : io_wdata; // @[RegFile.scala 75:16:@143430.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@143434.4]
  assign regs_25_io_enable = io_argOuts_22_valid | _T_3612; // @[RegFile.scala 74:20:@143428.4]
  assign regs_26_clock = clock; // @[:@143437.4]
  assign regs_26_reset = io_reset; // @[:@143438.4 RegFile.scala 76:16:@143445.4]
  assign regs_26_io_in = io_argOuts_23_valid ? io_argOuts_23_bits : io_wdata; // @[RegFile.scala 75:16:@143444.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@143448.4]
  assign regs_26_io_enable = io_argOuts_23_valid | _T_3619; // @[RegFile.scala 74:20:@143442.4]
  assign regs_27_clock = clock; // @[:@143451.4]
  assign regs_27_reset = io_reset; // @[:@143452.4 RegFile.scala 76:16:@143459.4]
  assign regs_27_io_in = io_argOuts_24_valid ? io_argOuts_24_bits : io_wdata; // @[RegFile.scala 75:16:@143458.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@143462.4]
  assign regs_27_io_enable = io_argOuts_24_valid | _T_3626; // @[RegFile.scala 74:20:@143456.4]
  assign regs_28_clock = clock; // @[:@143465.4]
  assign regs_28_reset = io_reset; // @[:@143466.4 RegFile.scala 76:16:@143473.4]
  assign regs_28_io_in = io_argOuts_25_valid ? io_argOuts_25_bits : io_wdata; // @[RegFile.scala 75:16:@143472.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@143476.4]
  assign regs_28_io_enable = io_argOuts_25_valid | _T_3633; // @[RegFile.scala 74:20:@143470.4]
  assign regs_29_clock = clock; // @[:@143479.4]
  assign regs_29_reset = io_reset; // @[:@143480.4 RegFile.scala 76:16:@143487.4]
  assign regs_29_io_in = io_argOuts_26_valid ? io_argOuts_26_bits : io_wdata; // @[RegFile.scala 75:16:@143486.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@143490.4]
  assign regs_29_io_enable = io_argOuts_26_valid | _T_3640; // @[RegFile.scala 74:20:@143484.4]
  assign regs_30_clock = clock; // @[:@143493.4]
  assign regs_30_reset = io_reset; // @[:@143494.4 RegFile.scala 76:16:@143501.4]
  assign regs_30_io_in = io_argOuts_27_valid ? io_argOuts_27_bits : io_wdata; // @[RegFile.scala 75:16:@143500.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@143504.4]
  assign regs_30_io_enable = io_argOuts_27_valid | _T_3647; // @[RegFile.scala 74:20:@143498.4]
  assign regs_31_clock = clock; // @[:@143507.4]
  assign regs_31_reset = io_reset; // @[:@143508.4 RegFile.scala 76:16:@143515.4]
  assign regs_31_io_in = io_argOuts_28_valid ? io_argOuts_28_bits : io_wdata; // @[RegFile.scala 75:16:@143514.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@143518.4]
  assign regs_31_io_enable = io_argOuts_28_valid | _T_3654; // @[RegFile.scala 74:20:@143512.4]
  assign regs_32_clock = clock; // @[:@143521.4]
  assign regs_32_reset = io_reset; // @[:@143522.4 RegFile.scala 76:16:@143529.4]
  assign regs_32_io_in = io_argOuts_29_valid ? io_argOuts_29_bits : io_wdata; // @[RegFile.scala 75:16:@143528.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@143532.4]
  assign regs_32_io_enable = io_argOuts_29_valid | _T_3661; // @[RegFile.scala 74:20:@143526.4]
  assign regs_33_clock = clock; // @[:@143535.4]
  assign regs_33_reset = io_reset; // @[:@143536.4 RegFile.scala 76:16:@143543.4]
  assign regs_33_io_in = io_argOuts_30_valid ? io_argOuts_30_bits : io_wdata; // @[RegFile.scala 75:16:@143542.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@143546.4]
  assign regs_33_io_enable = io_argOuts_30_valid | _T_3668; // @[RegFile.scala 74:20:@143540.4]
  assign regs_34_clock = clock; // @[:@143549.4]
  assign regs_34_reset = io_reset; // @[:@143550.4 RegFile.scala 76:16:@143557.4]
  assign regs_34_io_in = io_argOuts_31_valid ? io_argOuts_31_bits : io_wdata; // @[RegFile.scala 75:16:@143556.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@143560.4]
  assign regs_34_io_enable = io_argOuts_31_valid | _T_3675; // @[RegFile.scala 74:20:@143554.4]
  assign regs_35_clock = clock; // @[:@143563.4]
  assign regs_35_reset = io_reset; // @[:@143564.4 RegFile.scala 76:16:@143571.4]
  assign regs_35_io_in = io_argOuts_32_valid ? io_argOuts_32_bits : io_wdata; // @[RegFile.scala 75:16:@143570.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@143574.4]
  assign regs_35_io_enable = io_argOuts_32_valid | _T_3682; // @[RegFile.scala 74:20:@143568.4]
  assign regs_36_clock = clock; // @[:@143577.4]
  assign regs_36_reset = io_reset; // @[:@143578.4 RegFile.scala 76:16:@143585.4]
  assign regs_36_io_in = io_argOuts_33_valid ? io_argOuts_33_bits : io_wdata; // @[RegFile.scala 75:16:@143584.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@143588.4]
  assign regs_36_io_enable = io_argOuts_33_valid | _T_3689; // @[RegFile.scala 74:20:@143582.4]
  assign regs_37_clock = clock; // @[:@143591.4]
  assign regs_37_reset = io_reset; // @[:@143592.4 RegFile.scala 76:16:@143599.4]
  assign regs_37_io_in = io_argOuts_34_valid ? io_argOuts_34_bits : io_wdata; // @[RegFile.scala 75:16:@143598.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@143602.4]
  assign regs_37_io_enable = io_argOuts_34_valid | _T_3696; // @[RegFile.scala 74:20:@143596.4]
  assign regs_38_clock = clock; // @[:@143605.4]
  assign regs_38_reset = io_reset; // @[:@143606.4 RegFile.scala 76:16:@143613.4]
  assign regs_38_io_in = io_argOuts_35_valid ? io_argOuts_35_bits : io_wdata; // @[RegFile.scala 75:16:@143612.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@143616.4]
  assign regs_38_io_enable = io_argOuts_35_valid | _T_3703; // @[RegFile.scala 74:20:@143610.4]
  assign regs_39_clock = clock; // @[:@143619.4]
  assign regs_39_reset = io_reset; // @[:@143620.4 RegFile.scala 76:16:@143627.4]
  assign regs_39_io_in = io_argOuts_36_valid ? io_argOuts_36_bits : io_wdata; // @[RegFile.scala 75:16:@143626.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@143630.4]
  assign regs_39_io_enable = io_argOuts_36_valid | _T_3710; // @[RegFile.scala 74:20:@143624.4]
  assign regs_40_clock = clock; // @[:@143633.4]
  assign regs_40_reset = io_reset; // @[:@143634.4 RegFile.scala 76:16:@143641.4]
  assign regs_40_io_in = io_argOuts_37_valid ? io_argOuts_37_bits : io_wdata; // @[RegFile.scala 75:16:@143640.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@143644.4]
  assign regs_40_io_enable = io_argOuts_37_valid | _T_3717; // @[RegFile.scala 74:20:@143638.4]
  assign regs_41_clock = clock; // @[:@143647.4]
  assign regs_41_reset = io_reset; // @[:@143648.4 RegFile.scala 76:16:@143655.4]
  assign regs_41_io_in = io_argOuts_38_valid ? io_argOuts_38_bits : io_wdata; // @[RegFile.scala 75:16:@143654.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@143658.4]
  assign regs_41_io_enable = io_argOuts_38_valid | _T_3724; // @[RegFile.scala 74:20:@143652.4]
  assign regs_42_clock = clock; // @[:@143661.4]
  assign regs_42_reset = io_reset; // @[:@143662.4 RegFile.scala 76:16:@143669.4]
  assign regs_42_io_in = io_argOuts_39_valid ? io_argOuts_39_bits : io_wdata; // @[RegFile.scala 75:16:@143668.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@143672.4]
  assign regs_42_io_enable = io_argOuts_39_valid | _T_3731; // @[RegFile.scala 74:20:@143666.4]
  assign regs_43_clock = clock; // @[:@143675.4]
  assign regs_43_reset = io_reset; // @[:@143676.4 RegFile.scala 76:16:@143683.4]
  assign regs_43_io_in = io_argOuts_40_valid ? io_argOuts_40_bits : io_wdata; // @[RegFile.scala 75:16:@143682.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@143686.4]
  assign regs_43_io_enable = io_argOuts_40_valid | _T_3738; // @[RegFile.scala 74:20:@143680.4]
  assign regs_44_clock = clock; // @[:@143689.4]
  assign regs_44_reset = io_reset; // @[:@143690.4 RegFile.scala 76:16:@143697.4]
  assign regs_44_io_in = io_argOuts_41_valid ? io_argOuts_41_bits : io_wdata; // @[RegFile.scala 75:16:@143696.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@143700.4]
  assign regs_44_io_enable = io_argOuts_41_valid | _T_3745; // @[RegFile.scala 74:20:@143694.4]
  assign regs_45_clock = clock; // @[:@143703.4]
  assign regs_45_reset = io_reset; // @[:@143704.4 RegFile.scala 76:16:@143711.4]
  assign regs_45_io_in = io_argOuts_42_valid ? io_argOuts_42_bits : io_wdata; // @[RegFile.scala 75:16:@143710.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@143714.4]
  assign regs_45_io_enable = io_argOuts_42_valid | _T_3752; // @[RegFile.scala 74:20:@143708.4]
  assign regs_46_clock = clock; // @[:@143717.4]
  assign regs_46_reset = io_reset; // @[:@143718.4 RegFile.scala 76:16:@143725.4]
  assign regs_46_io_in = io_argOuts_43_valid ? io_argOuts_43_bits : io_wdata; // @[RegFile.scala 75:16:@143724.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@143728.4]
  assign regs_46_io_enable = io_argOuts_43_valid | _T_3759; // @[RegFile.scala 74:20:@143722.4]
  assign regs_47_clock = clock; // @[:@143731.4]
  assign regs_47_reset = io_reset; // @[:@143732.4 RegFile.scala 76:16:@143739.4]
  assign regs_47_io_in = io_argOuts_44_valid ? io_argOuts_44_bits : io_wdata; // @[RegFile.scala 75:16:@143738.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@143742.4]
  assign regs_47_io_enable = io_argOuts_44_valid | _T_3766; // @[RegFile.scala 74:20:@143736.4]
  assign regs_48_clock = clock; // @[:@143745.4]
  assign regs_48_reset = io_reset; // @[:@143746.4 RegFile.scala 76:16:@143753.4]
  assign regs_48_io_in = io_argOuts_45_valid ? io_argOuts_45_bits : io_wdata; // @[RegFile.scala 75:16:@143752.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@143756.4]
  assign regs_48_io_enable = io_argOuts_45_valid | _T_3773; // @[RegFile.scala 74:20:@143750.4]
  assign regs_49_clock = clock; // @[:@143759.4]
  assign regs_49_reset = io_reset; // @[:@143760.4 RegFile.scala 76:16:@143767.4]
  assign regs_49_io_in = io_argOuts_46_valid ? io_argOuts_46_bits : io_wdata; // @[RegFile.scala 75:16:@143766.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@143770.4]
  assign regs_49_io_enable = io_argOuts_46_valid | _T_3780; // @[RegFile.scala 74:20:@143764.4]
  assign regs_50_clock = clock; // @[:@143773.4]
  assign regs_50_reset = io_reset; // @[:@143774.4 RegFile.scala 76:16:@143781.4]
  assign regs_50_io_in = io_argOuts_47_valid ? io_argOuts_47_bits : io_wdata; // @[RegFile.scala 75:16:@143780.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@143784.4]
  assign regs_50_io_enable = io_argOuts_47_valid | _T_3787; // @[RegFile.scala 74:20:@143778.4]
  assign regs_51_clock = clock; // @[:@143787.4]
  assign regs_51_reset = io_reset; // @[:@143788.4 RegFile.scala 76:16:@143795.4]
  assign regs_51_io_in = io_argOuts_48_valid ? io_argOuts_48_bits : io_wdata; // @[RegFile.scala 75:16:@143794.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@143798.4]
  assign regs_51_io_enable = io_argOuts_48_valid | _T_3794; // @[RegFile.scala 74:20:@143792.4]
  assign regs_52_clock = clock; // @[:@143801.4]
  assign regs_52_reset = io_reset; // @[:@143802.4 RegFile.scala 76:16:@143809.4]
  assign regs_52_io_in = io_argOuts_49_valid ? io_argOuts_49_bits : io_wdata; // @[RegFile.scala 75:16:@143808.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@143812.4]
  assign regs_52_io_enable = io_argOuts_49_valid | _T_3801; // @[RegFile.scala 74:20:@143806.4]
  assign regs_53_clock = clock; // @[:@143815.4]
  assign regs_53_reset = io_reset; // @[:@143816.4 RegFile.scala 76:16:@143823.4]
  assign regs_53_io_in = io_argOuts_50_valid ? io_argOuts_50_bits : io_wdata; // @[RegFile.scala 75:16:@143822.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@143826.4]
  assign regs_53_io_enable = io_argOuts_50_valid | _T_3808; // @[RegFile.scala 74:20:@143820.4]
  assign regs_54_clock = clock; // @[:@143829.4]
  assign regs_54_reset = io_reset; // @[:@143830.4 RegFile.scala 76:16:@143837.4]
  assign regs_54_io_in = io_argOuts_51_valid ? io_argOuts_51_bits : io_wdata; // @[RegFile.scala 75:16:@143836.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@143840.4]
  assign regs_54_io_enable = io_argOuts_51_valid | _T_3815; // @[RegFile.scala 74:20:@143834.4]
  assign regs_55_clock = clock; // @[:@143843.4]
  assign regs_55_reset = io_reset; // @[:@143844.4 RegFile.scala 76:16:@143851.4]
  assign regs_55_io_in = io_argOuts_52_valid ? io_argOuts_52_bits : io_wdata; // @[RegFile.scala 75:16:@143850.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@143854.4]
  assign regs_55_io_enable = io_argOuts_52_valid | _T_3822; // @[RegFile.scala 74:20:@143848.4]
  assign regs_56_clock = clock; // @[:@143857.4]
  assign regs_56_reset = io_reset; // @[:@143858.4 RegFile.scala 76:16:@143865.4]
  assign regs_56_io_in = io_argOuts_53_valid ? io_argOuts_53_bits : io_wdata; // @[RegFile.scala 75:16:@143864.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@143868.4]
  assign regs_56_io_enable = io_argOuts_53_valid | _T_3829; // @[RegFile.scala 74:20:@143862.4]
  assign regs_57_clock = clock; // @[:@143871.4]
  assign regs_57_reset = io_reset; // @[:@143872.4 RegFile.scala 76:16:@143879.4]
  assign regs_57_io_in = io_argOuts_54_valid ? io_argOuts_54_bits : io_wdata; // @[RegFile.scala 75:16:@143878.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@143882.4]
  assign regs_57_io_enable = io_argOuts_54_valid | _T_3836; // @[RegFile.scala 74:20:@143876.4]
  assign regs_58_clock = clock; // @[:@143885.4]
  assign regs_58_reset = io_reset; // @[:@143886.4 RegFile.scala 76:16:@143893.4]
  assign regs_58_io_in = io_argOuts_55_valid ? io_argOuts_55_bits : io_wdata; // @[RegFile.scala 75:16:@143892.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@143896.4]
  assign regs_58_io_enable = io_argOuts_55_valid | _T_3843; // @[RegFile.scala 74:20:@143890.4]
  assign regs_59_clock = clock; // @[:@143899.4]
  assign regs_59_reset = io_reset; // @[:@143900.4 RegFile.scala 76:16:@143907.4]
  assign regs_59_io_in = io_argOuts_56_valid ? io_argOuts_56_bits : io_wdata; // @[RegFile.scala 75:16:@143906.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@143910.4]
  assign regs_59_io_enable = io_argOuts_56_valid | _T_3850; // @[RegFile.scala 74:20:@143904.4]
  assign regs_60_clock = clock; // @[:@143913.4]
  assign regs_60_reset = io_reset; // @[:@143914.4 RegFile.scala 76:16:@143921.4]
  assign regs_60_io_in = io_argOuts_57_valid ? io_argOuts_57_bits : io_wdata; // @[RegFile.scala 75:16:@143920.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@143924.4]
  assign regs_60_io_enable = io_argOuts_57_valid | _T_3857; // @[RegFile.scala 74:20:@143918.4]
  assign regs_61_clock = clock; // @[:@143927.4]
  assign regs_61_reset = io_reset; // @[:@143928.4 RegFile.scala 76:16:@143935.4]
  assign regs_61_io_in = io_argOuts_58_valid ? io_argOuts_58_bits : io_wdata; // @[RegFile.scala 75:16:@143934.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@143938.4]
  assign regs_61_io_enable = io_argOuts_58_valid | _T_3864; // @[RegFile.scala 74:20:@143932.4]
  assign regs_62_clock = clock; // @[:@143941.4]
  assign regs_62_reset = io_reset; // @[:@143942.4 RegFile.scala 76:16:@143949.4]
  assign regs_62_io_in = io_argOuts_59_valid ? io_argOuts_59_bits : io_wdata; // @[RegFile.scala 75:16:@143948.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@143952.4]
  assign regs_62_io_enable = io_argOuts_59_valid | _T_3871; // @[RegFile.scala 74:20:@143946.4]
  assign regs_63_clock = clock; // @[:@143955.4]
  assign regs_63_reset = io_reset; // @[:@143956.4 RegFile.scala 76:16:@143963.4]
  assign regs_63_io_in = io_argOuts_60_valid ? io_argOuts_60_bits : io_wdata; // @[RegFile.scala 75:16:@143962.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@143966.4]
  assign regs_63_io_enable = io_argOuts_60_valid | _T_3878; // @[RegFile.scala 74:20:@143960.4]
  assign regs_64_clock = clock; // @[:@143969.4]
  assign regs_64_reset = io_reset; // @[:@143970.4 RegFile.scala 76:16:@143977.4]
  assign regs_64_io_in = io_argOuts_61_bits; // @[RegFile.scala 75:16:@143976.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@143980.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@143974.4]
  assign regs_65_clock = clock; // @[:@143983.4]
  assign regs_65_reset = io_reset; // @[:@143984.4 RegFile.scala 76:16:@143991.4]
  assign regs_65_io_in = io_argOuts_62_bits; // @[RegFile.scala 75:16:@143990.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@143994.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@143988.4]
  assign regs_66_clock = clock; // @[:@143997.4]
  assign regs_66_reset = io_reset; // @[:@143998.4 RegFile.scala 76:16:@144005.4]
  assign regs_66_io_in = io_argOuts_63_bits; // @[RegFile.scala 75:16:@144004.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@144008.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@144002.4]
  assign regs_67_clock = clock; // @[:@144011.4]
  assign regs_67_reset = io_reset; // @[:@144012.4 RegFile.scala 76:16:@144019.4]
  assign regs_67_io_in = io_argOuts_64_bits; // @[RegFile.scala 75:16:@144018.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@144022.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@144016.4]
  assign regs_68_clock = clock; // @[:@144025.4]
  assign regs_68_reset = io_reset; // @[:@144026.4 RegFile.scala 76:16:@144033.4]
  assign regs_68_io_in = io_argOuts_65_bits; // @[RegFile.scala 75:16:@144032.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@144036.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@144030.4]
  assign regs_69_clock = clock; // @[:@144039.4]
  assign regs_69_reset = io_reset; // @[:@144040.4 RegFile.scala 76:16:@144047.4]
  assign regs_69_io_in = io_argOuts_66_bits; // @[RegFile.scala 75:16:@144046.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@144050.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@144044.4]
  assign regs_70_clock = clock; // @[:@144053.4]
  assign regs_70_reset = io_reset; // @[:@144054.4 RegFile.scala 76:16:@144061.4]
  assign regs_70_io_in = io_argOuts_67_bits; // @[RegFile.scala 75:16:@144060.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@144064.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@144058.4]
  assign regs_71_clock = clock; // @[:@144067.4]
  assign regs_71_reset = io_reset; // @[:@144068.4 RegFile.scala 76:16:@144075.4]
  assign regs_71_io_in = io_argOuts_68_bits; // @[RegFile.scala 75:16:@144074.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@144078.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@144072.4]
  assign regs_72_clock = clock; // @[:@144081.4]
  assign regs_72_reset = io_reset; // @[:@144082.4 RegFile.scala 76:16:@144089.4]
  assign regs_72_io_in = io_argOuts_69_bits; // @[RegFile.scala 75:16:@144088.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@144092.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@144086.4]
  assign regs_73_clock = clock; // @[:@144095.4]
  assign regs_73_reset = io_reset; // @[:@144096.4 RegFile.scala 76:16:@144103.4]
  assign regs_73_io_in = io_argOuts_70_bits; // @[RegFile.scala 75:16:@144102.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@144106.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@144100.4]
  assign regs_74_clock = clock; // @[:@144109.4]
  assign regs_74_reset = io_reset; // @[:@144110.4 RegFile.scala 76:16:@144117.4]
  assign regs_74_io_in = io_argOuts_71_bits; // @[RegFile.scala 75:16:@144116.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@144120.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@144114.4]
  assign regs_75_clock = clock; // @[:@144123.4]
  assign regs_75_reset = io_reset; // @[:@144124.4 RegFile.scala 76:16:@144131.4]
  assign regs_75_io_in = io_argOuts_72_bits; // @[RegFile.scala 75:16:@144130.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@144134.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@144128.4]
  assign regs_76_clock = clock; // @[:@144137.4]
  assign regs_76_reset = io_reset; // @[:@144138.4 RegFile.scala 76:16:@144145.4]
  assign regs_76_io_in = io_argOuts_73_bits; // @[RegFile.scala 75:16:@144144.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@144148.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@144142.4]
  assign regs_77_clock = clock; // @[:@144151.4]
  assign regs_77_reset = io_reset; // @[:@144152.4 RegFile.scala 76:16:@144159.4]
  assign regs_77_io_in = io_argOuts_74_bits; // @[RegFile.scala 75:16:@144158.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@144162.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@144156.4]
  assign regs_78_clock = clock; // @[:@144165.4]
  assign regs_78_reset = io_reset; // @[:@144166.4 RegFile.scala 76:16:@144173.4]
  assign regs_78_io_in = io_argOuts_75_bits; // @[RegFile.scala 75:16:@144172.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@144176.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@144170.4]
  assign regs_79_clock = clock; // @[:@144179.4]
  assign regs_79_reset = io_reset; // @[:@144180.4 RegFile.scala 76:16:@144187.4]
  assign regs_79_io_in = io_argOuts_76_bits; // @[RegFile.scala 75:16:@144186.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@144190.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@144184.4]
  assign regs_80_clock = clock; // @[:@144193.4]
  assign regs_80_reset = io_reset; // @[:@144194.4 RegFile.scala 76:16:@144201.4]
  assign regs_80_io_in = io_argOuts_77_bits; // @[RegFile.scala 75:16:@144200.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@144204.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@144198.4]
  assign regs_81_clock = clock; // @[:@144207.4]
  assign regs_81_reset = io_reset; // @[:@144208.4 RegFile.scala 76:16:@144215.4]
  assign regs_81_io_in = io_argOuts_78_bits; // @[RegFile.scala 75:16:@144214.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@144218.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@144212.4]
  assign regs_82_clock = clock; // @[:@144221.4]
  assign regs_82_reset = io_reset; // @[:@144222.4 RegFile.scala 76:16:@144229.4]
  assign regs_82_io_in = io_argOuts_79_bits; // @[RegFile.scala 75:16:@144228.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@144232.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@144226.4]
  assign regs_83_clock = clock; // @[:@144235.4]
  assign regs_83_reset = io_reset; // @[:@144236.4 RegFile.scala 76:16:@144243.4]
  assign regs_83_io_in = io_argOuts_80_bits; // @[RegFile.scala 75:16:@144242.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@144246.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@144240.4]
  assign regs_84_clock = clock; // @[:@144249.4]
  assign regs_84_reset = io_reset; // @[:@144250.4 RegFile.scala 76:16:@144257.4]
  assign regs_84_io_in = io_argOuts_81_bits; // @[RegFile.scala 75:16:@144256.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@144260.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@144254.4]
  assign regs_85_clock = clock; // @[:@144263.4]
  assign regs_85_reset = io_reset; // @[:@144264.4 RegFile.scala 76:16:@144271.4]
  assign regs_85_io_in = io_argOuts_82_bits; // @[RegFile.scala 75:16:@144270.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@144274.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@144268.4]
  assign regs_86_clock = clock; // @[:@144277.4]
  assign regs_86_reset = io_reset; // @[:@144278.4 RegFile.scala 76:16:@144285.4]
  assign regs_86_io_in = io_argOuts_83_bits; // @[RegFile.scala 75:16:@144284.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@144288.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@144282.4]
  assign regs_87_clock = clock; // @[:@144291.4]
  assign regs_87_reset = io_reset; // @[:@144292.4 RegFile.scala 76:16:@144299.4]
  assign regs_87_io_in = io_argOuts_84_bits; // @[RegFile.scala 75:16:@144298.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@144302.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@144296.4]
  assign regs_88_clock = clock; // @[:@144305.4]
  assign regs_88_reset = io_reset; // @[:@144306.4 RegFile.scala 76:16:@144313.4]
  assign regs_88_io_in = io_argOuts_85_bits; // @[RegFile.scala 75:16:@144312.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@144316.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@144310.4]
  assign regs_89_clock = clock; // @[:@144319.4]
  assign regs_89_reset = io_reset; // @[:@144320.4 RegFile.scala 76:16:@144327.4]
  assign regs_89_io_in = io_argOuts_86_bits; // @[RegFile.scala 75:16:@144326.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@144330.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@144324.4]
  assign regs_90_clock = clock; // @[:@144333.4]
  assign regs_90_reset = io_reset; // @[:@144334.4 RegFile.scala 76:16:@144341.4]
  assign regs_90_io_in = io_argOuts_87_bits; // @[RegFile.scala 75:16:@144340.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@144344.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@144338.4]
  assign regs_91_clock = clock; // @[:@144347.4]
  assign regs_91_reset = io_reset; // @[:@144348.4 RegFile.scala 76:16:@144355.4]
  assign regs_91_io_in = io_argOuts_88_bits; // @[RegFile.scala 75:16:@144354.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@144358.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@144352.4]
  assign regs_92_clock = clock; // @[:@144361.4]
  assign regs_92_reset = io_reset; // @[:@144362.4 RegFile.scala 76:16:@144369.4]
  assign regs_92_io_in = io_argOuts_89_bits; // @[RegFile.scala 75:16:@144368.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@144372.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@144366.4]
  assign regs_93_clock = clock; // @[:@144375.4]
  assign regs_93_reset = io_reset; // @[:@144376.4 RegFile.scala 76:16:@144383.4]
  assign regs_93_io_in = io_argOuts_90_bits; // @[RegFile.scala 75:16:@144382.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@144386.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@144380.4]
  assign regs_94_clock = clock; // @[:@144389.4]
  assign regs_94_reset = io_reset; // @[:@144390.4 RegFile.scala 76:16:@144397.4]
  assign regs_94_io_in = io_argOuts_91_bits; // @[RegFile.scala 75:16:@144396.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@144400.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@144394.4]
  assign regs_95_clock = clock; // @[:@144403.4]
  assign regs_95_reset = io_reset; // @[:@144404.4 RegFile.scala 76:16:@144411.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@144410.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@144414.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@144408.4]
  assign regs_96_clock = clock; // @[:@144417.4]
  assign regs_96_reset = io_reset; // @[:@144418.4 RegFile.scala 76:16:@144425.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@144424.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@144428.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@144422.4]
  assign regs_97_clock = clock; // @[:@144431.4]
  assign regs_97_reset = io_reset; // @[:@144432.4 RegFile.scala 76:16:@144439.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@144438.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@144442.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@144436.4]
  assign regs_98_clock = clock; // @[:@144445.4]
  assign regs_98_reset = io_reset; // @[:@144446.4 RegFile.scala 76:16:@144453.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@144452.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@144456.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@144450.4]
  assign regs_99_clock = clock; // @[:@144459.4]
  assign regs_99_reset = io_reset; // @[:@144460.4 RegFile.scala 76:16:@144467.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@144466.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@144470.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@144464.4]
  assign regs_100_clock = clock; // @[:@144473.4]
  assign regs_100_reset = io_reset; // @[:@144474.4 RegFile.scala 76:16:@144481.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@144480.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@144484.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@144478.4]
  assign regs_101_clock = clock; // @[:@144487.4]
  assign regs_101_reset = io_reset; // @[:@144488.4 RegFile.scala 76:16:@144495.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@144494.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@144498.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@144492.4]
  assign regs_102_clock = clock; // @[:@144501.4]
  assign regs_102_reset = io_reset; // @[:@144502.4 RegFile.scala 76:16:@144509.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@144508.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@144512.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@144506.4]
  assign regs_103_clock = clock; // @[:@144515.4]
  assign regs_103_reset = io_reset; // @[:@144516.4 RegFile.scala 76:16:@144523.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@144522.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@144526.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@144520.4]
  assign regs_104_clock = clock; // @[:@144529.4]
  assign regs_104_reset = io_reset; // @[:@144530.4 RegFile.scala 76:16:@144537.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@144536.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@144540.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@144534.4]
  assign regs_105_clock = clock; // @[:@144543.4]
  assign regs_105_reset = io_reset; // @[:@144544.4 RegFile.scala 76:16:@144551.4]
  assign regs_105_io_in = io_argOuts_102_bits; // @[RegFile.scala 75:16:@144550.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@144554.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@144548.4]
  assign regs_106_clock = clock; // @[:@144557.4]
  assign regs_106_reset = io_reset; // @[:@144558.4 RegFile.scala 76:16:@144565.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@144564.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@144568.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@144562.4]
  assign regs_107_clock = clock; // @[:@144571.4]
  assign regs_107_reset = io_reset; // @[:@144572.4 RegFile.scala 76:16:@144579.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@144578.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@144582.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@144576.4]
  assign regs_108_clock = clock; // @[:@144585.4]
  assign regs_108_reset = io_reset; // @[:@144586.4 RegFile.scala 76:16:@144593.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@144592.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@144596.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@144590.4]
  assign regs_109_clock = clock; // @[:@144599.4]
  assign regs_109_reset = io_reset; // @[:@144600.4 RegFile.scala 76:16:@144607.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@144606.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@144610.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@144604.4]
  assign regs_110_clock = clock; // @[:@144613.4]
  assign regs_110_reset = io_reset; // @[:@144614.4 RegFile.scala 76:16:@144621.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@144620.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@144624.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@144618.4]
  assign regs_111_clock = clock; // @[:@144627.4]
  assign regs_111_reset = io_reset; // @[:@144628.4 RegFile.scala 76:16:@144635.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@144634.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@144638.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@144632.4]
  assign regs_112_clock = clock; // @[:@144641.4]
  assign regs_112_reset = io_reset; // @[:@144642.4 RegFile.scala 76:16:@144649.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@144648.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@144652.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@144646.4]
  assign regs_113_clock = clock; // @[:@144655.4]
  assign regs_113_reset = io_reset; // @[:@144656.4 RegFile.scala 76:16:@144663.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@144662.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@144666.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@144660.4]
  assign regs_114_clock = clock; // @[:@144669.4]
  assign regs_114_reset = io_reset; // @[:@144670.4 RegFile.scala 76:16:@144677.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@144676.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@144680.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@144674.4]
  assign regs_115_clock = clock; // @[:@144683.4]
  assign regs_115_reset = io_reset; // @[:@144684.4 RegFile.scala 76:16:@144691.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@144690.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@144694.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@144688.4]
  assign regs_116_clock = clock; // @[:@144697.4]
  assign regs_116_reset = io_reset; // @[:@144698.4 RegFile.scala 76:16:@144705.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@144704.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@144708.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@144702.4]
  assign regs_117_clock = clock; // @[:@144711.4]
  assign regs_117_reset = io_reset; // @[:@144712.4 RegFile.scala 76:16:@144719.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@144718.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@144722.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@144716.4]
  assign regs_118_clock = clock; // @[:@144725.4]
  assign regs_118_reset = io_reset; // @[:@144726.4 RegFile.scala 76:16:@144733.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@144732.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@144736.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@144730.4]
  assign regs_119_clock = clock; // @[:@144739.4]
  assign regs_119_reset = io_reset; // @[:@144740.4 RegFile.scala 76:16:@144747.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@144746.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@144750.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@144744.4]
  assign regs_120_clock = clock; // @[:@144753.4]
  assign regs_120_reset = io_reset; // @[:@144754.4 RegFile.scala 76:16:@144761.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@144760.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@144764.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@144758.4]
  assign regs_121_clock = clock; // @[:@144767.4]
  assign regs_121_reset = io_reset; // @[:@144768.4 RegFile.scala 76:16:@144775.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@144774.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@144778.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@144772.4]
  assign regs_122_clock = clock; // @[:@144781.4]
  assign regs_122_reset = io_reset; // @[:@144782.4 RegFile.scala 76:16:@144789.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@144788.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@144792.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@144786.4]
  assign regs_123_clock = clock; // @[:@144795.4]
  assign regs_123_reset = io_reset; // @[:@144796.4 RegFile.scala 76:16:@144803.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@144802.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@144806.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@144800.4]
  assign regs_124_clock = clock; // @[:@144809.4]
  assign regs_124_reset = io_reset; // @[:@144810.4 RegFile.scala 76:16:@144817.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@144816.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@144820.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@144814.4]
  assign regs_125_clock = clock; // @[:@144823.4]
  assign regs_125_reset = io_reset; // @[:@144824.4 RegFile.scala 76:16:@144831.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@144830.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@144834.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@144828.4]
  assign regs_126_clock = clock; // @[:@144837.4]
  assign regs_126_reset = io_reset; // @[:@144838.4 RegFile.scala 76:16:@144845.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@144844.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@144848.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@144842.4]
  assign regs_127_clock = clock; // @[:@144851.4]
  assign regs_127_reset = io_reset; // @[:@144852.4 RegFile.scala 76:16:@144859.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@144858.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@144862.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@144856.4]
  assign regs_128_clock = clock; // @[:@144865.4]
  assign regs_128_reset = io_reset; // @[:@144866.4 RegFile.scala 76:16:@144873.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@144872.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@144876.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@144870.4]
  assign regs_129_clock = clock; // @[:@144879.4]
  assign regs_129_reset = io_reset; // @[:@144880.4 RegFile.scala 76:16:@144887.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@144886.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@144890.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@144884.4]
  assign regs_130_clock = clock; // @[:@144893.4]
  assign regs_130_reset = io_reset; // @[:@144894.4 RegFile.scala 76:16:@144901.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@144900.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@144904.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@144898.4]
  assign regs_131_clock = clock; // @[:@144907.4]
  assign regs_131_reset = io_reset; // @[:@144908.4 RegFile.scala 76:16:@144915.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@144914.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@144918.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@144912.4]
  assign regs_132_clock = clock; // @[:@144921.4]
  assign regs_132_reset = io_reset; // @[:@144922.4 RegFile.scala 76:16:@144929.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@144928.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@144932.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@144926.4]
  assign regs_133_clock = clock; // @[:@144935.4]
  assign regs_133_reset = io_reset; // @[:@144936.4 RegFile.scala 76:16:@144943.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@144942.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@144946.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@144940.4]
  assign regs_134_clock = clock; // @[:@144949.4]
  assign regs_134_reset = io_reset; // @[:@144950.4 RegFile.scala 76:16:@144957.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@144956.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@144960.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@144954.4]
  assign regs_135_clock = clock; // @[:@144963.4]
  assign regs_135_reset = io_reset; // @[:@144964.4 RegFile.scala 76:16:@144971.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@144970.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@144974.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@144968.4]
  assign regs_136_clock = clock; // @[:@144977.4]
  assign regs_136_reset = io_reset; // @[:@144978.4 RegFile.scala 76:16:@144985.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@144984.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@144988.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@144982.4]
  assign regs_137_clock = clock; // @[:@144991.4]
  assign regs_137_reset = io_reset; // @[:@144992.4 RegFile.scala 76:16:@144999.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@144998.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@145002.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@144996.4]
  assign regs_138_clock = clock; // @[:@145005.4]
  assign regs_138_reset = io_reset; // @[:@145006.4 RegFile.scala 76:16:@145013.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@145012.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@145016.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@145010.4]
  assign regs_139_clock = clock; // @[:@145019.4]
  assign regs_139_reset = io_reset; // @[:@145020.4 RegFile.scala 76:16:@145027.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@145026.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@145030.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@145024.4]
  assign regs_140_clock = clock; // @[:@145033.4]
  assign regs_140_reset = io_reset; // @[:@145034.4 RegFile.scala 76:16:@145041.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@145040.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@145044.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@145038.4]
  assign regs_141_clock = clock; // @[:@145047.4]
  assign regs_141_reset = io_reset; // @[:@145048.4 RegFile.scala 76:16:@145055.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@145054.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@145058.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@145052.4]
  assign regs_142_clock = clock; // @[:@145061.4]
  assign regs_142_reset = io_reset; // @[:@145062.4 RegFile.scala 76:16:@145069.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@145068.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@145072.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@145066.4]
  assign regs_143_clock = clock; // @[:@145075.4]
  assign regs_143_reset = io_reset; // @[:@145076.4 RegFile.scala 76:16:@145083.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@145082.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@145086.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@145080.4]
  assign regs_144_clock = clock; // @[:@145089.4]
  assign regs_144_reset = io_reset; // @[:@145090.4 RegFile.scala 76:16:@145097.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@145096.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@145100.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@145094.4]
  assign regs_145_clock = clock; // @[:@145103.4]
  assign regs_145_reset = io_reset; // @[:@145104.4 RegFile.scala 76:16:@145111.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@145110.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@145114.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@145108.4]
  assign regs_146_clock = clock; // @[:@145117.4]
  assign regs_146_reset = io_reset; // @[:@145118.4 RegFile.scala 76:16:@145125.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@145124.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@145128.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@145122.4]
  assign regs_147_clock = clock; // @[:@145131.4]
  assign regs_147_reset = io_reset; // @[:@145132.4 RegFile.scala 76:16:@145139.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@145138.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@145142.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@145136.4]
  assign regs_148_clock = clock; // @[:@145145.4]
  assign regs_148_reset = io_reset; // @[:@145146.4 RegFile.scala 76:16:@145153.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@145152.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@145156.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@145150.4]
  assign regs_149_clock = clock; // @[:@145159.4]
  assign regs_149_reset = io_reset; // @[:@145160.4 RegFile.scala 76:16:@145167.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@145166.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@145170.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@145164.4]
  assign regs_150_clock = clock; // @[:@145173.4]
  assign regs_150_reset = io_reset; // @[:@145174.4 RegFile.scala 76:16:@145181.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@145180.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@145184.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@145178.4]
  assign regs_151_clock = clock; // @[:@145187.4]
  assign regs_151_reset = io_reset; // @[:@145188.4 RegFile.scala 76:16:@145195.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@145194.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@145198.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@145192.4]
  assign regs_152_clock = clock; // @[:@145201.4]
  assign regs_152_reset = io_reset; // @[:@145202.4 RegFile.scala 76:16:@145209.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@145208.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@145212.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@145206.4]
  assign regs_153_clock = clock; // @[:@145215.4]
  assign regs_153_reset = io_reset; // @[:@145216.4 RegFile.scala 76:16:@145223.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@145222.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@145226.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@145220.4]
  assign regs_154_clock = clock; // @[:@145229.4]
  assign regs_154_reset = io_reset; // @[:@145230.4 RegFile.scala 76:16:@145237.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@145236.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@145240.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@145234.4]
  assign regs_155_clock = clock; // @[:@145243.4]
  assign regs_155_reset = io_reset; // @[:@145244.4 RegFile.scala 76:16:@145251.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@145250.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@145254.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@145248.4]
  assign regs_156_clock = clock; // @[:@145257.4]
  assign regs_156_reset = io_reset; // @[:@145258.4 RegFile.scala 76:16:@145265.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@145264.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@145268.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@145262.4]
  assign regs_157_clock = clock; // @[:@145271.4]
  assign regs_157_reset = io_reset; // @[:@145272.4 RegFile.scala 76:16:@145279.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@145278.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@145282.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@145276.4]
  assign regs_158_clock = clock; // @[:@145285.4]
  assign regs_158_reset = io_reset; // @[:@145286.4 RegFile.scala 76:16:@145293.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@145292.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@145296.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@145290.4]
  assign regs_159_clock = clock; // @[:@145299.4]
  assign regs_159_reset = io_reset; // @[:@145300.4 RegFile.scala 76:16:@145307.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@145306.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@145310.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@145304.4]
  assign regs_160_clock = clock; // @[:@145313.4]
  assign regs_160_reset = io_reset; // @[:@145314.4 RegFile.scala 76:16:@145321.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@145320.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@145324.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@145318.4]
  assign regs_161_clock = clock; // @[:@145327.4]
  assign regs_161_reset = io_reset; // @[:@145328.4 RegFile.scala 76:16:@145335.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@145334.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@145338.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@145332.4]
  assign regs_162_clock = clock; // @[:@145341.4]
  assign regs_162_reset = io_reset; // @[:@145342.4 RegFile.scala 76:16:@145349.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@145348.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@145352.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@145346.4]
  assign regs_163_clock = clock; // @[:@145355.4]
  assign regs_163_reset = io_reset; // @[:@145356.4 RegFile.scala 76:16:@145363.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@145362.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@145366.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@145360.4]
  assign regs_164_clock = clock; // @[:@145369.4]
  assign regs_164_reset = io_reset; // @[:@145370.4 RegFile.scala 76:16:@145377.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@145376.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@145380.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@145374.4]
  assign regs_165_clock = clock; // @[:@145383.4]
  assign regs_165_reset = io_reset; // @[:@145384.4 RegFile.scala 76:16:@145391.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@145390.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@145394.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@145388.4]
  assign regs_166_clock = clock; // @[:@145397.4]
  assign regs_166_reset = io_reset; // @[:@145398.4 RegFile.scala 76:16:@145405.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@145404.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@145408.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@145402.4]
  assign regs_167_clock = clock; // @[:@145411.4]
  assign regs_167_reset = io_reset; // @[:@145412.4 RegFile.scala 76:16:@145419.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@145418.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@145422.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@145416.4]
  assign regs_168_clock = clock; // @[:@145425.4]
  assign regs_168_reset = io_reset; // @[:@145426.4 RegFile.scala 76:16:@145433.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@145432.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@145436.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@145430.4]
  assign regs_169_clock = clock; // @[:@145439.4]
  assign regs_169_reset = io_reset; // @[:@145440.4 RegFile.scala 76:16:@145447.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@145446.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@145450.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@145444.4]
  assign regs_170_clock = clock; // @[:@145453.4]
  assign regs_170_reset = io_reset; // @[:@145454.4 RegFile.scala 76:16:@145461.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@145460.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@145464.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@145458.4]
  assign regs_171_clock = clock; // @[:@145467.4]
  assign regs_171_reset = io_reset; // @[:@145468.4 RegFile.scala 76:16:@145475.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@145474.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@145478.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@145472.4]
  assign regs_172_clock = clock; // @[:@145481.4]
  assign regs_172_reset = io_reset; // @[:@145482.4 RegFile.scala 76:16:@145489.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@145488.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@145492.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@145486.4]
  assign regs_173_clock = clock; // @[:@145495.4]
  assign regs_173_reset = io_reset; // @[:@145496.4 RegFile.scala 76:16:@145503.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@145502.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@145506.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@145500.4]
  assign regs_174_clock = clock; // @[:@145509.4]
  assign regs_174_reset = io_reset; // @[:@145510.4 RegFile.scala 76:16:@145517.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@145516.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@145520.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@145514.4]
  assign regs_175_clock = clock; // @[:@145523.4]
  assign regs_175_reset = io_reset; // @[:@145524.4 RegFile.scala 76:16:@145531.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@145530.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@145534.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@145528.4]
  assign regs_176_clock = clock; // @[:@145537.4]
  assign regs_176_reset = io_reset; // @[:@145538.4 RegFile.scala 76:16:@145545.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@145544.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@145548.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@145542.4]
  assign regs_177_clock = clock; // @[:@145551.4]
  assign regs_177_reset = io_reset; // @[:@145552.4 RegFile.scala 76:16:@145559.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@145558.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@145562.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@145556.4]
  assign regs_178_clock = clock; // @[:@145565.4]
  assign regs_178_reset = io_reset; // @[:@145566.4 RegFile.scala 76:16:@145573.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@145572.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@145576.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@145570.4]
  assign regs_179_clock = clock; // @[:@145579.4]
  assign regs_179_reset = io_reset; // @[:@145580.4 RegFile.scala 76:16:@145587.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@145586.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@145590.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@145584.4]
  assign regs_180_clock = clock; // @[:@145593.4]
  assign regs_180_reset = io_reset; // @[:@145594.4 RegFile.scala 76:16:@145601.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@145600.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@145604.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@145598.4]
  assign regs_181_clock = clock; // @[:@145607.4]
  assign regs_181_reset = io_reset; // @[:@145608.4 RegFile.scala 76:16:@145615.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@145614.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@145618.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@145612.4]
  assign regs_182_clock = clock; // @[:@145621.4]
  assign regs_182_reset = io_reset; // @[:@145622.4 RegFile.scala 76:16:@145629.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@145628.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@145632.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@145626.4]
  assign regs_183_clock = clock; // @[:@145635.4]
  assign regs_183_reset = io_reset; // @[:@145636.4 RegFile.scala 76:16:@145643.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@145642.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@145646.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@145640.4]
  assign regs_184_clock = clock; // @[:@145649.4]
  assign regs_184_reset = io_reset; // @[:@145650.4 RegFile.scala 76:16:@145657.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@145656.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@145660.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@145654.4]
  assign regs_185_clock = clock; // @[:@145663.4]
  assign regs_185_reset = io_reset; // @[:@145664.4 RegFile.scala 76:16:@145671.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@145670.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@145674.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@145668.4]
  assign regs_186_clock = clock; // @[:@145677.4]
  assign regs_186_reset = io_reset; // @[:@145678.4 RegFile.scala 76:16:@145685.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@145684.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@145688.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@145682.4]
  assign regs_187_clock = clock; // @[:@145691.4]
  assign regs_187_reset = io_reset; // @[:@145692.4 RegFile.scala 76:16:@145699.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@145698.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@145702.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@145696.4]
  assign regs_188_clock = clock; // @[:@145705.4]
  assign regs_188_reset = io_reset; // @[:@145706.4 RegFile.scala 76:16:@145713.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@145712.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@145716.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@145710.4]
  assign regs_189_clock = clock; // @[:@145719.4]
  assign regs_189_reset = io_reset; // @[:@145720.4 RegFile.scala 76:16:@145727.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@145726.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@145730.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@145724.4]
  assign regs_190_clock = clock; // @[:@145733.4]
  assign regs_190_reset = io_reset; // @[:@145734.4 RegFile.scala 76:16:@145741.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@145740.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@145744.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@145738.4]
  assign regs_191_clock = clock; // @[:@145747.4]
  assign regs_191_reset = io_reset; // @[:@145748.4 RegFile.scala 76:16:@145755.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@145754.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@145758.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@145752.4]
  assign regs_192_clock = clock; // @[:@145761.4]
  assign regs_192_reset = io_reset; // @[:@145762.4 RegFile.scala 76:16:@145769.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@145768.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@145772.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@145766.4]
  assign regs_193_clock = clock; // @[:@145775.4]
  assign regs_193_reset = io_reset; // @[:@145776.4 RegFile.scala 76:16:@145783.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@145782.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@145786.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@145780.4]
  assign regs_194_clock = clock; // @[:@145789.4]
  assign regs_194_reset = io_reset; // @[:@145790.4 RegFile.scala 76:16:@145797.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@145796.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@145800.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@145794.4]
  assign regs_195_clock = clock; // @[:@145803.4]
  assign regs_195_reset = io_reset; // @[:@145804.4 RegFile.scala 76:16:@145811.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@145810.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@145814.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@145808.4]
  assign regs_196_clock = clock; // @[:@145817.4]
  assign regs_196_reset = io_reset; // @[:@145818.4 RegFile.scala 76:16:@145825.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@145824.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@145828.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@145822.4]
  assign regs_197_clock = clock; // @[:@145831.4]
  assign regs_197_reset = io_reset; // @[:@145832.4 RegFile.scala 76:16:@145839.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@145838.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@145842.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@145836.4]
  assign regs_198_clock = clock; // @[:@145845.4]
  assign regs_198_reset = io_reset; // @[:@145846.4 RegFile.scala 76:16:@145853.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@145852.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@145856.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@145850.4]
  assign regs_199_clock = clock; // @[:@145859.4]
  assign regs_199_reset = io_reset; // @[:@145860.4 RegFile.scala 76:16:@145867.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@145866.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@145870.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@145864.4]
  assign regs_200_clock = clock; // @[:@145873.4]
  assign regs_200_reset = io_reset; // @[:@145874.4 RegFile.scala 76:16:@145881.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@145880.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@145884.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@145878.4]
  assign regs_201_clock = clock; // @[:@145887.4]
  assign regs_201_reset = io_reset; // @[:@145888.4 RegFile.scala 76:16:@145895.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@145894.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@145898.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@145892.4]
  assign regs_202_clock = clock; // @[:@145901.4]
  assign regs_202_reset = io_reset; // @[:@145902.4 RegFile.scala 76:16:@145909.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@145908.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@145912.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@145906.4]
  assign regs_203_clock = clock; // @[:@145915.4]
  assign regs_203_reset = io_reset; // @[:@145916.4 RegFile.scala 76:16:@145923.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@145922.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@145926.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@145920.4]
  assign regs_204_clock = clock; // @[:@145929.4]
  assign regs_204_reset = io_reset; // @[:@145930.4 RegFile.scala 76:16:@145937.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@145936.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@145940.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@145934.4]
  assign regs_205_clock = clock; // @[:@145943.4]
  assign regs_205_reset = io_reset; // @[:@145944.4 RegFile.scala 76:16:@145951.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@145950.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@145954.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@145948.4]
  assign regs_206_clock = clock; // @[:@145957.4]
  assign regs_206_reset = io_reset; // @[:@145958.4 RegFile.scala 76:16:@145965.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@145964.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@145968.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@145962.4]
  assign regs_207_clock = clock; // @[:@145971.4]
  assign regs_207_reset = io_reset; // @[:@145972.4 RegFile.scala 76:16:@145979.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@145978.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@145982.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@145976.4]
  assign regs_208_clock = clock; // @[:@145985.4]
  assign regs_208_reset = io_reset; // @[:@145986.4 RegFile.scala 76:16:@145993.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@145992.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@145996.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@145990.4]
  assign regs_209_clock = clock; // @[:@145999.4]
  assign regs_209_reset = io_reset; // @[:@146000.4 RegFile.scala 76:16:@146007.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@146006.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@146010.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@146004.4]
  assign regs_210_clock = clock; // @[:@146013.4]
  assign regs_210_reset = io_reset; // @[:@146014.4 RegFile.scala 76:16:@146021.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@146020.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@146024.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@146018.4]
  assign regs_211_clock = clock; // @[:@146027.4]
  assign regs_211_reset = io_reset; // @[:@146028.4 RegFile.scala 76:16:@146035.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@146034.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@146038.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@146032.4]
  assign regs_212_clock = clock; // @[:@146041.4]
  assign regs_212_reset = io_reset; // @[:@146042.4 RegFile.scala 76:16:@146049.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@146048.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@146052.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@146046.4]
  assign regs_213_clock = clock; // @[:@146055.4]
  assign regs_213_reset = io_reset; // @[:@146056.4 RegFile.scala 76:16:@146063.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@146062.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@146066.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@146060.4]
  assign regs_214_clock = clock; // @[:@146069.4]
  assign regs_214_reset = io_reset; // @[:@146070.4 RegFile.scala 76:16:@146077.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@146076.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@146080.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@146074.4]
  assign regs_215_clock = clock; // @[:@146083.4]
  assign regs_215_reset = io_reset; // @[:@146084.4 RegFile.scala 76:16:@146091.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@146090.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@146094.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@146088.4]
  assign regs_216_clock = clock; // @[:@146097.4]
  assign regs_216_reset = io_reset; // @[:@146098.4 RegFile.scala 76:16:@146105.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@146104.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@146108.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@146102.4]
  assign regs_217_clock = clock; // @[:@146111.4]
  assign regs_217_reset = io_reset; // @[:@146112.4 RegFile.scala 76:16:@146119.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@146118.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@146122.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@146116.4]
  assign regs_218_clock = clock; // @[:@146125.4]
  assign regs_218_reset = io_reset; // @[:@146126.4 RegFile.scala 76:16:@146133.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@146132.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@146136.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@146130.4]
  assign regs_219_clock = clock; // @[:@146139.4]
  assign regs_219_reset = io_reset; // @[:@146140.4 RegFile.scala 76:16:@146147.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@146146.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@146150.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@146144.4]
  assign regs_220_clock = clock; // @[:@146153.4]
  assign regs_220_reset = io_reset; // @[:@146154.4 RegFile.scala 76:16:@146161.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@146160.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@146164.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@146158.4]
  assign regs_221_clock = clock; // @[:@146167.4]
  assign regs_221_reset = io_reset; // @[:@146168.4 RegFile.scala 76:16:@146175.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@146174.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@146178.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@146172.4]
  assign regs_222_clock = clock; // @[:@146181.4]
  assign regs_222_reset = io_reset; // @[:@146182.4 RegFile.scala 76:16:@146189.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@146188.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@146192.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@146186.4]
  assign regs_223_clock = clock; // @[:@146195.4]
  assign regs_223_reset = io_reset; // @[:@146196.4 RegFile.scala 76:16:@146203.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@146202.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@146206.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@146200.4]
  assign regs_224_clock = clock; // @[:@146209.4]
  assign regs_224_reset = io_reset; // @[:@146210.4 RegFile.scala 76:16:@146217.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@146216.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@146220.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@146214.4]
  assign regs_225_clock = clock; // @[:@146223.4]
  assign regs_225_reset = io_reset; // @[:@146224.4 RegFile.scala 76:16:@146231.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@146230.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@146234.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@146228.4]
  assign regs_226_clock = clock; // @[:@146237.4]
  assign regs_226_reset = io_reset; // @[:@146238.4 RegFile.scala 76:16:@146245.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@146244.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@146248.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@146242.4]
  assign regs_227_clock = clock; // @[:@146251.4]
  assign regs_227_reset = io_reset; // @[:@146252.4 RegFile.scala 76:16:@146259.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@146258.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@146262.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@146256.4]
  assign regs_228_clock = clock; // @[:@146265.4]
  assign regs_228_reset = io_reset; // @[:@146266.4 RegFile.scala 76:16:@146273.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@146272.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@146276.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@146270.4]
  assign regs_229_clock = clock; // @[:@146279.4]
  assign regs_229_reset = io_reset; // @[:@146280.4 RegFile.scala 76:16:@146287.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@146286.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@146290.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@146284.4]
  assign regs_230_clock = clock; // @[:@146293.4]
  assign regs_230_reset = io_reset; // @[:@146294.4 RegFile.scala 76:16:@146301.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@146300.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@146304.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@146298.4]
  assign regs_231_clock = clock; // @[:@146307.4]
  assign regs_231_reset = io_reset; // @[:@146308.4 RegFile.scala 76:16:@146315.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@146314.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@146318.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@146312.4]
  assign regs_232_clock = clock; // @[:@146321.4]
  assign regs_232_reset = io_reset; // @[:@146322.4 RegFile.scala 76:16:@146329.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@146328.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@146332.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@146326.4]
  assign regs_233_clock = clock; // @[:@146335.4]
  assign regs_233_reset = io_reset; // @[:@146336.4 RegFile.scala 76:16:@146343.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@146342.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@146346.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@146340.4]
  assign regs_234_clock = clock; // @[:@146349.4]
  assign regs_234_reset = io_reset; // @[:@146350.4 RegFile.scala 76:16:@146357.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@146356.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@146360.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@146354.4]
  assign regs_235_clock = clock; // @[:@146363.4]
  assign regs_235_reset = io_reset; // @[:@146364.4 RegFile.scala 76:16:@146371.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@146370.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@146374.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@146368.4]
  assign regs_236_clock = clock; // @[:@146377.4]
  assign regs_236_reset = io_reset; // @[:@146378.4 RegFile.scala 76:16:@146385.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@146384.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@146388.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@146382.4]
  assign regs_237_clock = clock; // @[:@146391.4]
  assign regs_237_reset = io_reset; // @[:@146392.4 RegFile.scala 76:16:@146399.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@146398.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@146402.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@146396.4]
  assign regs_238_clock = clock; // @[:@146405.4]
  assign regs_238_reset = io_reset; // @[:@146406.4 RegFile.scala 76:16:@146413.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@146412.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@146416.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@146410.4]
  assign regs_239_clock = clock; // @[:@146419.4]
  assign regs_239_reset = io_reset; // @[:@146420.4 RegFile.scala 76:16:@146427.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@146426.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@146430.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@146424.4]
  assign regs_240_clock = clock; // @[:@146433.4]
  assign regs_240_reset = io_reset; // @[:@146434.4 RegFile.scala 76:16:@146441.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@146440.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@146444.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@146438.4]
  assign regs_241_clock = clock; // @[:@146447.4]
  assign regs_241_reset = io_reset; // @[:@146448.4 RegFile.scala 76:16:@146455.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@146454.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@146458.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@146452.4]
  assign regs_242_clock = clock; // @[:@146461.4]
  assign regs_242_reset = io_reset; // @[:@146462.4 RegFile.scala 76:16:@146469.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@146468.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@146472.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@146466.4]
  assign regs_243_clock = clock; // @[:@146475.4]
  assign regs_243_reset = io_reset; // @[:@146476.4 RegFile.scala 76:16:@146483.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@146482.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@146486.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@146480.4]
  assign regs_244_clock = clock; // @[:@146489.4]
  assign regs_244_reset = io_reset; // @[:@146490.4 RegFile.scala 76:16:@146497.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@146496.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@146500.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@146494.4]
  assign regs_245_clock = clock; // @[:@146503.4]
  assign regs_245_reset = io_reset; // @[:@146504.4 RegFile.scala 76:16:@146511.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@146510.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@146514.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@146508.4]
  assign regs_246_clock = clock; // @[:@146517.4]
  assign regs_246_reset = io_reset; // @[:@146518.4 RegFile.scala 76:16:@146525.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@146524.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@146528.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@146522.4]
  assign regs_247_clock = clock; // @[:@146531.4]
  assign regs_247_reset = io_reset; // @[:@146532.4 RegFile.scala 76:16:@146539.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@146538.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@146542.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@146536.4]
  assign regs_248_clock = clock; // @[:@146545.4]
  assign regs_248_reset = io_reset; // @[:@146546.4 RegFile.scala 76:16:@146553.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@146552.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@146556.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@146550.4]
  assign regs_249_clock = clock; // @[:@146559.4]
  assign regs_249_reset = io_reset; // @[:@146560.4 RegFile.scala 76:16:@146567.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@146566.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@146570.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@146564.4]
  assign regs_250_clock = clock; // @[:@146573.4]
  assign regs_250_reset = io_reset; // @[:@146574.4 RegFile.scala 76:16:@146581.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@146580.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@146584.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@146578.4]
  assign regs_251_clock = clock; // @[:@146587.4]
  assign regs_251_reset = io_reset; // @[:@146588.4 RegFile.scala 76:16:@146595.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@146594.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@146598.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@146592.4]
  assign regs_252_clock = clock; // @[:@146601.4]
  assign regs_252_reset = io_reset; // @[:@146602.4 RegFile.scala 76:16:@146609.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@146608.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@146612.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@146606.4]
  assign regs_253_clock = clock; // @[:@146615.4]
  assign regs_253_reset = io_reset; // @[:@146616.4 RegFile.scala 76:16:@146623.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@146622.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@146626.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@146620.4]
  assign regs_254_clock = clock; // @[:@146629.4]
  assign regs_254_reset = io_reset; // @[:@146630.4 RegFile.scala 76:16:@146637.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@146636.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@146640.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@146634.4]
  assign regs_255_clock = clock; // @[:@146643.4]
  assign regs_255_reset = io_reset; // @[:@146644.4 RegFile.scala 76:16:@146651.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@146650.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@146654.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@146648.4]
  assign regs_256_clock = clock; // @[:@146657.4]
  assign regs_256_reset = io_reset; // @[:@146658.4 RegFile.scala 76:16:@146665.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@146664.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@146668.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@146662.4]
  assign regs_257_clock = clock; // @[:@146671.4]
  assign regs_257_reset = io_reset; // @[:@146672.4 RegFile.scala 76:16:@146679.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@146678.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@146682.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@146676.4]
  assign regs_258_clock = clock; // @[:@146685.4]
  assign regs_258_reset = io_reset; // @[:@146686.4 RegFile.scala 76:16:@146693.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@146692.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@146696.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@146690.4]
  assign regs_259_clock = clock; // @[:@146699.4]
  assign regs_259_reset = io_reset; // @[:@146700.4 RegFile.scala 76:16:@146707.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@146706.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@146710.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@146704.4]
  assign regs_260_clock = clock; // @[:@146713.4]
  assign regs_260_reset = io_reset; // @[:@146714.4 RegFile.scala 76:16:@146721.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@146720.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@146724.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@146718.4]
  assign regs_261_clock = clock; // @[:@146727.4]
  assign regs_261_reset = io_reset; // @[:@146728.4 RegFile.scala 76:16:@146735.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@146734.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@146738.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@146732.4]
  assign regs_262_clock = clock; // @[:@146741.4]
  assign regs_262_reset = io_reset; // @[:@146742.4 RegFile.scala 76:16:@146749.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@146748.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@146752.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@146746.4]
  assign regs_263_clock = clock; // @[:@146755.4]
  assign regs_263_reset = io_reset; // @[:@146756.4 RegFile.scala 76:16:@146763.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@146762.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@146766.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@146760.4]
  assign regs_264_clock = clock; // @[:@146769.4]
  assign regs_264_reset = io_reset; // @[:@146770.4 RegFile.scala 76:16:@146777.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@146776.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@146780.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@146774.4]
  assign regs_265_clock = clock; // @[:@146783.4]
  assign regs_265_reset = io_reset; // @[:@146784.4 RegFile.scala 76:16:@146791.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@146790.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@146794.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@146788.4]
  assign regs_266_clock = clock; // @[:@146797.4]
  assign regs_266_reset = io_reset; // @[:@146798.4 RegFile.scala 76:16:@146805.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@146804.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@146808.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@146802.4]
  assign regs_267_clock = clock; // @[:@146811.4]
  assign regs_267_reset = io_reset; // @[:@146812.4 RegFile.scala 76:16:@146819.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@146818.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@146822.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@146816.4]
  assign regs_268_clock = clock; // @[:@146825.4]
  assign regs_268_reset = io_reset; // @[:@146826.4 RegFile.scala 76:16:@146833.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@146832.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@146836.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@146830.4]
  assign regs_269_clock = clock; // @[:@146839.4]
  assign regs_269_reset = io_reset; // @[:@146840.4 RegFile.scala 76:16:@146847.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@146846.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@146850.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@146844.4]
  assign regs_270_clock = clock; // @[:@146853.4]
  assign regs_270_reset = io_reset; // @[:@146854.4 RegFile.scala 76:16:@146861.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@146860.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@146864.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@146858.4]
  assign regs_271_clock = clock; // @[:@146867.4]
  assign regs_271_reset = io_reset; // @[:@146868.4 RegFile.scala 76:16:@146875.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@146874.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@146878.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@146872.4]
  assign regs_272_clock = clock; // @[:@146881.4]
  assign regs_272_reset = io_reset; // @[:@146882.4 RegFile.scala 76:16:@146889.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@146888.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@146892.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@146886.4]
  assign regs_273_clock = clock; // @[:@146895.4]
  assign regs_273_reset = io_reset; // @[:@146896.4 RegFile.scala 76:16:@146903.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@146902.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@146906.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@146900.4]
  assign regs_274_clock = clock; // @[:@146909.4]
  assign regs_274_reset = io_reset; // @[:@146910.4 RegFile.scala 76:16:@146917.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@146916.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@146920.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@146914.4]
  assign regs_275_clock = clock; // @[:@146923.4]
  assign regs_275_reset = io_reset; // @[:@146924.4 RegFile.scala 76:16:@146931.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@146930.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@146934.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@146928.4]
  assign regs_276_clock = clock; // @[:@146937.4]
  assign regs_276_reset = io_reset; // @[:@146938.4 RegFile.scala 76:16:@146945.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@146944.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@146948.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@146942.4]
  assign regs_277_clock = clock; // @[:@146951.4]
  assign regs_277_reset = io_reset; // @[:@146952.4 RegFile.scala 76:16:@146959.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@146958.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@146962.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@146956.4]
  assign regs_278_clock = clock; // @[:@146965.4]
  assign regs_278_reset = io_reset; // @[:@146966.4 RegFile.scala 76:16:@146973.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@146972.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@146976.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@146970.4]
  assign regs_279_clock = clock; // @[:@146979.4]
  assign regs_279_reset = io_reset; // @[:@146980.4 RegFile.scala 76:16:@146987.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@146986.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@146990.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@146984.4]
  assign regs_280_clock = clock; // @[:@146993.4]
  assign regs_280_reset = io_reset; // @[:@146994.4 RegFile.scala 76:16:@147001.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@147000.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@147004.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@146998.4]
  assign regs_281_clock = clock; // @[:@147007.4]
  assign regs_281_reset = io_reset; // @[:@147008.4 RegFile.scala 76:16:@147015.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@147014.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@147018.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@147012.4]
  assign regs_282_clock = clock; // @[:@147021.4]
  assign regs_282_reset = io_reset; // @[:@147022.4 RegFile.scala 76:16:@147029.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@147028.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@147032.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@147026.4]
  assign regs_283_clock = clock; // @[:@147035.4]
  assign regs_283_reset = io_reset; // @[:@147036.4 RegFile.scala 76:16:@147043.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@147042.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@147046.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@147040.4]
  assign regs_284_clock = clock; // @[:@147049.4]
  assign regs_284_reset = io_reset; // @[:@147050.4 RegFile.scala 76:16:@147057.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@147056.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@147060.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@147054.4]
  assign regs_285_clock = clock; // @[:@147063.4]
  assign regs_285_reset = io_reset; // @[:@147064.4 RegFile.scala 76:16:@147071.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@147070.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@147074.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@147068.4]
  assign regs_286_clock = clock; // @[:@147077.4]
  assign regs_286_reset = io_reset; // @[:@147078.4 RegFile.scala 76:16:@147085.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@147084.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@147088.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@147082.4]
  assign regs_287_clock = clock; // @[:@147091.4]
  assign regs_287_reset = io_reset; // @[:@147092.4 RegFile.scala 76:16:@147099.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@147098.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@147102.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@147096.4]
  assign regs_288_clock = clock; // @[:@147105.4]
  assign regs_288_reset = io_reset; // @[:@147106.4 RegFile.scala 76:16:@147113.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@147112.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@147116.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@147110.4]
  assign regs_289_clock = clock; // @[:@147119.4]
  assign regs_289_reset = io_reset; // @[:@147120.4 RegFile.scala 76:16:@147127.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@147126.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@147130.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@147124.4]
  assign regs_290_clock = clock; // @[:@147133.4]
  assign regs_290_reset = io_reset; // @[:@147134.4 RegFile.scala 76:16:@147141.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@147140.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@147144.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@147138.4]
  assign regs_291_clock = clock; // @[:@147147.4]
  assign regs_291_reset = io_reset; // @[:@147148.4 RegFile.scala 76:16:@147155.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@147154.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@147158.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@147152.4]
  assign regs_292_clock = clock; // @[:@147161.4]
  assign regs_292_reset = io_reset; // @[:@147162.4 RegFile.scala 76:16:@147169.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@147168.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@147172.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@147166.4]
  assign regs_293_clock = clock; // @[:@147175.4]
  assign regs_293_reset = io_reset; // @[:@147176.4 RegFile.scala 76:16:@147183.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@147182.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@147186.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@147180.4]
  assign regs_294_clock = clock; // @[:@147189.4]
  assign regs_294_reset = io_reset; // @[:@147190.4 RegFile.scala 76:16:@147197.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@147196.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@147200.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@147194.4]
  assign regs_295_clock = clock; // @[:@147203.4]
  assign regs_295_reset = io_reset; // @[:@147204.4 RegFile.scala 76:16:@147211.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@147210.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@147214.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@147208.4]
  assign regs_296_clock = clock; // @[:@147217.4]
  assign regs_296_reset = io_reset; // @[:@147218.4 RegFile.scala 76:16:@147225.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@147224.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@147228.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@147222.4]
  assign regs_297_clock = clock; // @[:@147231.4]
  assign regs_297_reset = io_reset; // @[:@147232.4 RegFile.scala 76:16:@147239.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@147238.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@147242.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@147236.4]
  assign regs_298_clock = clock; // @[:@147245.4]
  assign regs_298_reset = io_reset; // @[:@147246.4 RegFile.scala 76:16:@147253.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@147252.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@147256.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@147250.4]
  assign regs_299_clock = clock; // @[:@147259.4]
  assign regs_299_reset = io_reset; // @[:@147260.4 RegFile.scala 76:16:@147267.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@147266.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@147270.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@147264.4]
  assign regs_300_clock = clock; // @[:@147273.4]
  assign regs_300_reset = io_reset; // @[:@147274.4 RegFile.scala 76:16:@147281.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@147280.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@147284.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@147278.4]
  assign regs_301_clock = clock; // @[:@147287.4]
  assign regs_301_reset = io_reset; // @[:@147288.4 RegFile.scala 76:16:@147295.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@147294.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@147298.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@147292.4]
  assign regs_302_clock = clock; // @[:@147301.4]
  assign regs_302_reset = io_reset; // @[:@147302.4 RegFile.scala 76:16:@147309.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@147308.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@147312.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@147306.4]
  assign regs_303_clock = clock; // @[:@147315.4]
  assign regs_303_reset = io_reset; // @[:@147316.4 RegFile.scala 76:16:@147323.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@147322.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@147326.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@147320.4]
  assign regs_304_clock = clock; // @[:@147329.4]
  assign regs_304_reset = io_reset; // @[:@147330.4 RegFile.scala 76:16:@147337.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@147336.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@147340.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@147334.4]
  assign regs_305_clock = clock; // @[:@147343.4]
  assign regs_305_reset = io_reset; // @[:@147344.4 RegFile.scala 76:16:@147351.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@147350.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@147354.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@147348.4]
  assign regs_306_clock = clock; // @[:@147357.4]
  assign regs_306_reset = io_reset; // @[:@147358.4 RegFile.scala 76:16:@147365.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@147364.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@147368.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@147362.4]
  assign regs_307_clock = clock; // @[:@147371.4]
  assign regs_307_reset = io_reset; // @[:@147372.4 RegFile.scala 76:16:@147379.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@147378.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@147382.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@147376.4]
  assign regs_308_clock = clock; // @[:@147385.4]
  assign regs_308_reset = io_reset; // @[:@147386.4 RegFile.scala 76:16:@147393.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@147392.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@147396.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@147390.4]
  assign regs_309_clock = clock; // @[:@147399.4]
  assign regs_309_reset = io_reset; // @[:@147400.4 RegFile.scala 76:16:@147407.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@147406.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@147410.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@147404.4]
  assign regs_310_clock = clock; // @[:@147413.4]
  assign regs_310_reset = io_reset; // @[:@147414.4 RegFile.scala 76:16:@147421.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@147420.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@147424.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@147418.4]
  assign regs_311_clock = clock; // @[:@147427.4]
  assign regs_311_reset = io_reset; // @[:@147428.4 RegFile.scala 76:16:@147435.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@147434.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@147438.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@147432.4]
  assign regs_312_clock = clock; // @[:@147441.4]
  assign regs_312_reset = io_reset; // @[:@147442.4 RegFile.scala 76:16:@147449.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@147448.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@147452.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@147446.4]
  assign regs_313_clock = clock; // @[:@147455.4]
  assign regs_313_reset = io_reset; // @[:@147456.4 RegFile.scala 76:16:@147463.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@147462.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@147466.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@147460.4]
  assign regs_314_clock = clock; // @[:@147469.4]
  assign regs_314_reset = io_reset; // @[:@147470.4 RegFile.scala 76:16:@147477.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@147476.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@147480.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@147474.4]
  assign regs_315_clock = clock; // @[:@147483.4]
  assign regs_315_reset = io_reset; // @[:@147484.4 RegFile.scala 76:16:@147491.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@147490.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@147494.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@147488.4]
  assign regs_316_clock = clock; // @[:@147497.4]
  assign regs_316_reset = io_reset; // @[:@147498.4 RegFile.scala 76:16:@147505.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@147504.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@147508.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@147502.4]
  assign regs_317_clock = clock; // @[:@147511.4]
  assign regs_317_reset = io_reset; // @[:@147512.4 RegFile.scala 76:16:@147519.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@147518.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@147522.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@147516.4]
  assign regs_318_clock = clock; // @[:@147525.4]
  assign regs_318_reset = io_reset; // @[:@147526.4 RegFile.scala 76:16:@147533.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@147532.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@147536.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@147530.4]
  assign regs_319_clock = clock; // @[:@147539.4]
  assign regs_319_reset = io_reset; // @[:@147540.4 RegFile.scala 76:16:@147547.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@147546.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@147550.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@147544.4]
  assign regs_320_clock = clock; // @[:@147553.4]
  assign regs_320_reset = io_reset; // @[:@147554.4 RegFile.scala 76:16:@147561.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@147560.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@147564.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@147558.4]
  assign regs_321_clock = clock; // @[:@147567.4]
  assign regs_321_reset = io_reset; // @[:@147568.4 RegFile.scala 76:16:@147575.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@147574.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@147578.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@147572.4]
  assign regs_322_clock = clock; // @[:@147581.4]
  assign regs_322_reset = io_reset; // @[:@147582.4 RegFile.scala 76:16:@147589.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@147588.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@147592.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@147586.4]
  assign regs_323_clock = clock; // @[:@147595.4]
  assign regs_323_reset = io_reset; // @[:@147596.4 RegFile.scala 76:16:@147603.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@147602.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@147606.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@147600.4]
  assign regs_324_clock = clock; // @[:@147609.4]
  assign regs_324_reset = io_reset; // @[:@147610.4 RegFile.scala 76:16:@147617.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@147616.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@147620.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@147614.4]
  assign regs_325_clock = clock; // @[:@147623.4]
  assign regs_325_reset = io_reset; // @[:@147624.4 RegFile.scala 76:16:@147631.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@147630.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@147634.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@147628.4]
  assign regs_326_clock = clock; // @[:@147637.4]
  assign regs_326_reset = io_reset; // @[:@147638.4 RegFile.scala 76:16:@147645.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@147644.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@147648.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@147642.4]
  assign regs_327_clock = clock; // @[:@147651.4]
  assign regs_327_reset = io_reset; // @[:@147652.4 RegFile.scala 76:16:@147659.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@147658.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@147662.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@147656.4]
  assign regs_328_clock = clock; // @[:@147665.4]
  assign regs_328_reset = io_reset; // @[:@147666.4 RegFile.scala 76:16:@147673.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@147672.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@147676.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@147670.4]
  assign regs_329_clock = clock; // @[:@147679.4]
  assign regs_329_reset = io_reset; // @[:@147680.4 RegFile.scala 76:16:@147687.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@147686.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@147690.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@147684.4]
  assign regs_330_clock = clock; // @[:@147693.4]
  assign regs_330_reset = io_reset; // @[:@147694.4 RegFile.scala 76:16:@147701.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@147700.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@147704.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@147698.4]
  assign regs_331_clock = clock; // @[:@147707.4]
  assign regs_331_reset = io_reset; // @[:@147708.4 RegFile.scala 76:16:@147715.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@147714.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@147718.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@147712.4]
  assign regs_332_clock = clock; // @[:@147721.4]
  assign regs_332_reset = io_reset; // @[:@147722.4 RegFile.scala 76:16:@147729.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@147728.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@147732.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@147726.4]
  assign regs_333_clock = clock; // @[:@147735.4]
  assign regs_333_reset = io_reset; // @[:@147736.4 RegFile.scala 76:16:@147743.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@147742.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@147746.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@147740.4]
  assign regs_334_clock = clock; // @[:@147749.4]
  assign regs_334_reset = io_reset; // @[:@147750.4 RegFile.scala 76:16:@147757.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@147756.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@147760.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@147754.4]
  assign regs_335_clock = clock; // @[:@147763.4]
  assign regs_335_reset = io_reset; // @[:@147764.4 RegFile.scala 76:16:@147771.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@147770.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@147774.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@147768.4]
  assign regs_336_clock = clock; // @[:@147777.4]
  assign regs_336_reset = io_reset; // @[:@147778.4 RegFile.scala 76:16:@147785.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@147784.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@147788.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@147782.4]
  assign regs_337_clock = clock; // @[:@147791.4]
  assign regs_337_reset = io_reset; // @[:@147792.4 RegFile.scala 76:16:@147799.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@147798.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@147802.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@147796.4]
  assign regs_338_clock = clock; // @[:@147805.4]
  assign regs_338_reset = io_reset; // @[:@147806.4 RegFile.scala 76:16:@147813.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@147812.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@147816.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@147810.4]
  assign regs_339_clock = clock; // @[:@147819.4]
  assign regs_339_reset = io_reset; // @[:@147820.4 RegFile.scala 76:16:@147827.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@147826.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@147830.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@147824.4]
  assign regs_340_clock = clock; // @[:@147833.4]
  assign regs_340_reset = io_reset; // @[:@147834.4 RegFile.scala 76:16:@147841.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@147840.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@147844.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@147838.4]
  assign regs_341_clock = clock; // @[:@147847.4]
  assign regs_341_reset = io_reset; // @[:@147848.4 RegFile.scala 76:16:@147855.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@147854.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@147858.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@147852.4]
  assign regs_342_clock = clock; // @[:@147861.4]
  assign regs_342_reset = io_reset; // @[:@147862.4 RegFile.scala 76:16:@147869.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@147868.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@147872.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@147866.4]
  assign regs_343_clock = clock; // @[:@147875.4]
  assign regs_343_reset = io_reset; // @[:@147876.4 RegFile.scala 76:16:@147883.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@147882.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@147886.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@147880.4]
  assign regs_344_clock = clock; // @[:@147889.4]
  assign regs_344_reset = io_reset; // @[:@147890.4 RegFile.scala 76:16:@147897.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@147896.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@147900.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@147894.4]
  assign regs_345_clock = clock; // @[:@147903.4]
  assign regs_345_reset = io_reset; // @[:@147904.4 RegFile.scala 76:16:@147911.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@147910.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@147914.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@147908.4]
  assign regs_346_clock = clock; // @[:@147917.4]
  assign regs_346_reset = io_reset; // @[:@147918.4 RegFile.scala 76:16:@147925.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@147924.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@147928.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@147922.4]
  assign regs_347_clock = clock; // @[:@147931.4]
  assign regs_347_reset = io_reset; // @[:@147932.4 RegFile.scala 76:16:@147939.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@147938.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@147942.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@147936.4]
  assign regs_348_clock = clock; // @[:@147945.4]
  assign regs_348_reset = io_reset; // @[:@147946.4 RegFile.scala 76:16:@147953.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@147952.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@147956.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@147950.4]
  assign regs_349_clock = clock; // @[:@147959.4]
  assign regs_349_reset = io_reset; // @[:@147960.4 RegFile.scala 76:16:@147967.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@147966.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@147970.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@147964.4]
  assign regs_350_clock = clock; // @[:@147973.4]
  assign regs_350_reset = io_reset; // @[:@147974.4 RegFile.scala 76:16:@147981.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@147980.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@147984.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@147978.4]
  assign regs_351_clock = clock; // @[:@147987.4]
  assign regs_351_reset = io_reset; // @[:@147988.4 RegFile.scala 76:16:@147995.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@147994.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@147998.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@147992.4]
  assign regs_352_clock = clock; // @[:@148001.4]
  assign regs_352_reset = io_reset; // @[:@148002.4 RegFile.scala 76:16:@148009.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@148008.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@148012.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@148006.4]
  assign regs_353_clock = clock; // @[:@148015.4]
  assign regs_353_reset = io_reset; // @[:@148016.4 RegFile.scala 76:16:@148023.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@148022.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@148026.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@148020.4]
  assign regs_354_clock = clock; // @[:@148029.4]
  assign regs_354_reset = io_reset; // @[:@148030.4 RegFile.scala 76:16:@148037.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@148036.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@148040.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@148034.4]
  assign regs_355_clock = clock; // @[:@148043.4]
  assign regs_355_reset = io_reset; // @[:@148044.4 RegFile.scala 76:16:@148051.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@148050.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@148054.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@148048.4]
  assign regs_356_clock = clock; // @[:@148057.4]
  assign regs_356_reset = io_reset; // @[:@148058.4 RegFile.scala 76:16:@148065.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@148064.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@148068.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@148062.4]
  assign regs_357_clock = clock; // @[:@148071.4]
  assign regs_357_reset = io_reset; // @[:@148072.4 RegFile.scala 76:16:@148079.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@148078.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@148082.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@148076.4]
  assign regs_358_clock = clock; // @[:@148085.4]
  assign regs_358_reset = io_reset; // @[:@148086.4 RegFile.scala 76:16:@148093.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@148092.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@148096.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@148090.4]
  assign regs_359_clock = clock; // @[:@148099.4]
  assign regs_359_reset = io_reset; // @[:@148100.4 RegFile.scala 76:16:@148107.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@148106.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@148110.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@148104.4]
  assign regs_360_clock = clock; // @[:@148113.4]
  assign regs_360_reset = io_reset; // @[:@148114.4 RegFile.scala 76:16:@148121.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@148120.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@148124.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@148118.4]
  assign regs_361_clock = clock; // @[:@148127.4]
  assign regs_361_reset = io_reset; // @[:@148128.4 RegFile.scala 76:16:@148135.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@148134.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@148138.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@148132.4]
  assign regs_362_clock = clock; // @[:@148141.4]
  assign regs_362_reset = io_reset; // @[:@148142.4 RegFile.scala 76:16:@148149.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@148148.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@148152.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@148146.4]
  assign regs_363_clock = clock; // @[:@148155.4]
  assign regs_363_reset = io_reset; // @[:@148156.4 RegFile.scala 76:16:@148163.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@148162.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@148166.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@148160.4]
  assign regs_364_clock = clock; // @[:@148169.4]
  assign regs_364_reset = io_reset; // @[:@148170.4 RegFile.scala 76:16:@148177.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@148176.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@148180.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@148174.4]
  assign regs_365_clock = clock; // @[:@148183.4]
  assign regs_365_reset = io_reset; // @[:@148184.4 RegFile.scala 76:16:@148191.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@148190.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@148194.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@148188.4]
  assign regs_366_clock = clock; // @[:@148197.4]
  assign regs_366_reset = io_reset; // @[:@148198.4 RegFile.scala 76:16:@148205.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@148204.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@148208.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@148202.4]
  assign regs_367_clock = clock; // @[:@148211.4]
  assign regs_367_reset = io_reset; // @[:@148212.4 RegFile.scala 76:16:@148219.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@148218.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@148222.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@148216.4]
  assign regs_368_clock = clock; // @[:@148225.4]
  assign regs_368_reset = io_reset; // @[:@148226.4 RegFile.scala 76:16:@148233.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@148232.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@148236.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@148230.4]
  assign regs_369_clock = clock; // @[:@148239.4]
  assign regs_369_reset = io_reset; // @[:@148240.4 RegFile.scala 76:16:@148247.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@148246.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@148250.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@148244.4]
  assign regs_370_clock = clock; // @[:@148253.4]
  assign regs_370_reset = io_reset; // @[:@148254.4 RegFile.scala 76:16:@148261.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@148260.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@148264.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@148258.4]
  assign regs_371_clock = clock; // @[:@148267.4]
  assign regs_371_reset = io_reset; // @[:@148268.4 RegFile.scala 76:16:@148275.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@148274.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@148278.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@148272.4]
  assign regs_372_clock = clock; // @[:@148281.4]
  assign regs_372_reset = io_reset; // @[:@148282.4 RegFile.scala 76:16:@148289.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@148288.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@148292.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@148286.4]
  assign regs_373_clock = clock; // @[:@148295.4]
  assign regs_373_reset = io_reset; // @[:@148296.4 RegFile.scala 76:16:@148303.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@148302.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@148306.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@148300.4]
  assign regs_374_clock = clock; // @[:@148309.4]
  assign regs_374_reset = io_reset; // @[:@148310.4 RegFile.scala 76:16:@148317.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@148316.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@148320.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@148314.4]
  assign regs_375_clock = clock; // @[:@148323.4]
  assign regs_375_reset = io_reset; // @[:@148324.4 RegFile.scala 76:16:@148331.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@148330.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@148334.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@148328.4]
  assign regs_376_clock = clock; // @[:@148337.4]
  assign regs_376_reset = io_reset; // @[:@148338.4 RegFile.scala 76:16:@148345.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@148344.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@148348.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@148342.4]
  assign regs_377_clock = clock; // @[:@148351.4]
  assign regs_377_reset = io_reset; // @[:@148352.4 RegFile.scala 76:16:@148359.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@148358.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@148362.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@148356.4]
  assign regs_378_clock = clock; // @[:@148365.4]
  assign regs_378_reset = io_reset; // @[:@148366.4 RegFile.scala 76:16:@148373.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@148372.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@148376.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@148370.4]
  assign regs_379_clock = clock; // @[:@148379.4]
  assign regs_379_reset = io_reset; // @[:@148380.4 RegFile.scala 76:16:@148387.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@148386.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@148390.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@148384.4]
  assign regs_380_clock = clock; // @[:@148393.4]
  assign regs_380_reset = io_reset; // @[:@148394.4 RegFile.scala 76:16:@148401.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@148400.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@148404.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@148398.4]
  assign regs_381_clock = clock; // @[:@148407.4]
  assign regs_381_reset = io_reset; // @[:@148408.4 RegFile.scala 76:16:@148415.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@148414.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@148418.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@148412.4]
  assign regs_382_clock = clock; // @[:@148421.4]
  assign regs_382_reset = io_reset; // @[:@148422.4 RegFile.scala 76:16:@148429.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@148428.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@148432.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@148426.4]
  assign regs_383_clock = clock; // @[:@148435.4]
  assign regs_383_reset = io_reset; // @[:@148436.4 RegFile.scala 76:16:@148443.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@148442.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@148446.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@148440.4]
  assign regs_384_clock = clock; // @[:@148449.4]
  assign regs_384_reset = io_reset; // @[:@148450.4 RegFile.scala 76:16:@148457.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@148456.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@148460.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@148454.4]
  assign regs_385_clock = clock; // @[:@148463.4]
  assign regs_385_reset = io_reset; // @[:@148464.4 RegFile.scala 76:16:@148471.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@148470.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@148474.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@148468.4]
  assign regs_386_clock = clock; // @[:@148477.4]
  assign regs_386_reset = io_reset; // @[:@148478.4 RegFile.scala 76:16:@148485.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@148484.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@148488.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@148482.4]
  assign regs_387_clock = clock; // @[:@148491.4]
  assign regs_387_reset = io_reset; // @[:@148492.4 RegFile.scala 76:16:@148499.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@148498.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@148502.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@148496.4]
  assign regs_388_clock = clock; // @[:@148505.4]
  assign regs_388_reset = io_reset; // @[:@148506.4 RegFile.scala 76:16:@148513.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@148512.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@148516.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@148510.4]
  assign regs_389_clock = clock; // @[:@148519.4]
  assign regs_389_reset = io_reset; // @[:@148520.4 RegFile.scala 76:16:@148527.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@148526.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@148530.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@148524.4]
  assign regs_390_clock = clock; // @[:@148533.4]
  assign regs_390_reset = io_reset; // @[:@148534.4 RegFile.scala 76:16:@148541.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@148540.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@148544.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@148538.4]
  assign regs_391_clock = clock; // @[:@148547.4]
  assign regs_391_reset = io_reset; // @[:@148548.4 RegFile.scala 76:16:@148555.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@148554.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@148558.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@148552.4]
  assign regs_392_clock = clock; // @[:@148561.4]
  assign regs_392_reset = io_reset; // @[:@148562.4 RegFile.scala 76:16:@148569.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@148568.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@148572.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@148566.4]
  assign regs_393_clock = clock; // @[:@148575.4]
  assign regs_393_reset = io_reset; // @[:@148576.4 RegFile.scala 76:16:@148583.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@148582.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@148586.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@148580.4]
  assign regs_394_clock = clock; // @[:@148589.4]
  assign regs_394_reset = io_reset; // @[:@148590.4 RegFile.scala 76:16:@148597.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@148596.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@148600.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@148594.4]
  assign regs_395_clock = clock; // @[:@148603.4]
  assign regs_395_reset = io_reset; // @[:@148604.4 RegFile.scala 76:16:@148611.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@148610.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@148614.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@148608.4]
  assign regs_396_clock = clock; // @[:@148617.4]
  assign regs_396_reset = io_reset; // @[:@148618.4 RegFile.scala 76:16:@148625.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@148624.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@148628.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@148622.4]
  assign regs_397_clock = clock; // @[:@148631.4]
  assign regs_397_reset = io_reset; // @[:@148632.4 RegFile.scala 76:16:@148639.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@148638.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@148642.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@148636.4]
  assign regs_398_clock = clock; // @[:@148645.4]
  assign regs_398_reset = io_reset; // @[:@148646.4 RegFile.scala 76:16:@148653.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@148652.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@148656.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@148650.4]
  assign regs_399_clock = clock; // @[:@148659.4]
  assign regs_399_reset = io_reset; // @[:@148660.4 RegFile.scala 76:16:@148667.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@148666.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@148670.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@148664.4]
  assign regs_400_clock = clock; // @[:@148673.4]
  assign regs_400_reset = io_reset; // @[:@148674.4 RegFile.scala 76:16:@148681.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@148680.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@148684.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@148678.4]
  assign regs_401_clock = clock; // @[:@148687.4]
  assign regs_401_reset = io_reset; // @[:@148688.4 RegFile.scala 76:16:@148695.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@148694.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@148698.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@148692.4]
  assign regs_402_clock = clock; // @[:@148701.4]
  assign regs_402_reset = io_reset; // @[:@148702.4 RegFile.scala 76:16:@148709.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@148708.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@148712.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@148706.4]
  assign regs_403_clock = clock; // @[:@148715.4]
  assign regs_403_reset = io_reset; // @[:@148716.4 RegFile.scala 76:16:@148723.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@148722.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@148726.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@148720.4]
  assign regs_404_clock = clock; // @[:@148729.4]
  assign regs_404_reset = io_reset; // @[:@148730.4 RegFile.scala 76:16:@148737.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@148736.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@148740.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@148734.4]
  assign regs_405_clock = clock; // @[:@148743.4]
  assign regs_405_reset = io_reset; // @[:@148744.4 RegFile.scala 76:16:@148751.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@148750.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@148754.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@148748.4]
  assign regs_406_clock = clock; // @[:@148757.4]
  assign regs_406_reset = io_reset; // @[:@148758.4 RegFile.scala 76:16:@148765.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@148764.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@148768.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@148762.4]
  assign regs_407_clock = clock; // @[:@148771.4]
  assign regs_407_reset = io_reset; // @[:@148772.4 RegFile.scala 76:16:@148779.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@148778.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@148782.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@148776.4]
  assign regs_408_clock = clock; // @[:@148785.4]
  assign regs_408_reset = io_reset; // @[:@148786.4 RegFile.scala 76:16:@148793.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@148792.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@148796.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@148790.4]
  assign regs_409_clock = clock; // @[:@148799.4]
  assign regs_409_reset = io_reset; // @[:@148800.4 RegFile.scala 76:16:@148807.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@148806.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@148810.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@148804.4]
  assign regs_410_clock = clock; // @[:@148813.4]
  assign regs_410_reset = io_reset; // @[:@148814.4 RegFile.scala 76:16:@148821.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@148820.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@148824.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@148818.4]
  assign regs_411_clock = clock; // @[:@148827.4]
  assign regs_411_reset = io_reset; // @[:@148828.4 RegFile.scala 76:16:@148835.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@148834.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@148838.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@148832.4]
  assign regs_412_clock = clock; // @[:@148841.4]
  assign regs_412_reset = io_reset; // @[:@148842.4 RegFile.scala 76:16:@148849.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@148848.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@148852.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@148846.4]
  assign regs_413_clock = clock; // @[:@148855.4]
  assign regs_413_reset = io_reset; // @[:@148856.4 RegFile.scala 76:16:@148863.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@148862.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@148866.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@148860.4]
  assign regs_414_clock = clock; // @[:@148869.4]
  assign regs_414_reset = io_reset; // @[:@148870.4 RegFile.scala 76:16:@148877.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@148876.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@148880.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@148874.4]
  assign regs_415_clock = clock; // @[:@148883.4]
  assign regs_415_reset = io_reset; // @[:@148884.4 RegFile.scala 76:16:@148891.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@148890.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@148894.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@148888.4]
  assign regs_416_clock = clock; // @[:@148897.4]
  assign regs_416_reset = io_reset; // @[:@148898.4 RegFile.scala 76:16:@148905.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@148904.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@148908.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@148902.4]
  assign regs_417_clock = clock; // @[:@148911.4]
  assign regs_417_reset = io_reset; // @[:@148912.4 RegFile.scala 76:16:@148919.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@148918.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@148922.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@148916.4]
  assign regs_418_clock = clock; // @[:@148925.4]
  assign regs_418_reset = io_reset; // @[:@148926.4 RegFile.scala 76:16:@148933.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@148932.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@148936.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@148930.4]
  assign regs_419_clock = clock; // @[:@148939.4]
  assign regs_419_reset = io_reset; // @[:@148940.4 RegFile.scala 76:16:@148947.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@148946.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@148950.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@148944.4]
  assign regs_420_clock = clock; // @[:@148953.4]
  assign regs_420_reset = io_reset; // @[:@148954.4 RegFile.scala 76:16:@148961.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@148960.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@148964.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@148958.4]
  assign regs_421_clock = clock; // @[:@148967.4]
  assign regs_421_reset = io_reset; // @[:@148968.4 RegFile.scala 76:16:@148975.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@148974.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@148978.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@148972.4]
  assign regs_422_clock = clock; // @[:@148981.4]
  assign regs_422_reset = io_reset; // @[:@148982.4 RegFile.scala 76:16:@148989.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@148988.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@148992.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@148986.4]
  assign regs_423_clock = clock; // @[:@148995.4]
  assign regs_423_reset = io_reset; // @[:@148996.4 RegFile.scala 76:16:@149003.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@149002.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@149006.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@149000.4]
  assign regs_424_clock = clock; // @[:@149009.4]
  assign regs_424_reset = io_reset; // @[:@149010.4 RegFile.scala 76:16:@149017.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@149016.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@149020.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@149014.4]
  assign regs_425_clock = clock; // @[:@149023.4]
  assign regs_425_reset = io_reset; // @[:@149024.4 RegFile.scala 76:16:@149031.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@149030.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@149034.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@149028.4]
  assign regs_426_clock = clock; // @[:@149037.4]
  assign regs_426_reset = io_reset; // @[:@149038.4 RegFile.scala 76:16:@149045.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@149044.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@149048.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@149042.4]
  assign regs_427_clock = clock; // @[:@149051.4]
  assign regs_427_reset = io_reset; // @[:@149052.4 RegFile.scala 76:16:@149059.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@149058.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@149062.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@149056.4]
  assign regs_428_clock = clock; // @[:@149065.4]
  assign regs_428_reset = io_reset; // @[:@149066.4 RegFile.scala 76:16:@149073.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@149072.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@149076.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@149070.4]
  assign regs_429_clock = clock; // @[:@149079.4]
  assign regs_429_reset = io_reset; // @[:@149080.4 RegFile.scala 76:16:@149087.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@149086.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@149090.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@149084.4]
  assign regs_430_clock = clock; // @[:@149093.4]
  assign regs_430_reset = io_reset; // @[:@149094.4 RegFile.scala 76:16:@149101.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@149100.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@149104.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@149098.4]
  assign regs_431_clock = clock; // @[:@149107.4]
  assign regs_431_reset = io_reset; // @[:@149108.4 RegFile.scala 76:16:@149115.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@149114.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@149118.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@149112.4]
  assign regs_432_clock = clock; // @[:@149121.4]
  assign regs_432_reset = io_reset; // @[:@149122.4 RegFile.scala 76:16:@149129.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@149128.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@149132.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@149126.4]
  assign regs_433_clock = clock; // @[:@149135.4]
  assign regs_433_reset = io_reset; // @[:@149136.4 RegFile.scala 76:16:@149143.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@149142.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@149146.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@149140.4]
  assign regs_434_clock = clock; // @[:@149149.4]
  assign regs_434_reset = io_reset; // @[:@149150.4 RegFile.scala 76:16:@149157.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@149156.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@149160.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@149154.4]
  assign regs_435_clock = clock; // @[:@149163.4]
  assign regs_435_reset = io_reset; // @[:@149164.4 RegFile.scala 76:16:@149171.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@149170.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@149174.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@149168.4]
  assign regs_436_clock = clock; // @[:@149177.4]
  assign regs_436_reset = io_reset; // @[:@149178.4 RegFile.scala 76:16:@149185.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@149184.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@149188.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@149182.4]
  assign regs_437_clock = clock; // @[:@149191.4]
  assign regs_437_reset = io_reset; // @[:@149192.4 RegFile.scala 76:16:@149199.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@149198.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@149202.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@149196.4]
  assign regs_438_clock = clock; // @[:@149205.4]
  assign regs_438_reset = io_reset; // @[:@149206.4 RegFile.scala 76:16:@149213.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@149212.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@149216.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@149210.4]
  assign regs_439_clock = clock; // @[:@149219.4]
  assign regs_439_reset = io_reset; // @[:@149220.4 RegFile.scala 76:16:@149227.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@149226.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@149230.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@149224.4]
  assign regs_440_clock = clock; // @[:@149233.4]
  assign regs_440_reset = io_reset; // @[:@149234.4 RegFile.scala 76:16:@149241.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@149240.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@149244.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@149238.4]
  assign regs_441_clock = clock; // @[:@149247.4]
  assign regs_441_reset = io_reset; // @[:@149248.4 RegFile.scala 76:16:@149255.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@149254.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@149258.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@149252.4]
  assign regs_442_clock = clock; // @[:@149261.4]
  assign regs_442_reset = io_reset; // @[:@149262.4 RegFile.scala 76:16:@149269.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@149268.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@149272.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@149266.4]
  assign regs_443_clock = clock; // @[:@149275.4]
  assign regs_443_reset = io_reset; // @[:@149276.4 RegFile.scala 76:16:@149283.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@149282.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@149286.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@149280.4]
  assign regs_444_clock = clock; // @[:@149289.4]
  assign regs_444_reset = io_reset; // @[:@149290.4 RegFile.scala 76:16:@149297.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@149296.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@149300.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@149294.4]
  assign regs_445_clock = clock; // @[:@149303.4]
  assign regs_445_reset = io_reset; // @[:@149304.4 RegFile.scala 76:16:@149311.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@149310.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@149314.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@149308.4]
  assign regs_446_clock = clock; // @[:@149317.4]
  assign regs_446_reset = io_reset; // @[:@149318.4 RegFile.scala 76:16:@149325.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@149324.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@149328.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@149322.4]
  assign regs_447_clock = clock; // @[:@149331.4]
  assign regs_447_reset = io_reset; // @[:@149332.4 RegFile.scala 76:16:@149339.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@149338.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@149342.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@149336.4]
  assign regs_448_clock = clock; // @[:@149345.4]
  assign regs_448_reset = io_reset; // @[:@149346.4 RegFile.scala 76:16:@149353.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@149352.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@149356.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@149350.4]
  assign regs_449_clock = clock; // @[:@149359.4]
  assign regs_449_reset = io_reset; // @[:@149360.4 RegFile.scala 76:16:@149367.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@149366.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@149370.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@149364.4]
  assign regs_450_clock = clock; // @[:@149373.4]
  assign regs_450_reset = io_reset; // @[:@149374.4 RegFile.scala 76:16:@149381.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@149380.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@149384.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@149378.4]
  assign regs_451_clock = clock; // @[:@149387.4]
  assign regs_451_reset = io_reset; // @[:@149388.4 RegFile.scala 76:16:@149395.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@149394.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@149398.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@149392.4]
  assign regs_452_clock = clock; // @[:@149401.4]
  assign regs_452_reset = io_reset; // @[:@149402.4 RegFile.scala 76:16:@149409.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@149408.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@149412.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@149406.4]
  assign regs_453_clock = clock; // @[:@149415.4]
  assign regs_453_reset = io_reset; // @[:@149416.4 RegFile.scala 76:16:@149423.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@149422.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@149426.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@149420.4]
  assign regs_454_clock = clock; // @[:@149429.4]
  assign regs_454_reset = io_reset; // @[:@149430.4 RegFile.scala 76:16:@149437.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@149436.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@149440.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@149434.4]
  assign regs_455_clock = clock; // @[:@149443.4]
  assign regs_455_reset = io_reset; // @[:@149444.4 RegFile.scala 76:16:@149451.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@149450.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@149454.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@149448.4]
  assign regs_456_clock = clock; // @[:@149457.4]
  assign regs_456_reset = io_reset; // @[:@149458.4 RegFile.scala 76:16:@149465.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@149464.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@149468.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@149462.4]
  assign regs_457_clock = clock; // @[:@149471.4]
  assign regs_457_reset = io_reset; // @[:@149472.4 RegFile.scala 76:16:@149479.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@149478.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@149482.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@149476.4]
  assign regs_458_clock = clock; // @[:@149485.4]
  assign regs_458_reset = io_reset; // @[:@149486.4 RegFile.scala 76:16:@149493.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@149492.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@149496.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@149490.4]
  assign regs_459_clock = clock; // @[:@149499.4]
  assign regs_459_reset = io_reset; // @[:@149500.4 RegFile.scala 76:16:@149507.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@149506.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@149510.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@149504.4]
  assign regs_460_clock = clock; // @[:@149513.4]
  assign regs_460_reset = io_reset; // @[:@149514.4 RegFile.scala 76:16:@149521.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@149520.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@149524.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@149518.4]
  assign regs_461_clock = clock; // @[:@149527.4]
  assign regs_461_reset = io_reset; // @[:@149528.4 RegFile.scala 76:16:@149535.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@149534.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@149538.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@149532.4]
  assign regs_462_clock = clock; // @[:@149541.4]
  assign regs_462_reset = io_reset; // @[:@149542.4 RegFile.scala 76:16:@149549.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@149548.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@149552.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@149546.4]
  assign regs_463_clock = clock; // @[:@149555.4]
  assign regs_463_reset = io_reset; // @[:@149556.4 RegFile.scala 76:16:@149563.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@149562.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@149566.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@149560.4]
  assign regs_464_clock = clock; // @[:@149569.4]
  assign regs_464_reset = io_reset; // @[:@149570.4 RegFile.scala 76:16:@149577.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@149576.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@149580.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@149574.4]
  assign regs_465_clock = clock; // @[:@149583.4]
  assign regs_465_reset = io_reset; // @[:@149584.4 RegFile.scala 76:16:@149591.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@149590.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@149594.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@149588.4]
  assign regs_466_clock = clock; // @[:@149597.4]
  assign regs_466_reset = io_reset; // @[:@149598.4 RegFile.scala 76:16:@149605.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@149604.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@149608.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@149602.4]
  assign regs_467_clock = clock; // @[:@149611.4]
  assign regs_467_reset = io_reset; // @[:@149612.4 RegFile.scala 76:16:@149619.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@149618.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@149622.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@149616.4]
  assign regs_468_clock = clock; // @[:@149625.4]
  assign regs_468_reset = io_reset; // @[:@149626.4 RegFile.scala 76:16:@149633.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@149632.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@149636.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@149630.4]
  assign regs_469_clock = clock; // @[:@149639.4]
  assign regs_469_reset = io_reset; // @[:@149640.4 RegFile.scala 76:16:@149647.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@149646.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@149650.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@149644.4]
  assign regs_470_clock = clock; // @[:@149653.4]
  assign regs_470_reset = io_reset; // @[:@149654.4 RegFile.scala 76:16:@149661.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@149660.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@149664.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@149658.4]
  assign regs_471_clock = clock; // @[:@149667.4]
  assign regs_471_reset = io_reset; // @[:@149668.4 RegFile.scala 76:16:@149675.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@149674.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@149678.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@149672.4]
  assign regs_472_clock = clock; // @[:@149681.4]
  assign regs_472_reset = io_reset; // @[:@149682.4 RegFile.scala 76:16:@149689.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@149688.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@149692.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@149686.4]
  assign regs_473_clock = clock; // @[:@149695.4]
  assign regs_473_reset = io_reset; // @[:@149696.4 RegFile.scala 76:16:@149703.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@149702.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@149706.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@149700.4]
  assign regs_474_clock = clock; // @[:@149709.4]
  assign regs_474_reset = io_reset; // @[:@149710.4 RegFile.scala 76:16:@149717.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@149716.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@149720.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@149714.4]
  assign regs_475_clock = clock; // @[:@149723.4]
  assign regs_475_reset = io_reset; // @[:@149724.4 RegFile.scala 76:16:@149731.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@149730.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@149734.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@149728.4]
  assign regs_476_clock = clock; // @[:@149737.4]
  assign regs_476_reset = io_reset; // @[:@149738.4 RegFile.scala 76:16:@149745.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@149744.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@149748.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@149742.4]
  assign regs_477_clock = clock; // @[:@149751.4]
  assign regs_477_reset = io_reset; // @[:@149752.4 RegFile.scala 76:16:@149759.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@149758.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@149762.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@149756.4]
  assign regs_478_clock = clock; // @[:@149765.4]
  assign regs_478_reset = io_reset; // @[:@149766.4 RegFile.scala 76:16:@149773.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@149772.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@149776.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@149770.4]
  assign regs_479_clock = clock; // @[:@149779.4]
  assign regs_479_reset = io_reset; // @[:@149780.4 RegFile.scala 76:16:@149787.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@149786.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@149790.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@149784.4]
  assign regs_480_clock = clock; // @[:@149793.4]
  assign regs_480_reset = io_reset; // @[:@149794.4 RegFile.scala 76:16:@149801.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@149800.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@149804.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@149798.4]
  assign regs_481_clock = clock; // @[:@149807.4]
  assign regs_481_reset = io_reset; // @[:@149808.4 RegFile.scala 76:16:@149815.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@149814.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@149818.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@149812.4]
  assign regs_482_clock = clock; // @[:@149821.4]
  assign regs_482_reset = io_reset; // @[:@149822.4 RegFile.scala 76:16:@149829.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@149828.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@149832.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@149826.4]
  assign regs_483_clock = clock; // @[:@149835.4]
  assign regs_483_reset = io_reset; // @[:@149836.4 RegFile.scala 76:16:@149843.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@149842.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@149846.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@149840.4]
  assign regs_484_clock = clock; // @[:@149849.4]
  assign regs_484_reset = io_reset; // @[:@149850.4 RegFile.scala 76:16:@149857.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@149856.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@149860.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@149854.4]
  assign regs_485_clock = clock; // @[:@149863.4]
  assign regs_485_reset = io_reset; // @[:@149864.4 RegFile.scala 76:16:@149871.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@149870.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@149874.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@149868.4]
  assign regs_486_clock = clock; // @[:@149877.4]
  assign regs_486_reset = io_reset; // @[:@149878.4 RegFile.scala 76:16:@149885.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@149884.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@149888.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@149882.4]
  assign regs_487_clock = clock; // @[:@149891.4]
  assign regs_487_reset = io_reset; // @[:@149892.4 RegFile.scala 76:16:@149899.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@149898.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@149902.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@149896.4]
  assign regs_488_clock = clock; // @[:@149905.4]
  assign regs_488_reset = io_reset; // @[:@149906.4 RegFile.scala 76:16:@149913.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@149912.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@149916.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@149910.4]
  assign regs_489_clock = clock; // @[:@149919.4]
  assign regs_489_reset = io_reset; // @[:@149920.4 RegFile.scala 76:16:@149927.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@149926.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@149930.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@149924.4]
  assign regs_490_clock = clock; // @[:@149933.4]
  assign regs_490_reset = io_reset; // @[:@149934.4 RegFile.scala 76:16:@149941.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@149940.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@149944.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@149938.4]
  assign regs_491_clock = clock; // @[:@149947.4]
  assign regs_491_reset = io_reset; // @[:@149948.4 RegFile.scala 76:16:@149955.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@149954.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@149958.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@149952.4]
  assign regs_492_clock = clock; // @[:@149961.4]
  assign regs_492_reset = io_reset; // @[:@149962.4 RegFile.scala 76:16:@149969.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@149968.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@149972.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@149966.4]
  assign regs_493_clock = clock; // @[:@149975.4]
  assign regs_493_reset = io_reset; // @[:@149976.4 RegFile.scala 76:16:@149983.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@149982.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@149986.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@149980.4]
  assign regs_494_clock = clock; // @[:@149989.4]
  assign regs_494_reset = io_reset; // @[:@149990.4 RegFile.scala 76:16:@149997.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@149996.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@150000.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@149994.4]
  assign regs_495_clock = clock; // @[:@150003.4]
  assign regs_495_reset = io_reset; // @[:@150004.4 RegFile.scala 76:16:@150011.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@150010.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@150014.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@150008.4]
  assign regs_496_clock = clock; // @[:@150017.4]
  assign regs_496_reset = io_reset; // @[:@150018.4 RegFile.scala 76:16:@150025.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@150024.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@150028.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@150022.4]
  assign regs_497_clock = clock; // @[:@150031.4]
  assign regs_497_reset = io_reset; // @[:@150032.4 RegFile.scala 76:16:@150039.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@150038.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@150042.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@150036.4]
  assign regs_498_clock = clock; // @[:@150045.4]
  assign regs_498_reset = io_reset; // @[:@150046.4 RegFile.scala 76:16:@150053.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@150052.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@150056.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@150050.4]
  assign regs_499_clock = clock; // @[:@150059.4]
  assign regs_499_reset = io_reset; // @[:@150060.4 RegFile.scala 76:16:@150067.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@150066.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@150070.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@150064.4]
  assign regs_500_clock = clock; // @[:@150073.4]
  assign regs_500_reset = io_reset; // @[:@150074.4 RegFile.scala 76:16:@150081.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@150080.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@150084.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@150078.4]
  assign regs_501_clock = clock; // @[:@150087.4]
  assign regs_501_reset = io_reset; // @[:@150088.4 RegFile.scala 76:16:@150095.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@150094.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@150098.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@150092.4]
  assign regs_502_clock = clock; // @[:@150101.4]
  assign regs_502_reset = io_reset; // @[:@150102.4 RegFile.scala 76:16:@150109.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@150108.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@150112.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@150106.4]
  assign regs_503_clock = clock; // @[:@150115.4]
  assign regs_503_reset = io_reset; // @[:@150116.4 RegFile.scala 76:16:@150123.4]
  assign regs_503_io_in = 64'h0; // @[RegFile.scala 75:16:@150122.4]
  assign regs_503_io_reset = reset; // @[RegFile.scala 78:19:@150126.4]
  assign regs_503_io_enable = 1'h1; // @[RegFile.scala 74:20:@150120.4]
  assign regs_504_clock = clock; // @[:@150129.4]
  assign regs_504_reset = io_reset; // @[:@150130.4 RegFile.scala 76:16:@150137.4]
  assign regs_504_io_in = 64'h0; // @[RegFile.scala 75:16:@150136.4]
  assign regs_504_io_reset = reset; // @[RegFile.scala 78:19:@150140.4]
  assign regs_504_io_enable = 1'h1; // @[RegFile.scala 74:20:@150134.4]
  assign regs_505_clock = clock; // @[:@150143.4]
  assign regs_505_reset = io_reset; // @[:@150144.4 RegFile.scala 76:16:@150151.4]
  assign regs_505_io_in = 64'h0; // @[RegFile.scala 75:16:@150150.4]
  assign regs_505_io_reset = reset; // @[RegFile.scala 78:19:@150154.4]
  assign regs_505_io_enable = 1'h1; // @[RegFile.scala 74:20:@150148.4]
  assign regs_506_clock = clock; // @[:@150157.4]
  assign regs_506_reset = io_reset; // @[:@150158.4 RegFile.scala 76:16:@150165.4]
  assign regs_506_io_in = 64'h0; // @[RegFile.scala 75:16:@150164.4]
  assign regs_506_io_reset = reset; // @[RegFile.scala 78:19:@150168.4]
  assign regs_506_io_enable = 1'h1; // @[RegFile.scala 74:20:@150162.4]
  assign regs_507_clock = clock; // @[:@150171.4]
  assign regs_507_reset = io_reset; // @[:@150172.4 RegFile.scala 76:16:@150179.4]
  assign regs_507_io_in = 64'h0; // @[RegFile.scala 75:16:@150178.4]
  assign regs_507_io_reset = reset; // @[RegFile.scala 78:19:@150182.4]
  assign regs_507_io_enable = 1'h1; // @[RegFile.scala 74:20:@150176.4]
  assign regs_508_clock = clock; // @[:@150185.4]
  assign regs_508_reset = io_reset; // @[:@150186.4 RegFile.scala 76:16:@150193.4]
  assign regs_508_io_in = 64'h0; // @[RegFile.scala 75:16:@150192.4]
  assign regs_508_io_reset = reset; // @[RegFile.scala 78:19:@150196.4]
  assign regs_508_io_enable = 1'h1; // @[RegFile.scala 74:20:@150190.4]
  assign regs_509_clock = clock; // @[:@150199.4]
  assign regs_509_reset = io_reset; // @[:@150200.4 RegFile.scala 76:16:@150207.4]
  assign regs_509_io_in = 64'h0; // @[RegFile.scala 75:16:@150206.4]
  assign regs_509_io_reset = reset; // @[RegFile.scala 78:19:@150210.4]
  assign regs_509_io_enable = 1'h1; // @[RegFile.scala 74:20:@150204.4]
  assign regs_510_clock = clock; // @[:@150213.4]
  assign regs_510_reset = io_reset; // @[:@150214.4 RegFile.scala 76:16:@150221.4]
  assign regs_510_io_in = 64'h0; // @[RegFile.scala 75:16:@150220.4]
  assign regs_510_io_reset = reset; // @[RegFile.scala 78:19:@150224.4]
  assign regs_510_io_enable = 1'h1; // @[RegFile.scala 74:20:@150218.4]
  assign regs_511_clock = clock; // @[:@150227.4]
  assign regs_511_reset = io_reset; // @[:@150228.4 RegFile.scala 76:16:@150235.4]
  assign regs_511_io_in = 64'h0; // @[RegFile.scala 75:16:@150234.4]
  assign regs_511_io_reset = reset; // @[RegFile.scala 78:19:@150238.4]
  assign regs_511_io_enable = 1'h1; // @[RegFile.scala 74:20:@150232.4]
  assign regs_512_clock = clock; // @[:@150241.4]
  assign regs_512_reset = io_reset; // @[:@150242.4 RegFile.scala 76:16:@150249.4]
  assign regs_512_io_in = 64'h0; // @[RegFile.scala 75:16:@150248.4]
  assign regs_512_io_reset = reset; // @[RegFile.scala 78:19:@150252.4]
  assign regs_512_io_enable = 1'h1; // @[RegFile.scala 74:20:@150246.4]
  assign regs_513_clock = clock; // @[:@150255.4]
  assign regs_513_reset = io_reset; // @[:@150256.4 RegFile.scala 76:16:@150263.4]
  assign regs_513_io_in = 64'h0; // @[RegFile.scala 75:16:@150262.4]
  assign regs_513_io_reset = reset; // @[RegFile.scala 78:19:@150266.4]
  assign regs_513_io_enable = 1'h1; // @[RegFile.scala 74:20:@150260.4]
  assign regs_514_clock = clock; // @[:@150269.4]
  assign regs_514_reset = io_reset; // @[:@150270.4 RegFile.scala 76:16:@150277.4]
  assign regs_514_io_in = 64'h0; // @[RegFile.scala 75:16:@150276.4]
  assign regs_514_io_reset = reset; // @[RegFile.scala 78:19:@150280.4]
  assign regs_514_io_enable = 1'h1; // @[RegFile.scala 74:20:@150274.4]
  assign regs_515_clock = clock; // @[:@150283.4]
  assign regs_515_reset = io_reset; // @[:@150284.4 RegFile.scala 76:16:@150291.4]
  assign regs_515_io_in = 64'h0; // @[RegFile.scala 75:16:@150290.4]
  assign regs_515_io_reset = reset; // @[RegFile.scala 78:19:@150294.4]
  assign regs_515_io_enable = 1'h1; // @[RegFile.scala 74:20:@150288.4]
  assign regs_516_clock = clock; // @[:@150297.4]
  assign regs_516_reset = io_reset; // @[:@150298.4 RegFile.scala 76:16:@150305.4]
  assign regs_516_io_in = 64'h0; // @[RegFile.scala 75:16:@150304.4]
  assign regs_516_io_reset = reset; // @[RegFile.scala 78:19:@150308.4]
  assign regs_516_io_enable = 1'h1; // @[RegFile.scala 74:20:@150302.4]
  assign regs_517_clock = clock; // @[:@150311.4]
  assign regs_517_reset = io_reset; // @[:@150312.4 RegFile.scala 76:16:@150319.4]
  assign regs_517_io_in = 64'h0; // @[RegFile.scala 75:16:@150318.4]
  assign regs_517_io_reset = reset; // @[RegFile.scala 78:19:@150322.4]
  assign regs_517_io_enable = 1'h1; // @[RegFile.scala 74:20:@150316.4]
  assign regs_518_clock = clock; // @[:@150325.4]
  assign regs_518_reset = io_reset; // @[:@150326.4 RegFile.scala 76:16:@150333.4]
  assign regs_518_io_in = 64'h0; // @[RegFile.scala 75:16:@150332.4]
  assign regs_518_io_reset = reset; // @[RegFile.scala 78:19:@150336.4]
  assign regs_518_io_enable = 1'h1; // @[RegFile.scala 74:20:@150330.4]
  assign regs_519_clock = clock; // @[:@150339.4]
  assign regs_519_reset = io_reset; // @[:@150340.4 RegFile.scala 76:16:@150347.4]
  assign regs_519_io_in = 64'h0; // @[RegFile.scala 75:16:@150346.4]
  assign regs_519_io_reset = reset; // @[RegFile.scala 78:19:@150350.4]
  assign regs_519_io_enable = 1'h1; // @[RegFile.scala 74:20:@150344.4]
  assign regs_520_clock = clock; // @[:@150353.4]
  assign regs_520_reset = io_reset; // @[:@150354.4 RegFile.scala 76:16:@150361.4]
  assign regs_520_io_in = 64'h0; // @[RegFile.scala 75:16:@150360.4]
  assign regs_520_io_reset = reset; // @[RegFile.scala 78:19:@150364.4]
  assign regs_520_io_enable = 1'h1; // @[RegFile.scala 74:20:@150358.4]
  assign regs_521_clock = clock; // @[:@150367.4]
  assign regs_521_reset = io_reset; // @[:@150368.4 RegFile.scala 76:16:@150375.4]
  assign regs_521_io_in = 64'h0; // @[RegFile.scala 75:16:@150374.4]
  assign regs_521_io_reset = reset; // @[RegFile.scala 78:19:@150378.4]
  assign regs_521_io_enable = 1'h1; // @[RegFile.scala 74:20:@150372.4]
  assign regs_522_clock = clock; // @[:@150381.4]
  assign regs_522_reset = io_reset; // @[:@150382.4 RegFile.scala 76:16:@150389.4]
  assign regs_522_io_in = 64'h0; // @[RegFile.scala 75:16:@150388.4]
  assign regs_522_io_reset = reset; // @[RegFile.scala 78:19:@150392.4]
  assign regs_522_io_enable = 1'h1; // @[RegFile.scala 74:20:@150386.4]
  assign regs_523_clock = clock; // @[:@150395.4]
  assign regs_523_reset = io_reset; // @[:@150396.4 RegFile.scala 76:16:@150403.4]
  assign regs_523_io_in = 64'h0; // @[RegFile.scala 75:16:@150402.4]
  assign regs_523_io_reset = reset; // @[RegFile.scala 78:19:@150406.4]
  assign regs_523_io_enable = 1'h1; // @[RegFile.scala 74:20:@150400.4]
  assign regs_524_clock = clock; // @[:@150409.4]
  assign regs_524_reset = io_reset; // @[:@150410.4 RegFile.scala 76:16:@150417.4]
  assign regs_524_io_in = 64'h0; // @[RegFile.scala 75:16:@150416.4]
  assign regs_524_io_reset = reset; // @[RegFile.scala 78:19:@150420.4]
  assign regs_524_io_enable = 1'h1; // @[RegFile.scala 74:20:@150414.4]
  assign regs_525_clock = clock; // @[:@150423.4]
  assign regs_525_reset = io_reset; // @[:@150424.4 RegFile.scala 76:16:@150431.4]
  assign regs_525_io_in = 64'h0; // @[RegFile.scala 75:16:@150430.4]
  assign regs_525_io_reset = reset; // @[RegFile.scala 78:19:@150434.4]
  assign regs_525_io_enable = 1'h1; // @[RegFile.scala 74:20:@150428.4]
  assign regs_526_clock = clock; // @[:@150437.4]
  assign regs_526_reset = io_reset; // @[:@150438.4 RegFile.scala 76:16:@150445.4]
  assign regs_526_io_in = 64'h0; // @[RegFile.scala 75:16:@150444.4]
  assign regs_526_io_reset = reset; // @[RegFile.scala 78:19:@150448.4]
  assign regs_526_io_enable = 1'h1; // @[RegFile.scala 74:20:@150442.4]
  assign regs_527_clock = clock; // @[:@150451.4]
  assign regs_527_reset = io_reset; // @[:@150452.4 RegFile.scala 76:16:@150459.4]
  assign regs_527_io_in = 64'h0; // @[RegFile.scala 75:16:@150458.4]
  assign regs_527_io_reset = reset; // @[RegFile.scala 78:19:@150462.4]
  assign regs_527_io_enable = 1'h1; // @[RegFile.scala 74:20:@150456.4]
  assign regs_528_clock = clock; // @[:@150465.4]
  assign regs_528_reset = io_reset; // @[:@150466.4 RegFile.scala 76:16:@150473.4]
  assign regs_528_io_in = 64'h0; // @[RegFile.scala 75:16:@150472.4]
  assign regs_528_io_reset = reset; // @[RegFile.scala 78:19:@150476.4]
  assign regs_528_io_enable = 1'h1; // @[RegFile.scala 74:20:@150470.4]
  assign regs_529_clock = clock; // @[:@150479.4]
  assign regs_529_reset = io_reset; // @[:@150480.4 RegFile.scala 76:16:@150487.4]
  assign regs_529_io_in = 64'h0; // @[RegFile.scala 75:16:@150486.4]
  assign regs_529_io_reset = reset; // @[RegFile.scala 78:19:@150490.4]
  assign regs_529_io_enable = 1'h1; // @[RegFile.scala 74:20:@150484.4]
  assign regs_530_clock = clock; // @[:@150493.4]
  assign regs_530_reset = io_reset; // @[:@150494.4 RegFile.scala 76:16:@150501.4]
  assign regs_530_io_in = 64'h0; // @[RegFile.scala 75:16:@150500.4]
  assign regs_530_io_reset = reset; // @[RegFile.scala 78:19:@150504.4]
  assign regs_530_io_enable = 1'h1; // @[RegFile.scala 74:20:@150498.4]
  assign regs_531_clock = clock; // @[:@150507.4]
  assign regs_531_reset = io_reset; // @[:@150508.4 RegFile.scala 76:16:@150515.4]
  assign regs_531_io_in = 64'h0; // @[RegFile.scala 75:16:@150514.4]
  assign regs_531_io_reset = reset; // @[RegFile.scala 78:19:@150518.4]
  assign regs_531_io_enable = 1'h1; // @[RegFile.scala 74:20:@150512.4]
  assign regs_532_clock = clock; // @[:@150521.4]
  assign regs_532_reset = io_reset; // @[:@150522.4 RegFile.scala 76:16:@150529.4]
  assign regs_532_io_in = 64'h0; // @[RegFile.scala 75:16:@150528.4]
  assign regs_532_io_reset = reset; // @[RegFile.scala 78:19:@150532.4]
  assign regs_532_io_enable = 1'h1; // @[RegFile.scala 74:20:@150526.4]
  assign regs_533_clock = clock; // @[:@150535.4]
  assign regs_533_reset = io_reset; // @[:@150536.4 RegFile.scala 76:16:@150543.4]
  assign regs_533_io_in = 64'h0; // @[RegFile.scala 75:16:@150542.4]
  assign regs_533_io_reset = reset; // @[RegFile.scala 78:19:@150546.4]
  assign regs_533_io_enable = 1'h1; // @[RegFile.scala 74:20:@150540.4]
  assign regs_534_clock = clock; // @[:@150549.4]
  assign regs_534_reset = io_reset; // @[:@150550.4 RegFile.scala 76:16:@150557.4]
  assign regs_534_io_in = 64'h0; // @[RegFile.scala 75:16:@150556.4]
  assign regs_534_io_reset = reset; // @[RegFile.scala 78:19:@150560.4]
  assign regs_534_io_enable = 1'h1; // @[RegFile.scala 74:20:@150554.4]
  assign regs_535_clock = clock; // @[:@150563.4]
  assign regs_535_reset = io_reset; // @[:@150564.4 RegFile.scala 76:16:@150571.4]
  assign regs_535_io_in = 64'h0; // @[RegFile.scala 75:16:@150570.4]
  assign regs_535_io_reset = reset; // @[RegFile.scala 78:19:@150574.4]
  assign regs_535_io_enable = 1'h1; // @[RegFile.scala 74:20:@150568.4]
  assign regs_536_clock = clock; // @[:@150577.4]
  assign regs_536_reset = io_reset; // @[:@150578.4 RegFile.scala 76:16:@150585.4]
  assign regs_536_io_in = 64'h0; // @[RegFile.scala 75:16:@150584.4]
  assign regs_536_io_reset = reset; // @[RegFile.scala 78:19:@150588.4]
  assign regs_536_io_enable = 1'h1; // @[RegFile.scala 74:20:@150582.4]
  assign regs_537_clock = clock; // @[:@150591.4]
  assign regs_537_reset = io_reset; // @[:@150592.4 RegFile.scala 76:16:@150599.4]
  assign regs_537_io_in = 64'h0; // @[RegFile.scala 75:16:@150598.4]
  assign regs_537_io_reset = reset; // @[RegFile.scala 78:19:@150602.4]
  assign regs_537_io_enable = 1'h1; // @[RegFile.scala 74:20:@150596.4]
  assign regs_538_clock = clock; // @[:@150605.4]
  assign regs_538_reset = io_reset; // @[:@150606.4 RegFile.scala 76:16:@150613.4]
  assign regs_538_io_in = 64'h0; // @[RegFile.scala 75:16:@150612.4]
  assign regs_538_io_reset = reset; // @[RegFile.scala 78:19:@150616.4]
  assign regs_538_io_enable = 1'h1; // @[RegFile.scala 74:20:@150610.4]
  assign regs_539_clock = clock; // @[:@150619.4]
  assign regs_539_reset = io_reset; // @[:@150620.4 RegFile.scala 76:16:@150627.4]
  assign regs_539_io_in = 64'h0; // @[RegFile.scala 75:16:@150626.4]
  assign regs_539_io_reset = reset; // @[RegFile.scala 78:19:@150630.4]
  assign regs_539_io_enable = 1'h1; // @[RegFile.scala 74:20:@150624.4]
  assign regs_540_clock = clock; // @[:@150633.4]
  assign regs_540_reset = io_reset; // @[:@150634.4 RegFile.scala 76:16:@150641.4]
  assign regs_540_io_in = 64'h0; // @[RegFile.scala 75:16:@150640.4]
  assign regs_540_io_reset = reset; // @[RegFile.scala 78:19:@150644.4]
  assign regs_540_io_enable = 1'h1; // @[RegFile.scala 74:20:@150638.4]
  assign regs_541_clock = clock; // @[:@150647.4]
  assign regs_541_reset = io_reset; // @[:@150648.4 RegFile.scala 76:16:@150655.4]
  assign regs_541_io_in = 64'h0; // @[RegFile.scala 75:16:@150654.4]
  assign regs_541_io_reset = reset; // @[RegFile.scala 78:19:@150658.4]
  assign regs_541_io_enable = 1'h1; // @[RegFile.scala 74:20:@150652.4]
  assign regs_542_clock = clock; // @[:@150661.4]
  assign regs_542_reset = io_reset; // @[:@150662.4 RegFile.scala 76:16:@150669.4]
  assign regs_542_io_in = 64'h0; // @[RegFile.scala 75:16:@150668.4]
  assign regs_542_io_reset = reset; // @[RegFile.scala 78:19:@150672.4]
  assign regs_542_io_enable = 1'h1; // @[RegFile.scala 74:20:@150666.4]
  assign regs_543_clock = clock; // @[:@150675.4]
  assign regs_543_reset = io_reset; // @[:@150676.4 RegFile.scala 76:16:@150683.4]
  assign regs_543_io_in = 64'h0; // @[RegFile.scala 75:16:@150682.4]
  assign regs_543_io_reset = reset; // @[RegFile.scala 78:19:@150686.4]
  assign regs_543_io_enable = 1'h1; // @[RegFile.scala 74:20:@150680.4]
  assign regs_544_clock = clock; // @[:@150689.4]
  assign regs_544_reset = io_reset; // @[:@150690.4 RegFile.scala 76:16:@150697.4]
  assign regs_544_io_in = 64'h0; // @[RegFile.scala 75:16:@150696.4]
  assign regs_544_io_reset = reset; // @[RegFile.scala 78:19:@150700.4]
  assign regs_544_io_enable = 1'h1; // @[RegFile.scala 74:20:@150694.4]
  assign regs_545_clock = clock; // @[:@150703.4]
  assign regs_545_reset = io_reset; // @[:@150704.4 RegFile.scala 76:16:@150711.4]
  assign regs_545_io_in = 64'h0; // @[RegFile.scala 75:16:@150710.4]
  assign regs_545_io_reset = reset; // @[RegFile.scala 78:19:@150714.4]
  assign regs_545_io_enable = 1'h1; // @[RegFile.scala 74:20:@150708.4]
  assign regs_546_clock = clock; // @[:@150717.4]
  assign regs_546_reset = io_reset; // @[:@150718.4 RegFile.scala 76:16:@150725.4]
  assign regs_546_io_in = 64'h0; // @[RegFile.scala 75:16:@150724.4]
  assign regs_546_io_reset = reset; // @[RegFile.scala 78:19:@150728.4]
  assign regs_546_io_enable = 1'h1; // @[RegFile.scala 74:20:@150722.4]
  assign regs_547_clock = clock; // @[:@150731.4]
  assign regs_547_reset = io_reset; // @[:@150732.4 RegFile.scala 76:16:@150739.4]
  assign regs_547_io_in = 64'h0; // @[RegFile.scala 75:16:@150738.4]
  assign regs_547_io_reset = reset; // @[RegFile.scala 78:19:@150742.4]
  assign regs_547_io_enable = 1'h1; // @[RegFile.scala 74:20:@150736.4]
  assign regs_548_clock = clock; // @[:@150745.4]
  assign regs_548_reset = io_reset; // @[:@150746.4 RegFile.scala 76:16:@150753.4]
  assign regs_548_io_in = 64'h0; // @[RegFile.scala 75:16:@150752.4]
  assign regs_548_io_reset = reset; // @[RegFile.scala 78:19:@150756.4]
  assign regs_548_io_enable = 1'h1; // @[RegFile.scala 74:20:@150750.4]
  assign regs_549_clock = clock; // @[:@150759.4]
  assign regs_549_reset = io_reset; // @[:@150760.4 RegFile.scala 76:16:@150767.4]
  assign regs_549_io_in = 64'h0; // @[RegFile.scala 75:16:@150766.4]
  assign regs_549_io_reset = reset; // @[RegFile.scala 78:19:@150770.4]
  assign regs_549_io_enable = 1'h1; // @[RegFile.scala 74:20:@150764.4]
  assign regs_550_clock = clock; // @[:@150773.4]
  assign regs_550_reset = io_reset; // @[:@150774.4 RegFile.scala 76:16:@150781.4]
  assign regs_550_io_in = 64'h0; // @[RegFile.scala 75:16:@150780.4]
  assign regs_550_io_reset = reset; // @[RegFile.scala 78:19:@150784.4]
  assign regs_550_io_enable = 1'h1; // @[RegFile.scala 74:20:@150778.4]
  assign regs_551_clock = clock; // @[:@150787.4]
  assign regs_551_reset = io_reset; // @[:@150788.4 RegFile.scala 76:16:@150795.4]
  assign regs_551_io_in = 64'h0; // @[RegFile.scala 75:16:@150794.4]
  assign regs_551_io_reset = reset; // @[RegFile.scala 78:19:@150798.4]
  assign regs_551_io_enable = 1'h1; // @[RegFile.scala 74:20:@150792.4]
  assign regs_552_clock = clock; // @[:@150801.4]
  assign regs_552_reset = io_reset; // @[:@150802.4 RegFile.scala 76:16:@150809.4]
  assign regs_552_io_in = 64'h0; // @[RegFile.scala 75:16:@150808.4]
  assign regs_552_io_reset = reset; // @[RegFile.scala 78:19:@150812.4]
  assign regs_552_io_enable = 1'h1; // @[RegFile.scala 74:20:@150806.4]
  assign regs_553_clock = clock; // @[:@150815.4]
  assign regs_553_reset = io_reset; // @[:@150816.4 RegFile.scala 76:16:@150823.4]
  assign regs_553_io_in = 64'h0; // @[RegFile.scala 75:16:@150822.4]
  assign regs_553_io_reset = reset; // @[RegFile.scala 78:19:@150826.4]
  assign regs_553_io_enable = 1'h1; // @[RegFile.scala 74:20:@150820.4]
  assign regs_554_clock = clock; // @[:@150829.4]
  assign regs_554_reset = io_reset; // @[:@150830.4 RegFile.scala 76:16:@150837.4]
  assign regs_554_io_in = 64'h0; // @[RegFile.scala 75:16:@150836.4]
  assign regs_554_io_reset = reset; // @[RegFile.scala 78:19:@150840.4]
  assign regs_554_io_enable = 1'h1; // @[RegFile.scala 74:20:@150834.4]
  assign regs_555_clock = clock; // @[:@150843.4]
  assign regs_555_reset = io_reset; // @[:@150844.4 RegFile.scala 76:16:@150851.4]
  assign regs_555_io_in = 64'h0; // @[RegFile.scala 75:16:@150850.4]
  assign regs_555_io_reset = reset; // @[RegFile.scala 78:19:@150854.4]
  assign regs_555_io_enable = 1'h1; // @[RegFile.scala 74:20:@150848.4]
  assign regs_556_clock = clock; // @[:@150857.4]
  assign regs_556_reset = io_reset; // @[:@150858.4 RegFile.scala 76:16:@150865.4]
  assign regs_556_io_in = 64'h0; // @[RegFile.scala 75:16:@150864.4]
  assign regs_556_io_reset = reset; // @[RegFile.scala 78:19:@150868.4]
  assign regs_556_io_enable = 1'h1; // @[RegFile.scala 74:20:@150862.4]
  assign regs_557_clock = clock; // @[:@150871.4]
  assign regs_557_reset = io_reset; // @[:@150872.4 RegFile.scala 76:16:@150879.4]
  assign regs_557_io_in = 64'h0; // @[RegFile.scala 75:16:@150878.4]
  assign regs_557_io_reset = reset; // @[RegFile.scala 78:19:@150882.4]
  assign regs_557_io_enable = 1'h1; // @[RegFile.scala 74:20:@150876.4]
  assign regs_558_clock = clock; // @[:@150885.4]
  assign regs_558_reset = io_reset; // @[:@150886.4 RegFile.scala 76:16:@150893.4]
  assign regs_558_io_in = 64'h0; // @[RegFile.scala 75:16:@150892.4]
  assign regs_558_io_reset = reset; // @[RegFile.scala 78:19:@150896.4]
  assign regs_558_io_enable = 1'h1; // @[RegFile.scala 74:20:@150890.4]
  assign regs_559_clock = clock; // @[:@150899.4]
  assign regs_559_reset = io_reset; // @[:@150900.4 RegFile.scala 76:16:@150907.4]
  assign regs_559_io_in = 64'h0; // @[RegFile.scala 75:16:@150906.4]
  assign regs_559_io_reset = reset; // @[RegFile.scala 78:19:@150910.4]
  assign regs_559_io_enable = 1'h1; // @[RegFile.scala 74:20:@150904.4]
  assign regs_560_clock = clock; // @[:@150913.4]
  assign regs_560_reset = io_reset; // @[:@150914.4 RegFile.scala 76:16:@150921.4]
  assign regs_560_io_in = 64'h0; // @[RegFile.scala 75:16:@150920.4]
  assign regs_560_io_reset = reset; // @[RegFile.scala 78:19:@150924.4]
  assign regs_560_io_enable = 1'h1; // @[RegFile.scala 74:20:@150918.4]
  assign regs_561_clock = clock; // @[:@150927.4]
  assign regs_561_reset = io_reset; // @[:@150928.4 RegFile.scala 76:16:@150935.4]
  assign regs_561_io_in = 64'h0; // @[RegFile.scala 75:16:@150934.4]
  assign regs_561_io_reset = reset; // @[RegFile.scala 78:19:@150938.4]
  assign regs_561_io_enable = 1'h1; // @[RegFile.scala 74:20:@150932.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@151506.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@151507.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@151508.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@151509.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@151510.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@151511.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@151512.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@151513.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@151514.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@151515.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@151516.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@151517.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@151518.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@151519.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@151520.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@151521.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@151522.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@151523.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@151524.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@151525.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@151526.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@151527.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@151528.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@151529.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@151530.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@151531.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@151532.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@151533.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@151534.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@151535.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@151536.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@151537.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@151538.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@151539.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@151540.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@151541.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@151542.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@151543.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@151544.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@151545.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@151546.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@151547.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@151548.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@151549.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@151550.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@151551.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@151552.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@151553.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@151554.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@151555.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@151556.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@151557.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@151558.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@151559.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@151560.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@151561.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@151562.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@151563.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@151564.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@151565.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@151566.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@151567.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@151568.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@151569.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@151570.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@151571.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@151572.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@151573.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@151574.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@151575.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@151576.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@151577.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@151578.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@151579.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@151580.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@151581.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@151582.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@151583.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@151584.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@151585.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@151586.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@151587.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@151588.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@151589.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@151590.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@151591.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@151592.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@151593.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@151594.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@151595.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@151596.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@151597.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@151598.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@151599.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@151600.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@151601.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@151602.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@151603.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@151604.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@151605.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@151606.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@151607.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@151608.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@151609.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@151610.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@151611.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@151612.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@151613.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@151614.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@151615.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@151616.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@151617.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@151618.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@151619.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@151620.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@151621.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@151622.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@151623.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@151624.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@151625.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@151626.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@151627.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@151628.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@151629.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@151630.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@151631.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@151632.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@151633.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@151634.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@151635.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@151636.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@151637.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@151638.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@151639.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@151640.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@151641.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@151642.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@151643.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@151644.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@151645.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@151646.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@151647.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@151648.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@151649.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@151650.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@151651.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@151652.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@151653.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@151654.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@151655.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@151656.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@151657.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@151658.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@151659.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@151660.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@151661.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@151662.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@151663.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@151664.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@151665.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@151666.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@151667.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@151668.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@151669.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@151670.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@151671.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@151672.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@151673.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@151674.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@151675.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@151676.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@151677.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@151678.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@151679.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@151680.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@151681.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@151682.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@151683.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@151684.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@151685.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@151686.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@151687.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@151688.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@151689.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@151690.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@151691.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@151692.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@151693.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@151694.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@151695.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@151696.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@151697.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@151698.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@151699.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@151700.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@151701.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@151702.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@151703.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@151704.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@151705.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@151706.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@151707.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@151708.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@151709.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@151710.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@151711.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@151712.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@151713.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@151714.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@151715.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@151716.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@151717.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@151718.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@151719.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@151720.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@151721.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@151722.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@151723.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@151724.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@151725.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@151726.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@151727.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@151728.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@151729.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@151730.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@151731.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@151732.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@151733.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@151734.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@151735.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@151736.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@151737.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@151738.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@151739.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@151740.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@151741.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@151742.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@151743.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@151744.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@151745.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@151746.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@151747.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@151748.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@151749.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@151750.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@151751.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@151752.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@151753.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@151754.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@151755.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@151756.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@151757.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@151758.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@151759.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@151760.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@151761.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@151762.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@151763.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@151764.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@151765.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@151766.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@151767.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@151768.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@151769.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@151770.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@151771.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@151772.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@151773.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@151774.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@151775.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@151776.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@151777.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@151778.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@151779.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@151780.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@151781.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@151782.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@151783.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@151784.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@151785.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@151786.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@151787.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@151788.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@151789.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@151790.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@151791.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@151792.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@151793.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@151794.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@151795.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@151796.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@151797.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@151798.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@151799.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@151800.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@151801.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@151802.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@151803.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@151804.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@151805.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@151806.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@151807.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@151808.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@151809.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@151810.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@151811.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@151812.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@151813.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@151814.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@151815.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@151816.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@151817.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@151818.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@151819.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@151820.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@151821.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@151822.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@151823.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@151824.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@151825.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@151826.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@151827.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@151828.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@151829.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@151830.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@151831.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@151832.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@151833.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@151834.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@151835.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@151836.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@151837.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@151838.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@151839.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@151840.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@151841.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@151842.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@151843.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@151844.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@151845.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@151846.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@151847.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@151848.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@151849.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@151850.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@151851.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@151852.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@151853.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@151854.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@151855.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@151856.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@151857.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@151858.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@151859.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@151860.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@151861.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@151862.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@151863.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@151864.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@151865.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@151866.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@151867.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@151868.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@151869.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@151870.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@151871.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@151872.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@151873.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@151874.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@151875.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@151876.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@151877.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@151878.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@151879.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@151880.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@151881.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@151882.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@151883.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@151884.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@151885.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@151886.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@151887.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@151888.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@151889.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@151890.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@151891.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@151892.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@151893.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@151894.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@151895.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@151896.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@151897.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@151898.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@151899.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@151900.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@151901.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@151902.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@151903.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@151904.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@151905.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@151906.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@151907.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@151908.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@151909.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@151910.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@151911.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@151912.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@151913.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@151914.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@151915.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@151916.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@151917.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@151918.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@151919.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@151920.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@151921.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@151922.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@151923.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@151924.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@151925.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@151926.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@151927.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@151928.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@151929.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@151930.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@151931.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@151932.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@151933.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@151934.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@151935.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@151936.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@151937.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@151938.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@151939.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@151940.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@151941.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@151942.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@151943.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@151944.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@151945.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@151946.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@151947.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@151948.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@151949.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@151950.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@151951.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@151952.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@151953.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@151954.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@151955.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@151956.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@151957.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@151958.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@151959.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@151960.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@151961.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@151962.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@151963.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@151964.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@151965.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@151966.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@151967.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@151968.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@151969.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@151970.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@151971.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@151972.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@151973.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@151974.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@151975.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@151976.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@151977.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@151978.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@151979.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@151980.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@151981.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@151982.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@151983.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@151984.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@151985.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@151986.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@151987.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@151988.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@151989.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@151990.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@151991.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@151992.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@151993.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@151994.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@151995.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@151996.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@151997.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@151998.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@151999.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@152000.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@152001.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@152002.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@152003.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@152004.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@152005.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@152006.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@152007.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@152008.4]
  assign rport_io_ins_503 = regs_503_io_out; // @[RegFile.scala 97:16:@152009.4]
  assign rport_io_ins_504 = regs_504_io_out; // @[RegFile.scala 97:16:@152010.4]
  assign rport_io_ins_505 = regs_505_io_out; // @[RegFile.scala 97:16:@152011.4]
  assign rport_io_ins_506 = regs_506_io_out; // @[RegFile.scala 97:16:@152012.4]
  assign rport_io_ins_507 = regs_507_io_out; // @[RegFile.scala 97:16:@152013.4]
  assign rport_io_ins_508 = regs_508_io_out; // @[RegFile.scala 97:16:@152014.4]
  assign rport_io_ins_509 = regs_509_io_out; // @[RegFile.scala 97:16:@152015.4]
  assign rport_io_ins_510 = regs_510_io_out; // @[RegFile.scala 97:16:@152016.4]
  assign rport_io_ins_511 = regs_511_io_out; // @[RegFile.scala 97:16:@152017.4]
  assign rport_io_ins_512 = regs_512_io_out; // @[RegFile.scala 97:16:@152018.4]
  assign rport_io_ins_513 = regs_513_io_out; // @[RegFile.scala 97:16:@152019.4]
  assign rport_io_ins_514 = regs_514_io_out; // @[RegFile.scala 97:16:@152020.4]
  assign rport_io_ins_515 = regs_515_io_out; // @[RegFile.scala 97:16:@152021.4]
  assign rport_io_ins_516 = regs_516_io_out; // @[RegFile.scala 97:16:@152022.4]
  assign rport_io_ins_517 = regs_517_io_out; // @[RegFile.scala 97:16:@152023.4]
  assign rport_io_ins_518 = regs_518_io_out; // @[RegFile.scala 97:16:@152024.4]
  assign rport_io_ins_519 = regs_519_io_out; // @[RegFile.scala 97:16:@152025.4]
  assign rport_io_ins_520 = regs_520_io_out; // @[RegFile.scala 97:16:@152026.4]
  assign rport_io_ins_521 = regs_521_io_out; // @[RegFile.scala 97:16:@152027.4]
  assign rport_io_ins_522 = regs_522_io_out; // @[RegFile.scala 97:16:@152028.4]
  assign rport_io_ins_523 = regs_523_io_out; // @[RegFile.scala 97:16:@152029.4]
  assign rport_io_ins_524 = regs_524_io_out; // @[RegFile.scala 97:16:@152030.4]
  assign rport_io_ins_525 = regs_525_io_out; // @[RegFile.scala 97:16:@152031.4]
  assign rport_io_ins_526 = regs_526_io_out; // @[RegFile.scala 97:16:@152032.4]
  assign rport_io_ins_527 = regs_527_io_out; // @[RegFile.scala 97:16:@152033.4]
  assign rport_io_ins_528 = regs_528_io_out; // @[RegFile.scala 97:16:@152034.4]
  assign rport_io_ins_529 = regs_529_io_out; // @[RegFile.scala 97:16:@152035.4]
  assign rport_io_ins_530 = regs_530_io_out; // @[RegFile.scala 97:16:@152036.4]
  assign rport_io_ins_531 = regs_531_io_out; // @[RegFile.scala 97:16:@152037.4]
  assign rport_io_ins_532 = regs_532_io_out; // @[RegFile.scala 97:16:@152038.4]
  assign rport_io_ins_533 = regs_533_io_out; // @[RegFile.scala 97:16:@152039.4]
  assign rport_io_ins_534 = regs_534_io_out; // @[RegFile.scala 97:16:@152040.4]
  assign rport_io_ins_535 = regs_535_io_out; // @[RegFile.scala 97:16:@152041.4]
  assign rport_io_ins_536 = regs_536_io_out; // @[RegFile.scala 97:16:@152042.4]
  assign rport_io_ins_537 = regs_537_io_out; // @[RegFile.scala 97:16:@152043.4]
  assign rport_io_ins_538 = regs_538_io_out; // @[RegFile.scala 97:16:@152044.4]
  assign rport_io_ins_539 = regs_539_io_out; // @[RegFile.scala 97:16:@152045.4]
  assign rport_io_ins_540 = regs_540_io_out; // @[RegFile.scala 97:16:@152046.4]
  assign rport_io_ins_541 = regs_541_io_out; // @[RegFile.scala 97:16:@152047.4]
  assign rport_io_ins_542 = regs_542_io_out; // @[RegFile.scala 97:16:@152048.4]
  assign rport_io_ins_543 = regs_543_io_out; // @[RegFile.scala 97:16:@152049.4]
  assign rport_io_ins_544 = regs_544_io_out; // @[RegFile.scala 97:16:@152050.4]
  assign rport_io_ins_545 = regs_545_io_out; // @[RegFile.scala 97:16:@152051.4]
  assign rport_io_ins_546 = regs_546_io_out; // @[RegFile.scala 97:16:@152052.4]
  assign rport_io_ins_547 = regs_547_io_out; // @[RegFile.scala 97:16:@152053.4]
  assign rport_io_ins_548 = regs_548_io_out; // @[RegFile.scala 97:16:@152054.4]
  assign rport_io_ins_549 = regs_549_io_out; // @[RegFile.scala 97:16:@152055.4]
  assign rport_io_ins_550 = regs_550_io_out; // @[RegFile.scala 97:16:@152056.4]
  assign rport_io_ins_551 = regs_551_io_out; // @[RegFile.scala 97:16:@152057.4]
  assign rport_io_ins_552 = regs_552_io_out; // @[RegFile.scala 97:16:@152058.4]
  assign rport_io_ins_553 = regs_553_io_out; // @[RegFile.scala 97:16:@152059.4]
  assign rport_io_ins_554 = regs_554_io_out; // @[RegFile.scala 97:16:@152060.4]
  assign rport_io_ins_555 = regs_555_io_out; // @[RegFile.scala 97:16:@152061.4]
  assign rport_io_ins_556 = regs_556_io_out; // @[RegFile.scala 97:16:@152062.4]
  assign rport_io_ins_557 = regs_557_io_out; // @[RegFile.scala 97:16:@152063.4]
  assign rport_io_ins_558 = regs_558_io_out; // @[RegFile.scala 97:16:@152064.4]
  assign rport_io_ins_559 = regs_559_io_out; // @[RegFile.scala 97:16:@152065.4]
  assign rport_io_ins_560 = regs_560_io_out; // @[RegFile.scala 97:16:@152066.4]
  assign rport_io_ins_561 = regs_561_io_out; // @[RegFile.scala 97:16:@152067.4]
  assign rport_io_sel = io_raddr[9:0]; // @[RegFile.scala 106:18:@152068.4]
endmodule
module RetimeWrapper_1374( // @[:@152092.2]
  input         clock, // @[:@152093.4]
  input         reset, // @[:@152094.4]
  input  [39:0] io_in, // @[:@152095.4]
  output [39:0] io_out // @[:@152095.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@152097.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@152097.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@152097.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@152097.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@152097.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@152097.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@152097.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@152110.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@152109.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@152108.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@152107.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@152106.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@152104.4]
endmodule
module FringeFF_562( // @[:@152112.2]
  input         clock, // @[:@152113.4]
  input         reset, // @[:@152114.4]
  input  [39:0] io_in, // @[:@152115.4]
  output [39:0] io_out, // @[:@152115.4]
  input         io_enable // @[:@152115.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@152118.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@152118.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@152118.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@152118.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@152123.4 package.scala 96:25:@152124.4]
  RetimeWrapper_1374 RetimeWrapper ( // @[package.scala 93:22:@152118.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@152123.4 package.scala 96:25:@152124.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@152135.4]
  assign RetimeWrapper_clock = clock; // @[:@152119.4]
  assign RetimeWrapper_reset = reset; // @[:@152120.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@152121.4]
endmodule
module FringeCounter( // @[:@152137.2]
  input   clock, // @[:@152138.4]
  input   reset, // @[:@152139.4]
  input   io_enable, // @[:@152140.4]
  output  io_done // @[:@152140.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@152142.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@152142.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@152142.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@152142.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@152142.4]
  wire [40:0] count; // @[Cat.scala 30:58:@152149.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@152150.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@152151.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@152152.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@152154.4]
  FringeFF_562 reg$ ( // @[FringeCounter.scala 24:19:@152142.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@152149.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@152150.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@152151.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@152152.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@152154.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@152165.4]
  assign reg$_clock = clock; // @[:@152143.4]
  assign reg$_reset = reset; // @[:@152144.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@152156.6 FringeCounter.scala 37:15:@152159.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@152147.4]
endmodule
module FringeFF_563( // @[:@152199.2]
  input   clock, // @[:@152200.4]
  input   reset, // @[:@152201.4]
  input   io_in, // @[:@152202.4]
  input   io_reset, // @[:@152202.4]
  output  io_out, // @[:@152202.4]
  input   io_enable // @[:@152202.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@152205.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@152205.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@152205.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@152205.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@152205.4]
  wire  _T_18; // @[package.scala 96:25:@152210.4 package.scala 96:25:@152211.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@152216.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@152205.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@152210.4 package.scala 96:25:@152211.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@152216.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@152222.4]
  assign RetimeWrapper_clock = clock; // @[:@152206.4]
  assign RetimeWrapper_reset = reset; // @[:@152207.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@152209.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@152208.4]
endmodule
module Depulser( // @[:@152224.2]
  input   clock, // @[:@152225.4]
  input   reset, // @[:@152226.4]
  input   io_in, // @[:@152227.4]
  input   io_rst, // @[:@152227.4]
  output  io_out // @[:@152227.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@152229.4]
  wire  r_reset; // @[Depulser.scala 14:17:@152229.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@152229.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@152229.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@152229.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@152229.4]
  FringeFF_563 r ( // @[Depulser.scala 14:17:@152229.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@152238.4]
  assign r_clock = clock; // @[:@152230.4]
  assign r_reset = reset; // @[:@152231.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@152233.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@152237.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@152236.4]
endmodule
module Fringe( // @[:@152240.2]
  input         clock, // @[:@152241.4]
  input         reset, // @[:@152242.4]
  input  [31:0] io_raddr, // @[:@152243.4]
  input         io_wen, // @[:@152243.4]
  input  [31:0] io_waddr, // @[:@152243.4]
  input  [63:0] io_wdata, // @[:@152243.4]
  output [63:0] io_rdata, // @[:@152243.4]
  output        io_enable, // @[:@152243.4]
  input         io_done, // @[:@152243.4]
  output        io_reset, // @[:@152243.4]
  output [63:0] io_argIns_0, // @[:@152243.4]
  output [63:0] io_argIns_1, // @[:@152243.4]
  input         io_argOuts_0_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_0_bits, // @[:@152243.4]
  input         io_argOuts_1_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_1_bits, // @[:@152243.4]
  input         io_argOuts_2_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_2_bits, // @[:@152243.4]
  input         io_argOuts_3_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_3_bits, // @[:@152243.4]
  input         io_argOuts_4_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_4_bits, // @[:@152243.4]
  input         io_argOuts_5_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_5_bits, // @[:@152243.4]
  input         io_argOuts_6_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_6_bits, // @[:@152243.4]
  input         io_argOuts_7_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_7_bits, // @[:@152243.4]
  input         io_argOuts_8_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_8_bits, // @[:@152243.4]
  input         io_argOuts_9_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_9_bits, // @[:@152243.4]
  input         io_argOuts_10_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_10_bits, // @[:@152243.4]
  input         io_argOuts_11_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_11_bits, // @[:@152243.4]
  input         io_argOuts_12_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_12_bits, // @[:@152243.4]
  input         io_argOuts_13_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_13_bits, // @[:@152243.4]
  input         io_argOuts_14_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_14_bits, // @[:@152243.4]
  input         io_argOuts_15_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_15_bits, // @[:@152243.4]
  input         io_argOuts_16_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_16_bits, // @[:@152243.4]
  input         io_argOuts_17_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_17_bits, // @[:@152243.4]
  input         io_argOuts_18_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_18_bits, // @[:@152243.4]
  input         io_argOuts_19_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_19_bits, // @[:@152243.4]
  input         io_argOuts_20_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_20_bits, // @[:@152243.4]
  input         io_argOuts_21_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_21_bits, // @[:@152243.4]
  input         io_argOuts_22_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_22_bits, // @[:@152243.4]
  input         io_argOuts_23_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_23_bits, // @[:@152243.4]
  input         io_argOuts_24_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_24_bits, // @[:@152243.4]
  input         io_argOuts_25_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_25_bits, // @[:@152243.4]
  input         io_argOuts_26_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_26_bits, // @[:@152243.4]
  input         io_argOuts_27_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_27_bits, // @[:@152243.4]
  input         io_argOuts_28_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_28_bits, // @[:@152243.4]
  input         io_argOuts_29_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_29_bits, // @[:@152243.4]
  input         io_argOuts_30_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_30_bits, // @[:@152243.4]
  input         io_argOuts_31_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_31_bits, // @[:@152243.4]
  input         io_argOuts_32_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_32_bits, // @[:@152243.4]
  input         io_argOuts_33_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_33_bits, // @[:@152243.4]
  input         io_argOuts_34_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_34_bits, // @[:@152243.4]
  input         io_argOuts_35_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_35_bits, // @[:@152243.4]
  input         io_argOuts_36_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_36_bits, // @[:@152243.4]
  input         io_argOuts_37_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_37_bits, // @[:@152243.4]
  input         io_argOuts_38_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_38_bits, // @[:@152243.4]
  input         io_argOuts_39_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_39_bits, // @[:@152243.4]
  input         io_argOuts_40_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_40_bits, // @[:@152243.4]
  input         io_argOuts_41_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_41_bits, // @[:@152243.4]
  input         io_argOuts_42_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_42_bits, // @[:@152243.4]
  input         io_argOuts_43_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_43_bits, // @[:@152243.4]
  input         io_argOuts_44_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_44_bits, // @[:@152243.4]
  input         io_argOuts_45_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_45_bits, // @[:@152243.4]
  input         io_argOuts_46_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_46_bits, // @[:@152243.4]
  input         io_argOuts_47_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_47_bits, // @[:@152243.4]
  input         io_argOuts_48_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_48_bits, // @[:@152243.4]
  input         io_argOuts_49_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_49_bits, // @[:@152243.4]
  input         io_argOuts_50_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_50_bits, // @[:@152243.4]
  input         io_argOuts_51_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_51_bits, // @[:@152243.4]
  input         io_argOuts_52_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_52_bits, // @[:@152243.4]
  input         io_argOuts_53_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_53_bits, // @[:@152243.4]
  input         io_argOuts_54_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_54_bits, // @[:@152243.4]
  input         io_argOuts_55_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_55_bits, // @[:@152243.4]
  input         io_argOuts_56_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_56_bits, // @[:@152243.4]
  input         io_argOuts_57_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_57_bits, // @[:@152243.4]
  input         io_argOuts_58_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_58_bits, // @[:@152243.4]
  input         io_argOuts_59_valid, // @[:@152243.4]
  input  [63:0] io_argOuts_59_bits, // @[:@152243.4]
  output [63:0] io_argEchos_0, // @[:@152243.4]
  output [63:0] io_argEchos_1, // @[:@152243.4]
  output [63:0] io_argEchos_2, // @[:@152243.4]
  output [63:0] io_argEchos_3, // @[:@152243.4]
  output [63:0] io_argEchos_4, // @[:@152243.4]
  output [63:0] io_argEchos_5, // @[:@152243.4]
  output [63:0] io_argEchos_6, // @[:@152243.4]
  output [63:0] io_argEchos_7, // @[:@152243.4]
  output [63:0] io_argEchos_8, // @[:@152243.4]
  output [63:0] io_argEchos_9, // @[:@152243.4]
  output [63:0] io_argEchos_10, // @[:@152243.4]
  output [63:0] io_argEchos_11, // @[:@152243.4]
  output [63:0] io_argEchos_12, // @[:@152243.4]
  output [63:0] io_argEchos_13, // @[:@152243.4]
  output [63:0] io_argEchos_14, // @[:@152243.4]
  output [63:0] io_argEchos_15, // @[:@152243.4]
  output [63:0] io_argEchos_16, // @[:@152243.4]
  output [63:0] io_argEchos_17, // @[:@152243.4]
  output [63:0] io_argEchos_18, // @[:@152243.4]
  output [63:0] io_argEchos_19, // @[:@152243.4]
  output [63:0] io_argEchos_20, // @[:@152243.4]
  output [63:0] io_argEchos_21, // @[:@152243.4]
  output [63:0] io_argEchos_22, // @[:@152243.4]
  output [63:0] io_argEchos_23, // @[:@152243.4]
  output [63:0] io_argEchos_24, // @[:@152243.4]
  output [63:0] io_argEchos_25, // @[:@152243.4]
  output [63:0] io_argEchos_26, // @[:@152243.4]
  output [63:0] io_argEchos_27, // @[:@152243.4]
  output [63:0] io_argEchos_28, // @[:@152243.4]
  output [63:0] io_argEchos_29, // @[:@152243.4]
  output [63:0] io_argEchos_30, // @[:@152243.4]
  output [63:0] io_argEchos_31, // @[:@152243.4]
  output [63:0] io_argEchos_32, // @[:@152243.4]
  output [63:0] io_argEchos_33, // @[:@152243.4]
  output [63:0] io_argEchos_34, // @[:@152243.4]
  output [63:0] io_argEchos_35, // @[:@152243.4]
  output [63:0] io_argEchos_36, // @[:@152243.4]
  output [63:0] io_argEchos_37, // @[:@152243.4]
  output [63:0] io_argEchos_38, // @[:@152243.4]
  output [63:0] io_argEchos_39, // @[:@152243.4]
  output [63:0] io_argEchos_40, // @[:@152243.4]
  output [63:0] io_argEchos_41, // @[:@152243.4]
  output [63:0] io_argEchos_42, // @[:@152243.4]
  output [63:0] io_argEchos_43, // @[:@152243.4]
  output [63:0] io_argEchos_44, // @[:@152243.4]
  output [63:0] io_argEchos_45, // @[:@152243.4]
  output [63:0] io_argEchos_46, // @[:@152243.4]
  output [63:0] io_argEchos_47, // @[:@152243.4]
  output [63:0] io_argEchos_48, // @[:@152243.4]
  output [63:0] io_argEchos_49, // @[:@152243.4]
  output [63:0] io_argEchos_50, // @[:@152243.4]
  output [63:0] io_argEchos_51, // @[:@152243.4]
  output [63:0] io_argEchos_52, // @[:@152243.4]
  output [63:0] io_argEchos_53, // @[:@152243.4]
  output [63:0] io_argEchos_54, // @[:@152243.4]
  output [63:0] io_argEchos_55, // @[:@152243.4]
  output [63:0] io_argEchos_56, // @[:@152243.4]
  output [63:0] io_argEchos_57, // @[:@152243.4]
  output [63:0] io_argEchos_58, // @[:@152243.4]
  output [63:0] io_argEchos_59, // @[:@152243.4]
  output        io_memStreams_loads_0_cmd_ready, // @[:@152243.4]
  input         io_memStreams_loads_0_cmd_valid, // @[:@152243.4]
  input  [63:0] io_memStreams_loads_0_cmd_bits_addr, // @[:@152243.4]
  input  [31:0] io_memStreams_loads_0_cmd_bits_size, // @[:@152243.4]
  input         io_memStreams_loads_0_data_ready, // @[:@152243.4]
  output        io_memStreams_loads_0_data_valid, // @[:@152243.4]
  output [31:0] io_memStreams_loads_0_data_bits_rdata_0, // @[:@152243.4]
  output        io_memStreams_stores_0_cmd_ready, // @[:@152243.4]
  input         io_memStreams_stores_0_cmd_valid, // @[:@152243.4]
  input  [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@152243.4]
  input  [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@152243.4]
  output        io_memStreams_stores_0_data_ready, // @[:@152243.4]
  input         io_memStreams_stores_0_data_valid, // @[:@152243.4]
  input  [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@152243.4]
  input         io_memStreams_stores_0_data_bits_wstrb, // @[:@152243.4]
  input         io_memStreams_stores_0_wresp_ready, // @[:@152243.4]
  output        io_memStreams_stores_0_wresp_valid, // @[:@152243.4]
  output        io_memStreams_stores_0_wresp_bits, // @[:@152243.4]
  input         io_dram_0_cmd_ready, // @[:@152243.4]
  output        io_dram_0_cmd_valid, // @[:@152243.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@152243.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@152243.4]
  output [63:0] io_dram_0_cmd_bits_rawAddr, // @[:@152243.4]
  output        io_dram_0_cmd_bits_isWr, // @[:@152243.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@152243.4]
  input         io_dram_0_wdata_ready, // @[:@152243.4]
  output        io_dram_0_wdata_valid, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_0, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_1, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_2, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_3, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_4, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_5, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_6, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_7, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_8, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_9, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_10, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_11, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_12, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_13, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_14, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_15, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_16, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_17, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_18, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_19, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_20, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_21, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_22, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_23, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_24, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_25, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_26, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_27, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_28, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_29, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_30, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_31, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_32, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_33, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_34, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_35, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_36, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_37, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_38, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_39, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_40, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_41, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_42, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_43, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_44, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_45, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_46, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_47, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_48, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_49, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_50, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_51, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_52, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_53, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_54, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_55, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_56, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_57, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_58, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_59, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_60, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_61, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_62, // @[:@152243.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_63, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_0, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_1, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_2, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_3, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_4, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_5, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_6, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_7, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_8, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_9, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_10, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_11, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_12, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_13, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_14, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_15, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_16, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_17, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_18, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_19, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_20, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_21, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_22, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_23, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_24, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_25, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_26, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_27, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_28, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_29, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_30, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_31, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_32, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_33, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_34, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_35, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_36, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_37, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_38, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_39, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_40, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_41, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_42, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_43, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_44, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_45, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_46, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_47, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_48, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_49, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_50, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_51, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_52, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_53, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_54, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_55, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_56, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_57, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_58, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_59, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_60, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_61, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_62, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wstrb_63, // @[:@152243.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@152243.4]
  output        io_dram_0_rresp_ready, // @[:@152243.4]
  input         io_dram_0_rresp_valid, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_0, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_1, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_2, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_3, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_4, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_5, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_6, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_7, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_8, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_9, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_10, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_11, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_12, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_13, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_14, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_15, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_16, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_17, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_18, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_19, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_20, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_21, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_22, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_23, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_24, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_25, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_26, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_27, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_28, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_29, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_30, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_31, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_32, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_33, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_34, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_35, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_36, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_37, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_38, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_39, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_40, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_41, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_42, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_43, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_44, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_45, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_46, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_47, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_48, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_49, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_50, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_51, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_52, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_53, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_54, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_55, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_56, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_57, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_58, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_59, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_60, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_61, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_62, // @[:@152243.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_63, // @[:@152243.4]
  input  [31:0] io_dram_0_rresp_bits_tag, // @[:@152243.4]
  output        io_dram_0_wresp_ready, // @[:@152243.4]
  input         io_dram_0_wresp_valid, // @[:@152243.4]
  input  [31:0] io_dram_0_wresp_bits_tag, // @[:@152243.4]
  input         io_heap_0_req_valid, // @[:@152243.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@152243.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@152243.4]
  output        io_heap_0_resp_valid, // @[:@152243.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@152243.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@152243.4]
);
  wire  dramArbs_0_clock; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_reset; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_enable; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_app_loads_0_cmd_ready; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_app_loads_0_cmd_valid; // @[Fringe.scala 91:25:@152485.4]
  wire [63:0] dramArbs_0_io_app_loads_0_cmd_bits_addr; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_app_loads_0_cmd_bits_size; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_app_loads_0_data_ready; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_app_loads_0_data_valid; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_app_loads_0_data_bits_rdata_0; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_app_stores_0_cmd_valid; // @[Fringe.scala 91:25:@152485.4]
  wire [63:0] dramArbs_0_io_app_stores_0_cmd_bits_addr; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_app_stores_0_cmd_bits_size; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_app_stores_0_data_valid; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_app_stores_0_data_bits_wdata_0; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_app_stores_0_data_bits_wstrb; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_app_stores_0_wresp_ready; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_cmd_ready; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 91:25:@152485.4]
  wire [63:0] dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@152485.4]
  wire [63:0] dramArbs_0_io_dram_cmd_bits_rawAddr; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_ready; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_16; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_17; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_18; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_19; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_20; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_21; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_22; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_23; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_24; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_25; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_26; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_27; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_28; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_29; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_30; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_31; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_32; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_33; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_34; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_35; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_36; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_37; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_38; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_39; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_40; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_41; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_42; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_43; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_44; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_45; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_46; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_47; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_48; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_49; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_50; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_51; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_52; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_53; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_54; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_55; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_56; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_57; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_58; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_59; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_60; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_61; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_62; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_wdata_bits_wdata_63; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_rresp_valid; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_0; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_1; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_2; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_3; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_4; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_5; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_6; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_7; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_8; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_9; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_10; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_11; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_12; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_13; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_14; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_15; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_16; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_17; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_18; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_19; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_20; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_21; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_22; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_23; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_24; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_25; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_26; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_27; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_28; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_29; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_30; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_31; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_32; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_33; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_34; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_35; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_36; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_37; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_38; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_39; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_40; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_41; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_42; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_43; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_44; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_45; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_46; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_47; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_48; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_49; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_50; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_51; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_52; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_53; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_54; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_55; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_56; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_57; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_58; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_59; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_60; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_61; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_62; // @[Fringe.scala 91:25:@152485.4]
  wire [7:0] dramArbs_0_io_dram_rresp_bits_rdata_63; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_tag; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 91:25:@152485.4]
  wire  dramArbs_0_io_dram_wresp_valid; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_0; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_1; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_2; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_3; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_4; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_5; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_6; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_7; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_8; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_9; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_10; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_11; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_12; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_13; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_14; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_15; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_16; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_17; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_18; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_19; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_20; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_21; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_22; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_23; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_24; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_25; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_26; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_27; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_28; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_29; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_30; // @[Fringe.scala 91:25:@152485.4]
  wire [31:0] dramArbs_0_io_debugSignals_41; // @[Fringe.scala 91:25:@152485.4]
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@153928.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@153928.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@153928.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@153928.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@153928.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@153928.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@153928.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@153928.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@153928.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@153928.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@153928.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@153928.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@153937.4]
  wire [10:0] regs_io_raddr; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@153937.4]
  wire [10:0] regs_io_waddr; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argIns_3; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_2_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_2_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_3_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_3_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_4_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_4_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_5_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_5_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_6_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_6_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_7_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_7_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_8_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_8_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_9_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_9_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_10_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_10_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_11_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_11_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_12_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_12_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_13_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_13_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_14_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_14_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_15_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_15_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_16_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_16_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_17_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_17_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_18_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_18_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_19_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_19_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_20_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_20_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_21_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_21_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_22_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_22_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_23_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_23_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_24_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_24_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_25_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_25_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_26_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_26_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_27_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_27_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_28_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_28_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_29_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_29_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_30_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_30_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_31_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_31_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_32_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_32_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_33_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_33_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_34_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_34_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_35_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_35_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_36_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_36_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_37_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_37_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_38_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_38_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_39_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_39_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_40_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_40_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_41_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_41_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_42_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_42_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_43_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_43_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_44_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_44_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_45_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_45_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_46_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_46_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_47_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_47_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_48_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_48_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_49_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_49_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_50_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_50_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_51_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_51_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_52_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_52_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_53_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_53_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_54_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_54_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_55_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_55_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_56_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_56_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_57_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_57_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_58_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_58_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_59_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_59_bits; // @[Fringe.scala 116:20:@153937.4]
  wire  regs_io_argOuts_60_valid; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_60_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_61_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_62_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_63_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_64_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_65_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_66_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_67_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_68_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_69_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_70_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_71_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_72_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_73_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_74_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_75_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_76_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_77_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_78_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_79_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_80_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_81_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_82_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_83_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_84_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_85_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_86_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_87_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_88_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_89_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_90_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_91_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argOuts_102_bits; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_1; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_2; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_3; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_4; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_5; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_6; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_7; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_8; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_9; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_10; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_11; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_12; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_13; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_14; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_15; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_16; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_17; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_18; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_19; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_20; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_21; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_22; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_23; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_24; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_25; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_26; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_27; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_28; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_29; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_30; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_31; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_32; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_33; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_34; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_35; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_36; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_37; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_38; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_39; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_40; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_41; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_42; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_43; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_44; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_45; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_46; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_47; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_48; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_49; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_50; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_51; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_52; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_53; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_54; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_55; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_56; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_57; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_58; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_59; // @[Fringe.scala 116:20:@153937.4]
  wire [63:0] regs_io_argEchos_60; // @[Fringe.scala 116:20:@153937.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@156227.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@156227.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@156227.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@156227.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@156246.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@156246.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@156246.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@156246.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@156246.4]
  reg [63:0] _T_949; // @[Reg.scala 11:16:@156198.4]
  reg [63:0] _RAND_0;
  wire [63:0] _T_953; // @[:@156204.4 :@156205.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@156206.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@156208.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@156210.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@156212.4]
  wire  _T_958; // @[Fringe.scala 134:60:@156214.4]
  wire  _T_962; // @[Fringe.scala 134:74:@156216.4]
  wire  _T_963; // @[Fringe.scala 135:27:@156218.4]
  wire [63:0] _T_973; // @[Fringe.scala 156:22:@156254.4]
  reg  _T_980; // @[package.scala 152:20:@156257.4]
  reg [31:0] _RAND_1;
  wire  _T_981; // @[package.scala 153:13:@156259.4]
  wire  _T_982; // @[package.scala 153:8:@156260.4]
  wire  _T_985; // @[Fringe.scala 160:55:@156264.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@156265.4]
  wire  _T_988; // @[Fringe.scala 161:58:@156268.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@156269.4]
  wire [1:0] _T_992; // @[Fringe.scala 162:57:@156271.4]
  wire [1:0] _T_994; // @[Fringe.scala 162:34:@156272.4]
  wire [63:0] _T_996; // @[Fringe.scala 163:30:@156274.4]
  wire [1:0] _T_997; // @[Fringe.scala 171:37:@156277.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@156256.4 Fringe.scala 163:24:@156275.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@156256.4 Fringe.scala 162:28:@156273.4]
  wire [61:0] _T_998; // @[Fringe.scala 171:37:@156278.4]
  wire  alloc; // @[Fringe.scala 202:38:@157672.4]
  wire  dealloc; // @[Fringe.scala 203:40:@157673.4]
  wire  _T_1502; // @[Fringe.scala 204:37:@157674.4]
  reg  _T_1505; // @[package.scala 152:20:@157675.4]
  reg [31:0] _RAND_2;
  wire  _T_1506; // @[package.scala 153:13:@157677.4]
  DRAMArbiter dramArbs_0 ( // @[Fringe.scala 91:25:@152485.4]
    .clock(dramArbs_0_clock),
    .reset(dramArbs_0_reset),
    .io_enable(dramArbs_0_io_enable),
    .io_app_loads_0_cmd_ready(dramArbs_0_io_app_loads_0_cmd_ready),
    .io_app_loads_0_cmd_valid(dramArbs_0_io_app_loads_0_cmd_valid),
    .io_app_loads_0_cmd_bits_addr(dramArbs_0_io_app_loads_0_cmd_bits_addr),
    .io_app_loads_0_cmd_bits_size(dramArbs_0_io_app_loads_0_cmd_bits_size),
    .io_app_loads_0_data_ready(dramArbs_0_io_app_loads_0_data_ready),
    .io_app_loads_0_data_valid(dramArbs_0_io_app_loads_0_data_valid),
    .io_app_loads_0_data_bits_rdata_0(dramArbs_0_io_app_loads_0_data_bits_rdata_0),
    .io_app_stores_0_cmd_ready(dramArbs_0_io_app_stores_0_cmd_ready),
    .io_app_stores_0_cmd_valid(dramArbs_0_io_app_stores_0_cmd_valid),
    .io_app_stores_0_cmd_bits_addr(dramArbs_0_io_app_stores_0_cmd_bits_addr),
    .io_app_stores_0_cmd_bits_size(dramArbs_0_io_app_stores_0_cmd_bits_size),
    .io_app_stores_0_data_ready(dramArbs_0_io_app_stores_0_data_ready),
    .io_app_stores_0_data_valid(dramArbs_0_io_app_stores_0_data_valid),
    .io_app_stores_0_data_bits_wdata_0(dramArbs_0_io_app_stores_0_data_bits_wdata_0),
    .io_app_stores_0_data_bits_wstrb(dramArbs_0_io_app_stores_0_data_bits_wstrb),
    .io_app_stores_0_wresp_ready(dramArbs_0_io_app_stores_0_wresp_ready),
    .io_app_stores_0_wresp_valid(dramArbs_0_io_app_stores_0_wresp_valid),
    .io_app_stores_0_wresp_bits(dramArbs_0_io_app_stores_0_wresp_bits),
    .io_dram_cmd_ready(dramArbs_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_rawAddr(dramArbs_0_io_dram_cmd_bits_rawAddr),
    .io_dram_cmd_bits_isWr(dramArbs_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_0_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_0_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_0_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_0_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_0_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_0_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_0_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_0_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_0_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_0_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_0_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_0_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_0_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_0_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_0_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_0_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wdata_16(dramArbs_0_io_dram_wdata_bits_wdata_16),
    .io_dram_wdata_bits_wdata_17(dramArbs_0_io_dram_wdata_bits_wdata_17),
    .io_dram_wdata_bits_wdata_18(dramArbs_0_io_dram_wdata_bits_wdata_18),
    .io_dram_wdata_bits_wdata_19(dramArbs_0_io_dram_wdata_bits_wdata_19),
    .io_dram_wdata_bits_wdata_20(dramArbs_0_io_dram_wdata_bits_wdata_20),
    .io_dram_wdata_bits_wdata_21(dramArbs_0_io_dram_wdata_bits_wdata_21),
    .io_dram_wdata_bits_wdata_22(dramArbs_0_io_dram_wdata_bits_wdata_22),
    .io_dram_wdata_bits_wdata_23(dramArbs_0_io_dram_wdata_bits_wdata_23),
    .io_dram_wdata_bits_wdata_24(dramArbs_0_io_dram_wdata_bits_wdata_24),
    .io_dram_wdata_bits_wdata_25(dramArbs_0_io_dram_wdata_bits_wdata_25),
    .io_dram_wdata_bits_wdata_26(dramArbs_0_io_dram_wdata_bits_wdata_26),
    .io_dram_wdata_bits_wdata_27(dramArbs_0_io_dram_wdata_bits_wdata_27),
    .io_dram_wdata_bits_wdata_28(dramArbs_0_io_dram_wdata_bits_wdata_28),
    .io_dram_wdata_bits_wdata_29(dramArbs_0_io_dram_wdata_bits_wdata_29),
    .io_dram_wdata_bits_wdata_30(dramArbs_0_io_dram_wdata_bits_wdata_30),
    .io_dram_wdata_bits_wdata_31(dramArbs_0_io_dram_wdata_bits_wdata_31),
    .io_dram_wdata_bits_wdata_32(dramArbs_0_io_dram_wdata_bits_wdata_32),
    .io_dram_wdata_bits_wdata_33(dramArbs_0_io_dram_wdata_bits_wdata_33),
    .io_dram_wdata_bits_wdata_34(dramArbs_0_io_dram_wdata_bits_wdata_34),
    .io_dram_wdata_bits_wdata_35(dramArbs_0_io_dram_wdata_bits_wdata_35),
    .io_dram_wdata_bits_wdata_36(dramArbs_0_io_dram_wdata_bits_wdata_36),
    .io_dram_wdata_bits_wdata_37(dramArbs_0_io_dram_wdata_bits_wdata_37),
    .io_dram_wdata_bits_wdata_38(dramArbs_0_io_dram_wdata_bits_wdata_38),
    .io_dram_wdata_bits_wdata_39(dramArbs_0_io_dram_wdata_bits_wdata_39),
    .io_dram_wdata_bits_wdata_40(dramArbs_0_io_dram_wdata_bits_wdata_40),
    .io_dram_wdata_bits_wdata_41(dramArbs_0_io_dram_wdata_bits_wdata_41),
    .io_dram_wdata_bits_wdata_42(dramArbs_0_io_dram_wdata_bits_wdata_42),
    .io_dram_wdata_bits_wdata_43(dramArbs_0_io_dram_wdata_bits_wdata_43),
    .io_dram_wdata_bits_wdata_44(dramArbs_0_io_dram_wdata_bits_wdata_44),
    .io_dram_wdata_bits_wdata_45(dramArbs_0_io_dram_wdata_bits_wdata_45),
    .io_dram_wdata_bits_wdata_46(dramArbs_0_io_dram_wdata_bits_wdata_46),
    .io_dram_wdata_bits_wdata_47(dramArbs_0_io_dram_wdata_bits_wdata_47),
    .io_dram_wdata_bits_wdata_48(dramArbs_0_io_dram_wdata_bits_wdata_48),
    .io_dram_wdata_bits_wdata_49(dramArbs_0_io_dram_wdata_bits_wdata_49),
    .io_dram_wdata_bits_wdata_50(dramArbs_0_io_dram_wdata_bits_wdata_50),
    .io_dram_wdata_bits_wdata_51(dramArbs_0_io_dram_wdata_bits_wdata_51),
    .io_dram_wdata_bits_wdata_52(dramArbs_0_io_dram_wdata_bits_wdata_52),
    .io_dram_wdata_bits_wdata_53(dramArbs_0_io_dram_wdata_bits_wdata_53),
    .io_dram_wdata_bits_wdata_54(dramArbs_0_io_dram_wdata_bits_wdata_54),
    .io_dram_wdata_bits_wdata_55(dramArbs_0_io_dram_wdata_bits_wdata_55),
    .io_dram_wdata_bits_wdata_56(dramArbs_0_io_dram_wdata_bits_wdata_56),
    .io_dram_wdata_bits_wdata_57(dramArbs_0_io_dram_wdata_bits_wdata_57),
    .io_dram_wdata_bits_wdata_58(dramArbs_0_io_dram_wdata_bits_wdata_58),
    .io_dram_wdata_bits_wdata_59(dramArbs_0_io_dram_wdata_bits_wdata_59),
    .io_dram_wdata_bits_wdata_60(dramArbs_0_io_dram_wdata_bits_wdata_60),
    .io_dram_wdata_bits_wdata_61(dramArbs_0_io_dram_wdata_bits_wdata_61),
    .io_dram_wdata_bits_wdata_62(dramArbs_0_io_dram_wdata_bits_wdata_62),
    .io_dram_wdata_bits_wdata_63(dramArbs_0_io_dram_wdata_bits_wdata_63),
    .io_dram_wdata_bits_wstrb_0(dramArbs_0_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_0_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_0_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_0_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_0_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_0_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_0_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_0_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_0_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_0_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_0_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_0_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_0_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_0_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_0_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_0_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_0_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_0_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_0_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_0_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_0_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_0_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_0_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_0_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_0_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_0_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_0_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_0_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_0_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_0_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_0_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_0_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_0_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_0_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_0_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_0_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_0_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_0_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_0_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_0_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_0_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_0_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_0_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_0_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_0_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_0_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_0_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_0_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_0_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_0_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_0_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_0_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_0_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_0_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_0_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_0_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_0_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_0_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_0_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_0_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_0_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_0_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_0_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_0_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_0_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_0_io_dram_rresp_ready),
    .io_dram_rresp_valid(dramArbs_0_io_dram_rresp_valid),
    .io_dram_rresp_bits_rdata_0(dramArbs_0_io_dram_rresp_bits_rdata_0),
    .io_dram_rresp_bits_rdata_1(dramArbs_0_io_dram_rresp_bits_rdata_1),
    .io_dram_rresp_bits_rdata_2(dramArbs_0_io_dram_rresp_bits_rdata_2),
    .io_dram_rresp_bits_rdata_3(dramArbs_0_io_dram_rresp_bits_rdata_3),
    .io_dram_rresp_bits_rdata_4(dramArbs_0_io_dram_rresp_bits_rdata_4),
    .io_dram_rresp_bits_rdata_5(dramArbs_0_io_dram_rresp_bits_rdata_5),
    .io_dram_rresp_bits_rdata_6(dramArbs_0_io_dram_rresp_bits_rdata_6),
    .io_dram_rresp_bits_rdata_7(dramArbs_0_io_dram_rresp_bits_rdata_7),
    .io_dram_rresp_bits_rdata_8(dramArbs_0_io_dram_rresp_bits_rdata_8),
    .io_dram_rresp_bits_rdata_9(dramArbs_0_io_dram_rresp_bits_rdata_9),
    .io_dram_rresp_bits_rdata_10(dramArbs_0_io_dram_rresp_bits_rdata_10),
    .io_dram_rresp_bits_rdata_11(dramArbs_0_io_dram_rresp_bits_rdata_11),
    .io_dram_rresp_bits_rdata_12(dramArbs_0_io_dram_rresp_bits_rdata_12),
    .io_dram_rresp_bits_rdata_13(dramArbs_0_io_dram_rresp_bits_rdata_13),
    .io_dram_rresp_bits_rdata_14(dramArbs_0_io_dram_rresp_bits_rdata_14),
    .io_dram_rresp_bits_rdata_15(dramArbs_0_io_dram_rresp_bits_rdata_15),
    .io_dram_rresp_bits_rdata_16(dramArbs_0_io_dram_rresp_bits_rdata_16),
    .io_dram_rresp_bits_rdata_17(dramArbs_0_io_dram_rresp_bits_rdata_17),
    .io_dram_rresp_bits_rdata_18(dramArbs_0_io_dram_rresp_bits_rdata_18),
    .io_dram_rresp_bits_rdata_19(dramArbs_0_io_dram_rresp_bits_rdata_19),
    .io_dram_rresp_bits_rdata_20(dramArbs_0_io_dram_rresp_bits_rdata_20),
    .io_dram_rresp_bits_rdata_21(dramArbs_0_io_dram_rresp_bits_rdata_21),
    .io_dram_rresp_bits_rdata_22(dramArbs_0_io_dram_rresp_bits_rdata_22),
    .io_dram_rresp_bits_rdata_23(dramArbs_0_io_dram_rresp_bits_rdata_23),
    .io_dram_rresp_bits_rdata_24(dramArbs_0_io_dram_rresp_bits_rdata_24),
    .io_dram_rresp_bits_rdata_25(dramArbs_0_io_dram_rresp_bits_rdata_25),
    .io_dram_rresp_bits_rdata_26(dramArbs_0_io_dram_rresp_bits_rdata_26),
    .io_dram_rresp_bits_rdata_27(dramArbs_0_io_dram_rresp_bits_rdata_27),
    .io_dram_rresp_bits_rdata_28(dramArbs_0_io_dram_rresp_bits_rdata_28),
    .io_dram_rresp_bits_rdata_29(dramArbs_0_io_dram_rresp_bits_rdata_29),
    .io_dram_rresp_bits_rdata_30(dramArbs_0_io_dram_rresp_bits_rdata_30),
    .io_dram_rresp_bits_rdata_31(dramArbs_0_io_dram_rresp_bits_rdata_31),
    .io_dram_rresp_bits_rdata_32(dramArbs_0_io_dram_rresp_bits_rdata_32),
    .io_dram_rresp_bits_rdata_33(dramArbs_0_io_dram_rresp_bits_rdata_33),
    .io_dram_rresp_bits_rdata_34(dramArbs_0_io_dram_rresp_bits_rdata_34),
    .io_dram_rresp_bits_rdata_35(dramArbs_0_io_dram_rresp_bits_rdata_35),
    .io_dram_rresp_bits_rdata_36(dramArbs_0_io_dram_rresp_bits_rdata_36),
    .io_dram_rresp_bits_rdata_37(dramArbs_0_io_dram_rresp_bits_rdata_37),
    .io_dram_rresp_bits_rdata_38(dramArbs_0_io_dram_rresp_bits_rdata_38),
    .io_dram_rresp_bits_rdata_39(dramArbs_0_io_dram_rresp_bits_rdata_39),
    .io_dram_rresp_bits_rdata_40(dramArbs_0_io_dram_rresp_bits_rdata_40),
    .io_dram_rresp_bits_rdata_41(dramArbs_0_io_dram_rresp_bits_rdata_41),
    .io_dram_rresp_bits_rdata_42(dramArbs_0_io_dram_rresp_bits_rdata_42),
    .io_dram_rresp_bits_rdata_43(dramArbs_0_io_dram_rresp_bits_rdata_43),
    .io_dram_rresp_bits_rdata_44(dramArbs_0_io_dram_rresp_bits_rdata_44),
    .io_dram_rresp_bits_rdata_45(dramArbs_0_io_dram_rresp_bits_rdata_45),
    .io_dram_rresp_bits_rdata_46(dramArbs_0_io_dram_rresp_bits_rdata_46),
    .io_dram_rresp_bits_rdata_47(dramArbs_0_io_dram_rresp_bits_rdata_47),
    .io_dram_rresp_bits_rdata_48(dramArbs_0_io_dram_rresp_bits_rdata_48),
    .io_dram_rresp_bits_rdata_49(dramArbs_0_io_dram_rresp_bits_rdata_49),
    .io_dram_rresp_bits_rdata_50(dramArbs_0_io_dram_rresp_bits_rdata_50),
    .io_dram_rresp_bits_rdata_51(dramArbs_0_io_dram_rresp_bits_rdata_51),
    .io_dram_rresp_bits_rdata_52(dramArbs_0_io_dram_rresp_bits_rdata_52),
    .io_dram_rresp_bits_rdata_53(dramArbs_0_io_dram_rresp_bits_rdata_53),
    .io_dram_rresp_bits_rdata_54(dramArbs_0_io_dram_rresp_bits_rdata_54),
    .io_dram_rresp_bits_rdata_55(dramArbs_0_io_dram_rresp_bits_rdata_55),
    .io_dram_rresp_bits_rdata_56(dramArbs_0_io_dram_rresp_bits_rdata_56),
    .io_dram_rresp_bits_rdata_57(dramArbs_0_io_dram_rresp_bits_rdata_57),
    .io_dram_rresp_bits_rdata_58(dramArbs_0_io_dram_rresp_bits_rdata_58),
    .io_dram_rresp_bits_rdata_59(dramArbs_0_io_dram_rresp_bits_rdata_59),
    .io_dram_rresp_bits_rdata_60(dramArbs_0_io_dram_rresp_bits_rdata_60),
    .io_dram_rresp_bits_rdata_61(dramArbs_0_io_dram_rresp_bits_rdata_61),
    .io_dram_rresp_bits_rdata_62(dramArbs_0_io_dram_rresp_bits_rdata_62),
    .io_dram_rresp_bits_rdata_63(dramArbs_0_io_dram_rresp_bits_rdata_63),
    .io_dram_rresp_bits_tag(dramArbs_0_io_dram_rresp_bits_tag),
    .io_dram_wresp_ready(dramArbs_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_0_io_dram_wresp_bits_tag),
    .io_debugSignals_0(dramArbs_0_io_debugSignals_0),
    .io_debugSignals_1(dramArbs_0_io_debugSignals_1),
    .io_debugSignals_2(dramArbs_0_io_debugSignals_2),
    .io_debugSignals_3(dramArbs_0_io_debugSignals_3),
    .io_debugSignals_4(dramArbs_0_io_debugSignals_4),
    .io_debugSignals_5(dramArbs_0_io_debugSignals_5),
    .io_debugSignals_6(dramArbs_0_io_debugSignals_6),
    .io_debugSignals_7(dramArbs_0_io_debugSignals_7),
    .io_debugSignals_8(dramArbs_0_io_debugSignals_8),
    .io_debugSignals_9(dramArbs_0_io_debugSignals_9),
    .io_debugSignals_10(dramArbs_0_io_debugSignals_10),
    .io_debugSignals_11(dramArbs_0_io_debugSignals_11),
    .io_debugSignals_12(dramArbs_0_io_debugSignals_12),
    .io_debugSignals_13(dramArbs_0_io_debugSignals_13),
    .io_debugSignals_14(dramArbs_0_io_debugSignals_14),
    .io_debugSignals_15(dramArbs_0_io_debugSignals_15),
    .io_debugSignals_16(dramArbs_0_io_debugSignals_16),
    .io_debugSignals_17(dramArbs_0_io_debugSignals_17),
    .io_debugSignals_18(dramArbs_0_io_debugSignals_18),
    .io_debugSignals_19(dramArbs_0_io_debugSignals_19),
    .io_debugSignals_20(dramArbs_0_io_debugSignals_20),
    .io_debugSignals_21(dramArbs_0_io_debugSignals_21),
    .io_debugSignals_22(dramArbs_0_io_debugSignals_22),
    .io_debugSignals_23(dramArbs_0_io_debugSignals_23),
    .io_debugSignals_24(dramArbs_0_io_debugSignals_24),
    .io_debugSignals_25(dramArbs_0_io_debugSignals_25),
    .io_debugSignals_26(dramArbs_0_io_debugSignals_26),
    .io_debugSignals_27(dramArbs_0_io_debugSignals_27),
    .io_debugSignals_28(dramArbs_0_io_debugSignals_28),
    .io_debugSignals_29(dramArbs_0_io_debugSignals_29),
    .io_debugSignals_30(dramArbs_0_io_debugSignals_30),
    .io_debugSignals_41(dramArbs_0_io_debugSignals_41)
  );
  DRAMHeap heap ( // @[Fringe.scala 107:20:@153928.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@153937.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argIns_3(regs_io_argIns_3),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits),
    .io_argOuts_2_valid(regs_io_argOuts_2_valid),
    .io_argOuts_2_bits(regs_io_argOuts_2_bits),
    .io_argOuts_3_valid(regs_io_argOuts_3_valid),
    .io_argOuts_3_bits(regs_io_argOuts_3_bits),
    .io_argOuts_4_valid(regs_io_argOuts_4_valid),
    .io_argOuts_4_bits(regs_io_argOuts_4_bits),
    .io_argOuts_5_valid(regs_io_argOuts_5_valid),
    .io_argOuts_5_bits(regs_io_argOuts_5_bits),
    .io_argOuts_6_valid(regs_io_argOuts_6_valid),
    .io_argOuts_6_bits(regs_io_argOuts_6_bits),
    .io_argOuts_7_valid(regs_io_argOuts_7_valid),
    .io_argOuts_7_bits(regs_io_argOuts_7_bits),
    .io_argOuts_8_valid(regs_io_argOuts_8_valid),
    .io_argOuts_8_bits(regs_io_argOuts_8_bits),
    .io_argOuts_9_valid(regs_io_argOuts_9_valid),
    .io_argOuts_9_bits(regs_io_argOuts_9_bits),
    .io_argOuts_10_valid(regs_io_argOuts_10_valid),
    .io_argOuts_10_bits(regs_io_argOuts_10_bits),
    .io_argOuts_11_valid(regs_io_argOuts_11_valid),
    .io_argOuts_11_bits(regs_io_argOuts_11_bits),
    .io_argOuts_12_valid(regs_io_argOuts_12_valid),
    .io_argOuts_12_bits(regs_io_argOuts_12_bits),
    .io_argOuts_13_valid(regs_io_argOuts_13_valid),
    .io_argOuts_13_bits(regs_io_argOuts_13_bits),
    .io_argOuts_14_valid(regs_io_argOuts_14_valid),
    .io_argOuts_14_bits(regs_io_argOuts_14_bits),
    .io_argOuts_15_valid(regs_io_argOuts_15_valid),
    .io_argOuts_15_bits(regs_io_argOuts_15_bits),
    .io_argOuts_16_valid(regs_io_argOuts_16_valid),
    .io_argOuts_16_bits(regs_io_argOuts_16_bits),
    .io_argOuts_17_valid(regs_io_argOuts_17_valid),
    .io_argOuts_17_bits(regs_io_argOuts_17_bits),
    .io_argOuts_18_valid(regs_io_argOuts_18_valid),
    .io_argOuts_18_bits(regs_io_argOuts_18_bits),
    .io_argOuts_19_valid(regs_io_argOuts_19_valid),
    .io_argOuts_19_bits(regs_io_argOuts_19_bits),
    .io_argOuts_20_valid(regs_io_argOuts_20_valid),
    .io_argOuts_20_bits(regs_io_argOuts_20_bits),
    .io_argOuts_21_valid(regs_io_argOuts_21_valid),
    .io_argOuts_21_bits(regs_io_argOuts_21_bits),
    .io_argOuts_22_valid(regs_io_argOuts_22_valid),
    .io_argOuts_22_bits(regs_io_argOuts_22_bits),
    .io_argOuts_23_valid(regs_io_argOuts_23_valid),
    .io_argOuts_23_bits(regs_io_argOuts_23_bits),
    .io_argOuts_24_valid(regs_io_argOuts_24_valid),
    .io_argOuts_24_bits(regs_io_argOuts_24_bits),
    .io_argOuts_25_valid(regs_io_argOuts_25_valid),
    .io_argOuts_25_bits(regs_io_argOuts_25_bits),
    .io_argOuts_26_valid(regs_io_argOuts_26_valid),
    .io_argOuts_26_bits(regs_io_argOuts_26_bits),
    .io_argOuts_27_valid(regs_io_argOuts_27_valid),
    .io_argOuts_27_bits(regs_io_argOuts_27_bits),
    .io_argOuts_28_valid(regs_io_argOuts_28_valid),
    .io_argOuts_28_bits(regs_io_argOuts_28_bits),
    .io_argOuts_29_valid(regs_io_argOuts_29_valid),
    .io_argOuts_29_bits(regs_io_argOuts_29_bits),
    .io_argOuts_30_valid(regs_io_argOuts_30_valid),
    .io_argOuts_30_bits(regs_io_argOuts_30_bits),
    .io_argOuts_31_valid(regs_io_argOuts_31_valid),
    .io_argOuts_31_bits(regs_io_argOuts_31_bits),
    .io_argOuts_32_valid(regs_io_argOuts_32_valid),
    .io_argOuts_32_bits(regs_io_argOuts_32_bits),
    .io_argOuts_33_valid(regs_io_argOuts_33_valid),
    .io_argOuts_33_bits(regs_io_argOuts_33_bits),
    .io_argOuts_34_valid(regs_io_argOuts_34_valid),
    .io_argOuts_34_bits(regs_io_argOuts_34_bits),
    .io_argOuts_35_valid(regs_io_argOuts_35_valid),
    .io_argOuts_35_bits(regs_io_argOuts_35_bits),
    .io_argOuts_36_valid(regs_io_argOuts_36_valid),
    .io_argOuts_36_bits(regs_io_argOuts_36_bits),
    .io_argOuts_37_valid(regs_io_argOuts_37_valid),
    .io_argOuts_37_bits(regs_io_argOuts_37_bits),
    .io_argOuts_38_valid(regs_io_argOuts_38_valid),
    .io_argOuts_38_bits(regs_io_argOuts_38_bits),
    .io_argOuts_39_valid(regs_io_argOuts_39_valid),
    .io_argOuts_39_bits(regs_io_argOuts_39_bits),
    .io_argOuts_40_valid(regs_io_argOuts_40_valid),
    .io_argOuts_40_bits(regs_io_argOuts_40_bits),
    .io_argOuts_41_valid(regs_io_argOuts_41_valid),
    .io_argOuts_41_bits(regs_io_argOuts_41_bits),
    .io_argOuts_42_valid(regs_io_argOuts_42_valid),
    .io_argOuts_42_bits(regs_io_argOuts_42_bits),
    .io_argOuts_43_valid(regs_io_argOuts_43_valid),
    .io_argOuts_43_bits(regs_io_argOuts_43_bits),
    .io_argOuts_44_valid(regs_io_argOuts_44_valid),
    .io_argOuts_44_bits(regs_io_argOuts_44_bits),
    .io_argOuts_45_valid(regs_io_argOuts_45_valid),
    .io_argOuts_45_bits(regs_io_argOuts_45_bits),
    .io_argOuts_46_valid(regs_io_argOuts_46_valid),
    .io_argOuts_46_bits(regs_io_argOuts_46_bits),
    .io_argOuts_47_valid(regs_io_argOuts_47_valid),
    .io_argOuts_47_bits(regs_io_argOuts_47_bits),
    .io_argOuts_48_valid(regs_io_argOuts_48_valid),
    .io_argOuts_48_bits(regs_io_argOuts_48_bits),
    .io_argOuts_49_valid(regs_io_argOuts_49_valid),
    .io_argOuts_49_bits(regs_io_argOuts_49_bits),
    .io_argOuts_50_valid(regs_io_argOuts_50_valid),
    .io_argOuts_50_bits(regs_io_argOuts_50_bits),
    .io_argOuts_51_valid(regs_io_argOuts_51_valid),
    .io_argOuts_51_bits(regs_io_argOuts_51_bits),
    .io_argOuts_52_valid(regs_io_argOuts_52_valid),
    .io_argOuts_52_bits(regs_io_argOuts_52_bits),
    .io_argOuts_53_valid(regs_io_argOuts_53_valid),
    .io_argOuts_53_bits(regs_io_argOuts_53_bits),
    .io_argOuts_54_valid(regs_io_argOuts_54_valid),
    .io_argOuts_54_bits(regs_io_argOuts_54_bits),
    .io_argOuts_55_valid(regs_io_argOuts_55_valid),
    .io_argOuts_55_bits(regs_io_argOuts_55_bits),
    .io_argOuts_56_valid(regs_io_argOuts_56_valid),
    .io_argOuts_56_bits(regs_io_argOuts_56_bits),
    .io_argOuts_57_valid(regs_io_argOuts_57_valid),
    .io_argOuts_57_bits(regs_io_argOuts_57_bits),
    .io_argOuts_58_valid(regs_io_argOuts_58_valid),
    .io_argOuts_58_bits(regs_io_argOuts_58_bits),
    .io_argOuts_59_valid(regs_io_argOuts_59_valid),
    .io_argOuts_59_bits(regs_io_argOuts_59_bits),
    .io_argOuts_60_valid(regs_io_argOuts_60_valid),
    .io_argOuts_60_bits(regs_io_argOuts_60_bits),
    .io_argOuts_61_bits(regs_io_argOuts_61_bits),
    .io_argOuts_62_bits(regs_io_argOuts_62_bits),
    .io_argOuts_63_bits(regs_io_argOuts_63_bits),
    .io_argOuts_64_bits(regs_io_argOuts_64_bits),
    .io_argOuts_65_bits(regs_io_argOuts_65_bits),
    .io_argOuts_66_bits(regs_io_argOuts_66_bits),
    .io_argOuts_67_bits(regs_io_argOuts_67_bits),
    .io_argOuts_68_bits(regs_io_argOuts_68_bits),
    .io_argOuts_69_bits(regs_io_argOuts_69_bits),
    .io_argOuts_70_bits(regs_io_argOuts_70_bits),
    .io_argOuts_71_bits(regs_io_argOuts_71_bits),
    .io_argOuts_72_bits(regs_io_argOuts_72_bits),
    .io_argOuts_73_bits(regs_io_argOuts_73_bits),
    .io_argOuts_74_bits(regs_io_argOuts_74_bits),
    .io_argOuts_75_bits(regs_io_argOuts_75_bits),
    .io_argOuts_76_bits(regs_io_argOuts_76_bits),
    .io_argOuts_77_bits(regs_io_argOuts_77_bits),
    .io_argOuts_78_bits(regs_io_argOuts_78_bits),
    .io_argOuts_79_bits(regs_io_argOuts_79_bits),
    .io_argOuts_80_bits(regs_io_argOuts_80_bits),
    .io_argOuts_81_bits(regs_io_argOuts_81_bits),
    .io_argOuts_82_bits(regs_io_argOuts_82_bits),
    .io_argOuts_83_bits(regs_io_argOuts_83_bits),
    .io_argOuts_84_bits(regs_io_argOuts_84_bits),
    .io_argOuts_85_bits(regs_io_argOuts_85_bits),
    .io_argOuts_86_bits(regs_io_argOuts_86_bits),
    .io_argOuts_87_bits(regs_io_argOuts_87_bits),
    .io_argOuts_88_bits(regs_io_argOuts_88_bits),
    .io_argOuts_89_bits(regs_io_argOuts_89_bits),
    .io_argOuts_90_bits(regs_io_argOuts_90_bits),
    .io_argOuts_91_bits(regs_io_argOuts_91_bits),
    .io_argOuts_102_bits(regs_io_argOuts_102_bits),
    .io_argEchos_1(regs_io_argEchos_1),
    .io_argEchos_2(regs_io_argEchos_2),
    .io_argEchos_3(regs_io_argEchos_3),
    .io_argEchos_4(regs_io_argEchos_4),
    .io_argEchos_5(regs_io_argEchos_5),
    .io_argEchos_6(regs_io_argEchos_6),
    .io_argEchos_7(regs_io_argEchos_7),
    .io_argEchos_8(regs_io_argEchos_8),
    .io_argEchos_9(regs_io_argEchos_9),
    .io_argEchos_10(regs_io_argEchos_10),
    .io_argEchos_11(regs_io_argEchos_11),
    .io_argEchos_12(regs_io_argEchos_12),
    .io_argEchos_13(regs_io_argEchos_13),
    .io_argEchos_14(regs_io_argEchos_14),
    .io_argEchos_15(regs_io_argEchos_15),
    .io_argEchos_16(regs_io_argEchos_16),
    .io_argEchos_17(regs_io_argEchos_17),
    .io_argEchos_18(regs_io_argEchos_18),
    .io_argEchos_19(regs_io_argEchos_19),
    .io_argEchos_20(regs_io_argEchos_20),
    .io_argEchos_21(regs_io_argEchos_21),
    .io_argEchos_22(regs_io_argEchos_22),
    .io_argEchos_23(regs_io_argEchos_23),
    .io_argEchos_24(regs_io_argEchos_24),
    .io_argEchos_25(regs_io_argEchos_25),
    .io_argEchos_26(regs_io_argEchos_26),
    .io_argEchos_27(regs_io_argEchos_27),
    .io_argEchos_28(regs_io_argEchos_28),
    .io_argEchos_29(regs_io_argEchos_29),
    .io_argEchos_30(regs_io_argEchos_30),
    .io_argEchos_31(regs_io_argEchos_31),
    .io_argEchos_32(regs_io_argEchos_32),
    .io_argEchos_33(regs_io_argEchos_33),
    .io_argEchos_34(regs_io_argEchos_34),
    .io_argEchos_35(regs_io_argEchos_35),
    .io_argEchos_36(regs_io_argEchos_36),
    .io_argEchos_37(regs_io_argEchos_37),
    .io_argEchos_38(regs_io_argEchos_38),
    .io_argEchos_39(regs_io_argEchos_39),
    .io_argEchos_40(regs_io_argEchos_40),
    .io_argEchos_41(regs_io_argEchos_41),
    .io_argEchos_42(regs_io_argEchos_42),
    .io_argEchos_43(regs_io_argEchos_43),
    .io_argEchos_44(regs_io_argEchos_44),
    .io_argEchos_45(regs_io_argEchos_45),
    .io_argEchos_46(regs_io_argEchos_46),
    .io_argEchos_47(regs_io_argEchos_47),
    .io_argEchos_48(regs_io_argEchos_48),
    .io_argEchos_49(regs_io_argEchos_49),
    .io_argEchos_50(regs_io_argEchos_50),
    .io_argEchos_51(regs_io_argEchos_51),
    .io_argEchos_52(regs_io_argEchos_52),
    .io_argEchos_53(regs_io_argEchos_53),
    .io_argEchos_54(regs_io_argEchos_54),
    .io_argEchos_55(regs_io_argEchos_55),
    .io_argEchos_56(regs_io_argEchos_56),
    .io_argEchos_57(regs_io_argEchos_57),
    .io_argEchos_58(regs_io_argEchos_58),
    .io_argEchos_59(regs_io_argEchos_59),
    .io_argEchos_60(regs_io_argEchos_60)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@156227.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@156246.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_953 = regs_io_argIns_1; // @[:@156204.4 :@156205.4]
  assign curStatus_done = _T_953[0]; // @[Fringe.scala 133:45:@156206.4]
  assign curStatus_timeout = _T_953[1]; // @[Fringe.scala 133:45:@156208.4]
  assign curStatus_allocDealloc = _T_953[4:2]; // @[Fringe.scala 133:45:@156210.4]
  assign curStatus_sizeAddr = _T_953[63:5]; // @[Fringe.scala 133:45:@156212.4]
  assign _T_958 = regs_io_argIns_0[0]; // @[Fringe.scala 134:60:@156214.4]
  assign _T_962 = curStatus_done == 1'h0; // @[Fringe.scala 134:74:@156216.4]
  assign _T_963 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@156218.4]
  assign _T_973 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@156254.4]
  assign _T_981 = _T_980 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@156259.4]
  assign _T_982 = heap_io_host_0_req_valid & _T_981; // @[package.scala 153:8:@156260.4]
  assign _T_985 = _T_958 & depulser_io_out; // @[Fringe.scala 160:55:@156264.4]
  assign status_bits_done = depulser_io_out ? _T_985 : curStatus_done; // @[Fringe.scala 160:26:@156265.4]
  assign _T_988 = _T_958 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@156268.4]
  assign status_bits_timeout = depulser_io_out ? _T_988 : curStatus_timeout; // @[Fringe.scala 161:29:@156269.4]
  assign _T_992 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@156271.4]
  assign _T_994 = heap_io_host_0_req_valid ? _T_992 : 2'h0; // @[Fringe.scala 162:34:@156272.4]
  assign _T_996 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@156274.4]
  assign _T_997 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@156277.4]
  assign status_bits_sizeAddr = _T_996[58:0]; // @[Fringe.scala 158:20:@156256.4 Fringe.scala 163:24:@156275.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_994}; // @[Fringe.scala 158:20:@156256.4 Fringe.scala 162:28:@156273.4]
  assign _T_998 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@156278.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@157672.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@157673.4]
  assign _T_1502 = alloc | dealloc; // @[Fringe.scala 204:37:@157674.4]
  assign _T_1506 = _T_1505 ^ _T_1502; // @[package.scala 153:13:@157677.4]
  assign io_rdata = _T_949; // @[Fringe.scala 128:14:@156202.4]
  assign io_enable = _T_958 & _T_962; // @[Fringe.scala 136:13:@156222.4]
  assign io_reset = _T_963 | reset; // @[Fringe.scala 137:12:@156223.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@156244.4]
  assign io_argIns_1 = regs_io_argIns_3; // @[Fringe.scala 151:51:@156245.4]
  assign io_argEchos_0 = regs_io_argEchos_1; // @[Fringe.scala 174:24:@156281.4]
  assign io_argEchos_1 = regs_io_argEchos_2; // @[Fringe.scala 174:24:@156284.4]
  assign io_argEchos_2 = regs_io_argEchos_3; // @[Fringe.scala 174:24:@156287.4]
  assign io_argEchos_3 = regs_io_argEchos_4; // @[Fringe.scala 174:24:@156290.4]
  assign io_argEchos_4 = regs_io_argEchos_5; // @[Fringe.scala 174:24:@156293.4]
  assign io_argEchos_5 = regs_io_argEchos_6; // @[Fringe.scala 174:24:@156296.4]
  assign io_argEchos_6 = regs_io_argEchos_7; // @[Fringe.scala 174:24:@156299.4]
  assign io_argEchos_7 = regs_io_argEchos_8; // @[Fringe.scala 174:24:@156302.4]
  assign io_argEchos_8 = regs_io_argEchos_9; // @[Fringe.scala 174:24:@156305.4]
  assign io_argEchos_9 = regs_io_argEchos_10; // @[Fringe.scala 174:24:@156308.4]
  assign io_argEchos_10 = regs_io_argEchos_11; // @[Fringe.scala 174:24:@156311.4]
  assign io_argEchos_11 = regs_io_argEchos_12; // @[Fringe.scala 174:24:@156314.4]
  assign io_argEchos_12 = regs_io_argEchos_13; // @[Fringe.scala 174:24:@156317.4]
  assign io_argEchos_13 = regs_io_argEchos_14; // @[Fringe.scala 174:24:@156320.4]
  assign io_argEchos_14 = regs_io_argEchos_15; // @[Fringe.scala 174:24:@156323.4]
  assign io_argEchos_15 = regs_io_argEchos_16; // @[Fringe.scala 174:24:@156326.4]
  assign io_argEchos_16 = regs_io_argEchos_17; // @[Fringe.scala 174:24:@156329.4]
  assign io_argEchos_17 = regs_io_argEchos_18; // @[Fringe.scala 174:24:@156332.4]
  assign io_argEchos_18 = regs_io_argEchos_19; // @[Fringe.scala 174:24:@156335.4]
  assign io_argEchos_19 = regs_io_argEchos_20; // @[Fringe.scala 174:24:@156338.4]
  assign io_argEchos_20 = regs_io_argEchos_21; // @[Fringe.scala 174:24:@156341.4]
  assign io_argEchos_21 = regs_io_argEchos_22; // @[Fringe.scala 174:24:@156344.4]
  assign io_argEchos_22 = regs_io_argEchos_23; // @[Fringe.scala 174:24:@156347.4]
  assign io_argEchos_23 = regs_io_argEchos_24; // @[Fringe.scala 174:24:@156350.4]
  assign io_argEchos_24 = regs_io_argEchos_25; // @[Fringe.scala 174:24:@156353.4]
  assign io_argEchos_25 = regs_io_argEchos_26; // @[Fringe.scala 174:24:@156356.4]
  assign io_argEchos_26 = regs_io_argEchos_27; // @[Fringe.scala 174:24:@156359.4]
  assign io_argEchos_27 = regs_io_argEchos_28; // @[Fringe.scala 174:24:@156362.4]
  assign io_argEchos_28 = regs_io_argEchos_29; // @[Fringe.scala 174:24:@156365.4]
  assign io_argEchos_29 = regs_io_argEchos_30; // @[Fringe.scala 174:24:@156368.4]
  assign io_argEchos_30 = regs_io_argEchos_31; // @[Fringe.scala 174:24:@156371.4]
  assign io_argEchos_31 = regs_io_argEchos_32; // @[Fringe.scala 174:24:@156374.4]
  assign io_argEchos_32 = regs_io_argEchos_33; // @[Fringe.scala 174:24:@156377.4]
  assign io_argEchos_33 = regs_io_argEchos_34; // @[Fringe.scala 174:24:@156380.4]
  assign io_argEchos_34 = regs_io_argEchos_35; // @[Fringe.scala 174:24:@156383.4]
  assign io_argEchos_35 = regs_io_argEchos_36; // @[Fringe.scala 174:24:@156386.4]
  assign io_argEchos_36 = regs_io_argEchos_37; // @[Fringe.scala 174:24:@156389.4]
  assign io_argEchos_37 = regs_io_argEchos_38; // @[Fringe.scala 174:24:@156392.4]
  assign io_argEchos_38 = regs_io_argEchos_39; // @[Fringe.scala 174:24:@156395.4]
  assign io_argEchos_39 = regs_io_argEchos_40; // @[Fringe.scala 174:24:@156398.4]
  assign io_argEchos_40 = regs_io_argEchos_41; // @[Fringe.scala 174:24:@156401.4]
  assign io_argEchos_41 = regs_io_argEchos_42; // @[Fringe.scala 174:24:@156404.4]
  assign io_argEchos_42 = regs_io_argEchos_43; // @[Fringe.scala 174:24:@156407.4]
  assign io_argEchos_43 = regs_io_argEchos_44; // @[Fringe.scala 174:24:@156410.4]
  assign io_argEchos_44 = regs_io_argEchos_45; // @[Fringe.scala 174:24:@156413.4]
  assign io_argEchos_45 = regs_io_argEchos_46; // @[Fringe.scala 174:24:@156416.4]
  assign io_argEchos_46 = regs_io_argEchos_47; // @[Fringe.scala 174:24:@156419.4]
  assign io_argEchos_47 = regs_io_argEchos_48; // @[Fringe.scala 174:24:@156422.4]
  assign io_argEchos_48 = regs_io_argEchos_49; // @[Fringe.scala 174:24:@156425.4]
  assign io_argEchos_49 = regs_io_argEchos_50; // @[Fringe.scala 174:24:@156428.4]
  assign io_argEchos_50 = regs_io_argEchos_51; // @[Fringe.scala 174:24:@156431.4]
  assign io_argEchos_51 = regs_io_argEchos_52; // @[Fringe.scala 174:24:@156434.4]
  assign io_argEchos_52 = regs_io_argEchos_53; // @[Fringe.scala 174:24:@156437.4]
  assign io_argEchos_53 = regs_io_argEchos_54; // @[Fringe.scala 174:24:@156440.4]
  assign io_argEchos_54 = regs_io_argEchos_55; // @[Fringe.scala 174:24:@156443.4]
  assign io_argEchos_55 = regs_io_argEchos_56; // @[Fringe.scala 174:24:@156446.4]
  assign io_argEchos_56 = regs_io_argEchos_57; // @[Fringe.scala 174:24:@156449.4]
  assign io_argEchos_57 = regs_io_argEchos_58; // @[Fringe.scala 174:24:@156452.4]
  assign io_argEchos_58 = regs_io_argEchos_59; // @[Fringe.scala 174:24:@156455.4]
  assign io_argEchos_59 = regs_io_argEchos_60; // @[Fringe.scala 174:24:@156458.4]
  assign io_memStreams_loads_0_cmd_ready = dramArbs_0_io_app_loads_0_cmd_ready; // @[Fringe.scala 100:70:@153651.4]
  assign io_memStreams_loads_0_data_valid = dramArbs_0_io_app_loads_0_data_valid; // @[Fringe.scala 100:70:@153646.4]
  assign io_memStreams_loads_0_data_bits_rdata_0 = dramArbs_0_io_app_loads_0_data_bits_rdata_0; // @[Fringe.scala 100:70:@153645.4]
  assign io_memStreams_stores_0_cmd_ready = dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 101:72:@153662.4]
  assign io_memStreams_stores_0_data_ready = dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 101:72:@153658.4]
  assign io_memStreams_stores_0_wresp_valid = dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 101:72:@153653.4]
  assign io_memStreams_stores_0_wresp_bits = dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 101:72:@153652.4]
  assign io_dram_0_cmd_valid = dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 195:72:@157670.4]
  assign io_dram_0_cmd_bits_addr = dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@157669.4]
  assign io_dram_0_cmd_bits_size = dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@157668.4]
  assign io_dram_0_cmd_bits_rawAddr = dramArbs_0_io_dram_cmd_bits_rawAddr; // @[Fringe.scala 195:72:@157667.4]
  assign io_dram_0_cmd_bits_isWr = dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@157666.4]
  assign io_dram_0_cmd_bits_tag = dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@157665.4]
  assign io_dram_0_wdata_valid = dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 195:72:@157663.4]
  assign io_dram_0_wdata_bits_wdata_0 = dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@157599.4]
  assign io_dram_0_wdata_bits_wdata_1 = dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@157600.4]
  assign io_dram_0_wdata_bits_wdata_2 = dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@157601.4]
  assign io_dram_0_wdata_bits_wdata_3 = dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@157602.4]
  assign io_dram_0_wdata_bits_wdata_4 = dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@157603.4]
  assign io_dram_0_wdata_bits_wdata_5 = dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@157604.4]
  assign io_dram_0_wdata_bits_wdata_6 = dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@157605.4]
  assign io_dram_0_wdata_bits_wdata_7 = dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@157606.4]
  assign io_dram_0_wdata_bits_wdata_8 = dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@157607.4]
  assign io_dram_0_wdata_bits_wdata_9 = dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@157608.4]
  assign io_dram_0_wdata_bits_wdata_10 = dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@157609.4]
  assign io_dram_0_wdata_bits_wdata_11 = dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@157610.4]
  assign io_dram_0_wdata_bits_wdata_12 = dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@157611.4]
  assign io_dram_0_wdata_bits_wdata_13 = dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@157612.4]
  assign io_dram_0_wdata_bits_wdata_14 = dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@157613.4]
  assign io_dram_0_wdata_bits_wdata_15 = dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@157614.4]
  assign io_dram_0_wdata_bits_wdata_16 = dramArbs_0_io_dram_wdata_bits_wdata_16; // @[Fringe.scala 195:72:@157615.4]
  assign io_dram_0_wdata_bits_wdata_17 = dramArbs_0_io_dram_wdata_bits_wdata_17; // @[Fringe.scala 195:72:@157616.4]
  assign io_dram_0_wdata_bits_wdata_18 = dramArbs_0_io_dram_wdata_bits_wdata_18; // @[Fringe.scala 195:72:@157617.4]
  assign io_dram_0_wdata_bits_wdata_19 = dramArbs_0_io_dram_wdata_bits_wdata_19; // @[Fringe.scala 195:72:@157618.4]
  assign io_dram_0_wdata_bits_wdata_20 = dramArbs_0_io_dram_wdata_bits_wdata_20; // @[Fringe.scala 195:72:@157619.4]
  assign io_dram_0_wdata_bits_wdata_21 = dramArbs_0_io_dram_wdata_bits_wdata_21; // @[Fringe.scala 195:72:@157620.4]
  assign io_dram_0_wdata_bits_wdata_22 = dramArbs_0_io_dram_wdata_bits_wdata_22; // @[Fringe.scala 195:72:@157621.4]
  assign io_dram_0_wdata_bits_wdata_23 = dramArbs_0_io_dram_wdata_bits_wdata_23; // @[Fringe.scala 195:72:@157622.4]
  assign io_dram_0_wdata_bits_wdata_24 = dramArbs_0_io_dram_wdata_bits_wdata_24; // @[Fringe.scala 195:72:@157623.4]
  assign io_dram_0_wdata_bits_wdata_25 = dramArbs_0_io_dram_wdata_bits_wdata_25; // @[Fringe.scala 195:72:@157624.4]
  assign io_dram_0_wdata_bits_wdata_26 = dramArbs_0_io_dram_wdata_bits_wdata_26; // @[Fringe.scala 195:72:@157625.4]
  assign io_dram_0_wdata_bits_wdata_27 = dramArbs_0_io_dram_wdata_bits_wdata_27; // @[Fringe.scala 195:72:@157626.4]
  assign io_dram_0_wdata_bits_wdata_28 = dramArbs_0_io_dram_wdata_bits_wdata_28; // @[Fringe.scala 195:72:@157627.4]
  assign io_dram_0_wdata_bits_wdata_29 = dramArbs_0_io_dram_wdata_bits_wdata_29; // @[Fringe.scala 195:72:@157628.4]
  assign io_dram_0_wdata_bits_wdata_30 = dramArbs_0_io_dram_wdata_bits_wdata_30; // @[Fringe.scala 195:72:@157629.4]
  assign io_dram_0_wdata_bits_wdata_31 = dramArbs_0_io_dram_wdata_bits_wdata_31; // @[Fringe.scala 195:72:@157630.4]
  assign io_dram_0_wdata_bits_wdata_32 = dramArbs_0_io_dram_wdata_bits_wdata_32; // @[Fringe.scala 195:72:@157631.4]
  assign io_dram_0_wdata_bits_wdata_33 = dramArbs_0_io_dram_wdata_bits_wdata_33; // @[Fringe.scala 195:72:@157632.4]
  assign io_dram_0_wdata_bits_wdata_34 = dramArbs_0_io_dram_wdata_bits_wdata_34; // @[Fringe.scala 195:72:@157633.4]
  assign io_dram_0_wdata_bits_wdata_35 = dramArbs_0_io_dram_wdata_bits_wdata_35; // @[Fringe.scala 195:72:@157634.4]
  assign io_dram_0_wdata_bits_wdata_36 = dramArbs_0_io_dram_wdata_bits_wdata_36; // @[Fringe.scala 195:72:@157635.4]
  assign io_dram_0_wdata_bits_wdata_37 = dramArbs_0_io_dram_wdata_bits_wdata_37; // @[Fringe.scala 195:72:@157636.4]
  assign io_dram_0_wdata_bits_wdata_38 = dramArbs_0_io_dram_wdata_bits_wdata_38; // @[Fringe.scala 195:72:@157637.4]
  assign io_dram_0_wdata_bits_wdata_39 = dramArbs_0_io_dram_wdata_bits_wdata_39; // @[Fringe.scala 195:72:@157638.4]
  assign io_dram_0_wdata_bits_wdata_40 = dramArbs_0_io_dram_wdata_bits_wdata_40; // @[Fringe.scala 195:72:@157639.4]
  assign io_dram_0_wdata_bits_wdata_41 = dramArbs_0_io_dram_wdata_bits_wdata_41; // @[Fringe.scala 195:72:@157640.4]
  assign io_dram_0_wdata_bits_wdata_42 = dramArbs_0_io_dram_wdata_bits_wdata_42; // @[Fringe.scala 195:72:@157641.4]
  assign io_dram_0_wdata_bits_wdata_43 = dramArbs_0_io_dram_wdata_bits_wdata_43; // @[Fringe.scala 195:72:@157642.4]
  assign io_dram_0_wdata_bits_wdata_44 = dramArbs_0_io_dram_wdata_bits_wdata_44; // @[Fringe.scala 195:72:@157643.4]
  assign io_dram_0_wdata_bits_wdata_45 = dramArbs_0_io_dram_wdata_bits_wdata_45; // @[Fringe.scala 195:72:@157644.4]
  assign io_dram_0_wdata_bits_wdata_46 = dramArbs_0_io_dram_wdata_bits_wdata_46; // @[Fringe.scala 195:72:@157645.4]
  assign io_dram_0_wdata_bits_wdata_47 = dramArbs_0_io_dram_wdata_bits_wdata_47; // @[Fringe.scala 195:72:@157646.4]
  assign io_dram_0_wdata_bits_wdata_48 = dramArbs_0_io_dram_wdata_bits_wdata_48; // @[Fringe.scala 195:72:@157647.4]
  assign io_dram_0_wdata_bits_wdata_49 = dramArbs_0_io_dram_wdata_bits_wdata_49; // @[Fringe.scala 195:72:@157648.4]
  assign io_dram_0_wdata_bits_wdata_50 = dramArbs_0_io_dram_wdata_bits_wdata_50; // @[Fringe.scala 195:72:@157649.4]
  assign io_dram_0_wdata_bits_wdata_51 = dramArbs_0_io_dram_wdata_bits_wdata_51; // @[Fringe.scala 195:72:@157650.4]
  assign io_dram_0_wdata_bits_wdata_52 = dramArbs_0_io_dram_wdata_bits_wdata_52; // @[Fringe.scala 195:72:@157651.4]
  assign io_dram_0_wdata_bits_wdata_53 = dramArbs_0_io_dram_wdata_bits_wdata_53; // @[Fringe.scala 195:72:@157652.4]
  assign io_dram_0_wdata_bits_wdata_54 = dramArbs_0_io_dram_wdata_bits_wdata_54; // @[Fringe.scala 195:72:@157653.4]
  assign io_dram_0_wdata_bits_wdata_55 = dramArbs_0_io_dram_wdata_bits_wdata_55; // @[Fringe.scala 195:72:@157654.4]
  assign io_dram_0_wdata_bits_wdata_56 = dramArbs_0_io_dram_wdata_bits_wdata_56; // @[Fringe.scala 195:72:@157655.4]
  assign io_dram_0_wdata_bits_wdata_57 = dramArbs_0_io_dram_wdata_bits_wdata_57; // @[Fringe.scala 195:72:@157656.4]
  assign io_dram_0_wdata_bits_wdata_58 = dramArbs_0_io_dram_wdata_bits_wdata_58; // @[Fringe.scala 195:72:@157657.4]
  assign io_dram_0_wdata_bits_wdata_59 = dramArbs_0_io_dram_wdata_bits_wdata_59; // @[Fringe.scala 195:72:@157658.4]
  assign io_dram_0_wdata_bits_wdata_60 = dramArbs_0_io_dram_wdata_bits_wdata_60; // @[Fringe.scala 195:72:@157659.4]
  assign io_dram_0_wdata_bits_wdata_61 = dramArbs_0_io_dram_wdata_bits_wdata_61; // @[Fringe.scala 195:72:@157660.4]
  assign io_dram_0_wdata_bits_wdata_62 = dramArbs_0_io_dram_wdata_bits_wdata_62; // @[Fringe.scala 195:72:@157661.4]
  assign io_dram_0_wdata_bits_wdata_63 = dramArbs_0_io_dram_wdata_bits_wdata_63; // @[Fringe.scala 195:72:@157662.4]
  assign io_dram_0_wdata_bits_wstrb_0 = dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@157535.4]
  assign io_dram_0_wdata_bits_wstrb_1 = dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@157536.4]
  assign io_dram_0_wdata_bits_wstrb_2 = dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@157537.4]
  assign io_dram_0_wdata_bits_wstrb_3 = dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@157538.4]
  assign io_dram_0_wdata_bits_wstrb_4 = dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@157539.4]
  assign io_dram_0_wdata_bits_wstrb_5 = dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@157540.4]
  assign io_dram_0_wdata_bits_wstrb_6 = dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@157541.4]
  assign io_dram_0_wdata_bits_wstrb_7 = dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@157542.4]
  assign io_dram_0_wdata_bits_wstrb_8 = dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@157543.4]
  assign io_dram_0_wdata_bits_wstrb_9 = dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@157544.4]
  assign io_dram_0_wdata_bits_wstrb_10 = dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@157545.4]
  assign io_dram_0_wdata_bits_wstrb_11 = dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@157546.4]
  assign io_dram_0_wdata_bits_wstrb_12 = dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@157547.4]
  assign io_dram_0_wdata_bits_wstrb_13 = dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@157548.4]
  assign io_dram_0_wdata_bits_wstrb_14 = dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@157549.4]
  assign io_dram_0_wdata_bits_wstrb_15 = dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@157550.4]
  assign io_dram_0_wdata_bits_wstrb_16 = dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@157551.4]
  assign io_dram_0_wdata_bits_wstrb_17 = dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@157552.4]
  assign io_dram_0_wdata_bits_wstrb_18 = dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@157553.4]
  assign io_dram_0_wdata_bits_wstrb_19 = dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@157554.4]
  assign io_dram_0_wdata_bits_wstrb_20 = dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@157555.4]
  assign io_dram_0_wdata_bits_wstrb_21 = dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@157556.4]
  assign io_dram_0_wdata_bits_wstrb_22 = dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@157557.4]
  assign io_dram_0_wdata_bits_wstrb_23 = dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@157558.4]
  assign io_dram_0_wdata_bits_wstrb_24 = dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@157559.4]
  assign io_dram_0_wdata_bits_wstrb_25 = dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@157560.4]
  assign io_dram_0_wdata_bits_wstrb_26 = dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@157561.4]
  assign io_dram_0_wdata_bits_wstrb_27 = dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@157562.4]
  assign io_dram_0_wdata_bits_wstrb_28 = dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@157563.4]
  assign io_dram_0_wdata_bits_wstrb_29 = dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@157564.4]
  assign io_dram_0_wdata_bits_wstrb_30 = dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@157565.4]
  assign io_dram_0_wdata_bits_wstrb_31 = dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@157566.4]
  assign io_dram_0_wdata_bits_wstrb_32 = dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@157567.4]
  assign io_dram_0_wdata_bits_wstrb_33 = dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@157568.4]
  assign io_dram_0_wdata_bits_wstrb_34 = dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@157569.4]
  assign io_dram_0_wdata_bits_wstrb_35 = dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@157570.4]
  assign io_dram_0_wdata_bits_wstrb_36 = dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@157571.4]
  assign io_dram_0_wdata_bits_wstrb_37 = dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@157572.4]
  assign io_dram_0_wdata_bits_wstrb_38 = dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@157573.4]
  assign io_dram_0_wdata_bits_wstrb_39 = dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@157574.4]
  assign io_dram_0_wdata_bits_wstrb_40 = dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@157575.4]
  assign io_dram_0_wdata_bits_wstrb_41 = dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@157576.4]
  assign io_dram_0_wdata_bits_wstrb_42 = dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@157577.4]
  assign io_dram_0_wdata_bits_wstrb_43 = dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@157578.4]
  assign io_dram_0_wdata_bits_wstrb_44 = dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@157579.4]
  assign io_dram_0_wdata_bits_wstrb_45 = dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@157580.4]
  assign io_dram_0_wdata_bits_wstrb_46 = dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@157581.4]
  assign io_dram_0_wdata_bits_wstrb_47 = dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@157582.4]
  assign io_dram_0_wdata_bits_wstrb_48 = dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@157583.4]
  assign io_dram_0_wdata_bits_wstrb_49 = dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@157584.4]
  assign io_dram_0_wdata_bits_wstrb_50 = dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@157585.4]
  assign io_dram_0_wdata_bits_wstrb_51 = dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@157586.4]
  assign io_dram_0_wdata_bits_wstrb_52 = dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@157587.4]
  assign io_dram_0_wdata_bits_wstrb_53 = dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@157588.4]
  assign io_dram_0_wdata_bits_wstrb_54 = dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@157589.4]
  assign io_dram_0_wdata_bits_wstrb_55 = dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@157590.4]
  assign io_dram_0_wdata_bits_wstrb_56 = dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@157591.4]
  assign io_dram_0_wdata_bits_wstrb_57 = dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@157592.4]
  assign io_dram_0_wdata_bits_wstrb_58 = dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@157593.4]
  assign io_dram_0_wdata_bits_wstrb_59 = dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@157594.4]
  assign io_dram_0_wdata_bits_wstrb_60 = dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@157595.4]
  assign io_dram_0_wdata_bits_wstrb_61 = dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@157596.4]
  assign io_dram_0_wdata_bits_wstrb_62 = dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@157597.4]
  assign io_dram_0_wdata_bits_wstrb_63 = dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@157598.4]
  assign io_dram_0_wdata_bits_wlast = dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@157534.4]
  assign io_dram_0_rresp_ready = dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 195:72:@157533.4]
  assign io_dram_0_wresp_ready = dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 195:72:@157466.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@153933.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@153932.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@153931.4]
  assign dramArbs_0_clock = clock; // @[:@152486.4]
  assign dramArbs_0_reset = _T_963 | reset; // @[:@152487.4 Fringe.scala 187:30:@157462.4]
  assign dramArbs_0_io_enable = _T_958 & _T_962; // @[Fringe.scala 192:36:@157463.4]
  assign dramArbs_0_io_app_loads_0_cmd_valid = io_memStreams_loads_0_cmd_valid; // @[Fringe.scala 100:70:@153650.4]
  assign dramArbs_0_io_app_loads_0_cmd_bits_addr = io_memStreams_loads_0_cmd_bits_addr; // @[Fringe.scala 100:70:@153649.4]
  assign dramArbs_0_io_app_loads_0_cmd_bits_size = io_memStreams_loads_0_cmd_bits_size; // @[Fringe.scala 100:70:@153648.4]
  assign dramArbs_0_io_app_loads_0_data_ready = io_memStreams_loads_0_data_ready; // @[Fringe.scala 100:70:@153647.4]
  assign dramArbs_0_io_app_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[Fringe.scala 101:72:@153661.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[Fringe.scala 101:72:@153660.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[Fringe.scala 101:72:@153659.4]
  assign dramArbs_0_io_app_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[Fringe.scala 101:72:@153657.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[Fringe.scala 101:72:@153656.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[Fringe.scala 101:72:@153655.4]
  assign dramArbs_0_io_app_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[Fringe.scala 101:72:@153654.4]
  assign dramArbs_0_io_dram_cmd_ready = io_dram_0_cmd_ready; // @[Fringe.scala 195:72:@157671.4]
  assign dramArbs_0_io_dram_wdata_ready = io_dram_0_wdata_ready; // @[Fringe.scala 195:72:@157664.4]
  assign dramArbs_0_io_dram_rresp_valid = io_dram_0_rresp_valid; // @[Fringe.scala 195:72:@157532.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_0 = io_dram_0_rresp_bits_rdata_0; // @[Fringe.scala 195:72:@157468.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_1 = io_dram_0_rresp_bits_rdata_1; // @[Fringe.scala 195:72:@157469.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_2 = io_dram_0_rresp_bits_rdata_2; // @[Fringe.scala 195:72:@157470.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_3 = io_dram_0_rresp_bits_rdata_3; // @[Fringe.scala 195:72:@157471.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_4 = io_dram_0_rresp_bits_rdata_4; // @[Fringe.scala 195:72:@157472.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_5 = io_dram_0_rresp_bits_rdata_5; // @[Fringe.scala 195:72:@157473.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_6 = io_dram_0_rresp_bits_rdata_6; // @[Fringe.scala 195:72:@157474.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_7 = io_dram_0_rresp_bits_rdata_7; // @[Fringe.scala 195:72:@157475.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_8 = io_dram_0_rresp_bits_rdata_8; // @[Fringe.scala 195:72:@157476.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_9 = io_dram_0_rresp_bits_rdata_9; // @[Fringe.scala 195:72:@157477.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_10 = io_dram_0_rresp_bits_rdata_10; // @[Fringe.scala 195:72:@157478.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_11 = io_dram_0_rresp_bits_rdata_11; // @[Fringe.scala 195:72:@157479.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_12 = io_dram_0_rresp_bits_rdata_12; // @[Fringe.scala 195:72:@157480.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_13 = io_dram_0_rresp_bits_rdata_13; // @[Fringe.scala 195:72:@157481.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_14 = io_dram_0_rresp_bits_rdata_14; // @[Fringe.scala 195:72:@157482.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_15 = io_dram_0_rresp_bits_rdata_15; // @[Fringe.scala 195:72:@157483.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_16 = io_dram_0_rresp_bits_rdata_16; // @[Fringe.scala 195:72:@157484.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_17 = io_dram_0_rresp_bits_rdata_17; // @[Fringe.scala 195:72:@157485.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_18 = io_dram_0_rresp_bits_rdata_18; // @[Fringe.scala 195:72:@157486.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_19 = io_dram_0_rresp_bits_rdata_19; // @[Fringe.scala 195:72:@157487.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_20 = io_dram_0_rresp_bits_rdata_20; // @[Fringe.scala 195:72:@157488.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_21 = io_dram_0_rresp_bits_rdata_21; // @[Fringe.scala 195:72:@157489.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_22 = io_dram_0_rresp_bits_rdata_22; // @[Fringe.scala 195:72:@157490.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_23 = io_dram_0_rresp_bits_rdata_23; // @[Fringe.scala 195:72:@157491.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_24 = io_dram_0_rresp_bits_rdata_24; // @[Fringe.scala 195:72:@157492.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_25 = io_dram_0_rresp_bits_rdata_25; // @[Fringe.scala 195:72:@157493.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_26 = io_dram_0_rresp_bits_rdata_26; // @[Fringe.scala 195:72:@157494.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_27 = io_dram_0_rresp_bits_rdata_27; // @[Fringe.scala 195:72:@157495.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_28 = io_dram_0_rresp_bits_rdata_28; // @[Fringe.scala 195:72:@157496.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_29 = io_dram_0_rresp_bits_rdata_29; // @[Fringe.scala 195:72:@157497.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_30 = io_dram_0_rresp_bits_rdata_30; // @[Fringe.scala 195:72:@157498.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_31 = io_dram_0_rresp_bits_rdata_31; // @[Fringe.scala 195:72:@157499.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_32 = io_dram_0_rresp_bits_rdata_32; // @[Fringe.scala 195:72:@157500.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_33 = io_dram_0_rresp_bits_rdata_33; // @[Fringe.scala 195:72:@157501.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_34 = io_dram_0_rresp_bits_rdata_34; // @[Fringe.scala 195:72:@157502.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_35 = io_dram_0_rresp_bits_rdata_35; // @[Fringe.scala 195:72:@157503.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_36 = io_dram_0_rresp_bits_rdata_36; // @[Fringe.scala 195:72:@157504.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_37 = io_dram_0_rresp_bits_rdata_37; // @[Fringe.scala 195:72:@157505.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_38 = io_dram_0_rresp_bits_rdata_38; // @[Fringe.scala 195:72:@157506.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_39 = io_dram_0_rresp_bits_rdata_39; // @[Fringe.scala 195:72:@157507.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_40 = io_dram_0_rresp_bits_rdata_40; // @[Fringe.scala 195:72:@157508.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_41 = io_dram_0_rresp_bits_rdata_41; // @[Fringe.scala 195:72:@157509.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_42 = io_dram_0_rresp_bits_rdata_42; // @[Fringe.scala 195:72:@157510.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_43 = io_dram_0_rresp_bits_rdata_43; // @[Fringe.scala 195:72:@157511.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_44 = io_dram_0_rresp_bits_rdata_44; // @[Fringe.scala 195:72:@157512.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_45 = io_dram_0_rresp_bits_rdata_45; // @[Fringe.scala 195:72:@157513.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_46 = io_dram_0_rresp_bits_rdata_46; // @[Fringe.scala 195:72:@157514.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_47 = io_dram_0_rresp_bits_rdata_47; // @[Fringe.scala 195:72:@157515.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_48 = io_dram_0_rresp_bits_rdata_48; // @[Fringe.scala 195:72:@157516.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_49 = io_dram_0_rresp_bits_rdata_49; // @[Fringe.scala 195:72:@157517.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_50 = io_dram_0_rresp_bits_rdata_50; // @[Fringe.scala 195:72:@157518.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_51 = io_dram_0_rresp_bits_rdata_51; // @[Fringe.scala 195:72:@157519.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_52 = io_dram_0_rresp_bits_rdata_52; // @[Fringe.scala 195:72:@157520.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_53 = io_dram_0_rresp_bits_rdata_53; // @[Fringe.scala 195:72:@157521.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_54 = io_dram_0_rresp_bits_rdata_54; // @[Fringe.scala 195:72:@157522.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_55 = io_dram_0_rresp_bits_rdata_55; // @[Fringe.scala 195:72:@157523.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_56 = io_dram_0_rresp_bits_rdata_56; // @[Fringe.scala 195:72:@157524.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_57 = io_dram_0_rresp_bits_rdata_57; // @[Fringe.scala 195:72:@157525.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_58 = io_dram_0_rresp_bits_rdata_58; // @[Fringe.scala 195:72:@157526.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_59 = io_dram_0_rresp_bits_rdata_59; // @[Fringe.scala 195:72:@157527.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_60 = io_dram_0_rresp_bits_rdata_60; // @[Fringe.scala 195:72:@157528.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_61 = io_dram_0_rresp_bits_rdata_61; // @[Fringe.scala 195:72:@157529.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_62 = io_dram_0_rresp_bits_rdata_62; // @[Fringe.scala 195:72:@157530.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_63 = io_dram_0_rresp_bits_rdata_63; // @[Fringe.scala 195:72:@157531.4]
  assign dramArbs_0_io_dram_rresp_bits_tag = io_dram_0_rresp_bits_tag; // @[Fringe.scala 195:72:@157467.4]
  assign dramArbs_0_io_dram_wresp_valid = io_dram_0_wresp_valid; // @[Fringe.scala 195:72:@157465.4]
  assign dramArbs_0_io_dram_wresp_bits_tag = io_dram_0_wresp_bits_tag; // @[Fringe.scala 195:72:@157464.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@153936.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@153935.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@153934.4]
  assign heap_io_host_0_resp_valid = _T_1502 & _T_1506; // @[Fringe.scala 204:22:@157679.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@157680.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@157681.4]
  assign regs_clock = clock; // @[:@153938.4]
  assign regs_reset = reset; // @[:@153939.4 Fringe.scala 139:14:@156226.4]
  assign regs_io_raddr = io_raddr[10:0]; // @[Fringe.scala 118:17:@156194.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@156196.4]
  assign regs_io_waddr = io_waddr[10:0]; // @[Fringe.scala 119:17:@156195.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@156197.4]
  assign regs_io_reset = _T_963 | reset; // @[Fringe.scala 138:17:@156224.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_982; // @[Fringe.scala 170:23:@156276.4]
  assign regs_io_argOuts_0_bits = {_T_998,_T_997}; // @[Fringe.scala 171:22:@156280.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@156283.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@156282.4]
  assign regs_io_argOuts_2_valid = io_argOuts_1_valid; // @[Fringe.scala 176:23:@156286.4]
  assign regs_io_argOuts_2_bits = io_argOuts_1_bits; // @[Fringe.scala 175:22:@156285.4]
  assign regs_io_argOuts_3_valid = io_argOuts_2_valid; // @[Fringe.scala 176:23:@156289.4]
  assign regs_io_argOuts_3_bits = io_argOuts_2_bits; // @[Fringe.scala 175:22:@156288.4]
  assign regs_io_argOuts_4_valid = io_argOuts_3_valid; // @[Fringe.scala 176:23:@156292.4]
  assign regs_io_argOuts_4_bits = io_argOuts_3_bits; // @[Fringe.scala 175:22:@156291.4]
  assign regs_io_argOuts_5_valid = io_argOuts_4_valid; // @[Fringe.scala 176:23:@156295.4]
  assign regs_io_argOuts_5_bits = io_argOuts_4_bits; // @[Fringe.scala 175:22:@156294.4]
  assign regs_io_argOuts_6_valid = io_argOuts_5_valid; // @[Fringe.scala 176:23:@156298.4]
  assign regs_io_argOuts_6_bits = io_argOuts_5_bits; // @[Fringe.scala 175:22:@156297.4]
  assign regs_io_argOuts_7_valid = io_argOuts_6_valid; // @[Fringe.scala 176:23:@156301.4]
  assign regs_io_argOuts_7_bits = io_argOuts_6_bits; // @[Fringe.scala 175:22:@156300.4]
  assign regs_io_argOuts_8_valid = io_argOuts_7_valid; // @[Fringe.scala 176:23:@156304.4]
  assign regs_io_argOuts_8_bits = io_argOuts_7_bits; // @[Fringe.scala 175:22:@156303.4]
  assign regs_io_argOuts_9_valid = io_argOuts_8_valid; // @[Fringe.scala 176:23:@156307.4]
  assign regs_io_argOuts_9_bits = io_argOuts_8_bits; // @[Fringe.scala 175:22:@156306.4]
  assign regs_io_argOuts_10_valid = io_argOuts_9_valid; // @[Fringe.scala 176:23:@156310.4]
  assign regs_io_argOuts_10_bits = io_argOuts_9_bits; // @[Fringe.scala 175:22:@156309.4]
  assign regs_io_argOuts_11_valid = io_argOuts_10_valid; // @[Fringe.scala 176:23:@156313.4]
  assign regs_io_argOuts_11_bits = io_argOuts_10_bits; // @[Fringe.scala 175:22:@156312.4]
  assign regs_io_argOuts_12_valid = io_argOuts_11_valid; // @[Fringe.scala 176:23:@156316.4]
  assign regs_io_argOuts_12_bits = io_argOuts_11_bits; // @[Fringe.scala 175:22:@156315.4]
  assign regs_io_argOuts_13_valid = io_argOuts_12_valid; // @[Fringe.scala 176:23:@156319.4]
  assign regs_io_argOuts_13_bits = io_argOuts_12_bits; // @[Fringe.scala 175:22:@156318.4]
  assign regs_io_argOuts_14_valid = io_argOuts_13_valid; // @[Fringe.scala 176:23:@156322.4]
  assign regs_io_argOuts_14_bits = io_argOuts_13_bits; // @[Fringe.scala 175:22:@156321.4]
  assign regs_io_argOuts_15_valid = io_argOuts_14_valid; // @[Fringe.scala 176:23:@156325.4]
  assign regs_io_argOuts_15_bits = io_argOuts_14_bits; // @[Fringe.scala 175:22:@156324.4]
  assign regs_io_argOuts_16_valid = io_argOuts_15_valid; // @[Fringe.scala 176:23:@156328.4]
  assign regs_io_argOuts_16_bits = io_argOuts_15_bits; // @[Fringe.scala 175:22:@156327.4]
  assign regs_io_argOuts_17_valid = io_argOuts_16_valid; // @[Fringe.scala 176:23:@156331.4]
  assign regs_io_argOuts_17_bits = io_argOuts_16_bits; // @[Fringe.scala 175:22:@156330.4]
  assign regs_io_argOuts_18_valid = io_argOuts_17_valid; // @[Fringe.scala 176:23:@156334.4]
  assign regs_io_argOuts_18_bits = io_argOuts_17_bits; // @[Fringe.scala 175:22:@156333.4]
  assign regs_io_argOuts_19_valid = io_argOuts_18_valid; // @[Fringe.scala 176:23:@156337.4]
  assign regs_io_argOuts_19_bits = io_argOuts_18_bits; // @[Fringe.scala 175:22:@156336.4]
  assign regs_io_argOuts_20_valid = io_argOuts_19_valid; // @[Fringe.scala 176:23:@156340.4]
  assign regs_io_argOuts_20_bits = io_argOuts_19_bits; // @[Fringe.scala 175:22:@156339.4]
  assign regs_io_argOuts_21_valid = io_argOuts_20_valid; // @[Fringe.scala 176:23:@156343.4]
  assign regs_io_argOuts_21_bits = io_argOuts_20_bits; // @[Fringe.scala 175:22:@156342.4]
  assign regs_io_argOuts_22_valid = io_argOuts_21_valid; // @[Fringe.scala 176:23:@156346.4]
  assign regs_io_argOuts_22_bits = io_argOuts_21_bits; // @[Fringe.scala 175:22:@156345.4]
  assign regs_io_argOuts_23_valid = io_argOuts_22_valid; // @[Fringe.scala 176:23:@156349.4]
  assign regs_io_argOuts_23_bits = io_argOuts_22_bits; // @[Fringe.scala 175:22:@156348.4]
  assign regs_io_argOuts_24_valid = io_argOuts_23_valid; // @[Fringe.scala 176:23:@156352.4]
  assign regs_io_argOuts_24_bits = io_argOuts_23_bits; // @[Fringe.scala 175:22:@156351.4]
  assign regs_io_argOuts_25_valid = io_argOuts_24_valid; // @[Fringe.scala 176:23:@156355.4]
  assign regs_io_argOuts_25_bits = io_argOuts_24_bits; // @[Fringe.scala 175:22:@156354.4]
  assign regs_io_argOuts_26_valid = io_argOuts_25_valid; // @[Fringe.scala 176:23:@156358.4]
  assign regs_io_argOuts_26_bits = io_argOuts_25_bits; // @[Fringe.scala 175:22:@156357.4]
  assign regs_io_argOuts_27_valid = io_argOuts_26_valid; // @[Fringe.scala 176:23:@156361.4]
  assign regs_io_argOuts_27_bits = io_argOuts_26_bits; // @[Fringe.scala 175:22:@156360.4]
  assign regs_io_argOuts_28_valid = io_argOuts_27_valid; // @[Fringe.scala 176:23:@156364.4]
  assign regs_io_argOuts_28_bits = io_argOuts_27_bits; // @[Fringe.scala 175:22:@156363.4]
  assign regs_io_argOuts_29_valid = io_argOuts_28_valid; // @[Fringe.scala 176:23:@156367.4]
  assign regs_io_argOuts_29_bits = io_argOuts_28_bits; // @[Fringe.scala 175:22:@156366.4]
  assign regs_io_argOuts_30_valid = io_argOuts_29_valid; // @[Fringe.scala 176:23:@156370.4]
  assign regs_io_argOuts_30_bits = io_argOuts_29_bits; // @[Fringe.scala 175:22:@156369.4]
  assign regs_io_argOuts_31_valid = io_argOuts_30_valid; // @[Fringe.scala 176:23:@156373.4]
  assign regs_io_argOuts_31_bits = io_argOuts_30_bits; // @[Fringe.scala 175:22:@156372.4]
  assign regs_io_argOuts_32_valid = io_argOuts_31_valid; // @[Fringe.scala 176:23:@156376.4]
  assign regs_io_argOuts_32_bits = io_argOuts_31_bits; // @[Fringe.scala 175:22:@156375.4]
  assign regs_io_argOuts_33_valid = io_argOuts_32_valid; // @[Fringe.scala 176:23:@156379.4]
  assign regs_io_argOuts_33_bits = io_argOuts_32_bits; // @[Fringe.scala 175:22:@156378.4]
  assign regs_io_argOuts_34_valid = io_argOuts_33_valid; // @[Fringe.scala 176:23:@156382.4]
  assign regs_io_argOuts_34_bits = io_argOuts_33_bits; // @[Fringe.scala 175:22:@156381.4]
  assign regs_io_argOuts_35_valid = io_argOuts_34_valid; // @[Fringe.scala 176:23:@156385.4]
  assign regs_io_argOuts_35_bits = io_argOuts_34_bits; // @[Fringe.scala 175:22:@156384.4]
  assign regs_io_argOuts_36_valid = io_argOuts_35_valid; // @[Fringe.scala 176:23:@156388.4]
  assign regs_io_argOuts_36_bits = io_argOuts_35_bits; // @[Fringe.scala 175:22:@156387.4]
  assign regs_io_argOuts_37_valid = io_argOuts_36_valid; // @[Fringe.scala 176:23:@156391.4]
  assign regs_io_argOuts_37_bits = io_argOuts_36_bits; // @[Fringe.scala 175:22:@156390.4]
  assign regs_io_argOuts_38_valid = io_argOuts_37_valid; // @[Fringe.scala 176:23:@156394.4]
  assign regs_io_argOuts_38_bits = io_argOuts_37_bits; // @[Fringe.scala 175:22:@156393.4]
  assign regs_io_argOuts_39_valid = io_argOuts_38_valid; // @[Fringe.scala 176:23:@156397.4]
  assign regs_io_argOuts_39_bits = io_argOuts_38_bits; // @[Fringe.scala 175:22:@156396.4]
  assign regs_io_argOuts_40_valid = io_argOuts_39_valid; // @[Fringe.scala 176:23:@156400.4]
  assign regs_io_argOuts_40_bits = io_argOuts_39_bits; // @[Fringe.scala 175:22:@156399.4]
  assign regs_io_argOuts_41_valid = io_argOuts_40_valid; // @[Fringe.scala 176:23:@156403.4]
  assign regs_io_argOuts_41_bits = io_argOuts_40_bits; // @[Fringe.scala 175:22:@156402.4]
  assign regs_io_argOuts_42_valid = io_argOuts_41_valid; // @[Fringe.scala 176:23:@156406.4]
  assign regs_io_argOuts_42_bits = io_argOuts_41_bits; // @[Fringe.scala 175:22:@156405.4]
  assign regs_io_argOuts_43_valid = io_argOuts_42_valid; // @[Fringe.scala 176:23:@156409.4]
  assign regs_io_argOuts_43_bits = io_argOuts_42_bits; // @[Fringe.scala 175:22:@156408.4]
  assign regs_io_argOuts_44_valid = io_argOuts_43_valid; // @[Fringe.scala 176:23:@156412.4]
  assign regs_io_argOuts_44_bits = io_argOuts_43_bits; // @[Fringe.scala 175:22:@156411.4]
  assign regs_io_argOuts_45_valid = io_argOuts_44_valid; // @[Fringe.scala 176:23:@156415.4]
  assign regs_io_argOuts_45_bits = io_argOuts_44_bits; // @[Fringe.scala 175:22:@156414.4]
  assign regs_io_argOuts_46_valid = io_argOuts_45_valid; // @[Fringe.scala 176:23:@156418.4]
  assign regs_io_argOuts_46_bits = io_argOuts_45_bits; // @[Fringe.scala 175:22:@156417.4]
  assign regs_io_argOuts_47_valid = io_argOuts_46_valid; // @[Fringe.scala 176:23:@156421.4]
  assign regs_io_argOuts_47_bits = io_argOuts_46_bits; // @[Fringe.scala 175:22:@156420.4]
  assign regs_io_argOuts_48_valid = io_argOuts_47_valid; // @[Fringe.scala 176:23:@156424.4]
  assign regs_io_argOuts_48_bits = io_argOuts_47_bits; // @[Fringe.scala 175:22:@156423.4]
  assign regs_io_argOuts_49_valid = io_argOuts_48_valid; // @[Fringe.scala 176:23:@156427.4]
  assign regs_io_argOuts_49_bits = io_argOuts_48_bits; // @[Fringe.scala 175:22:@156426.4]
  assign regs_io_argOuts_50_valid = io_argOuts_49_valid; // @[Fringe.scala 176:23:@156430.4]
  assign regs_io_argOuts_50_bits = io_argOuts_49_bits; // @[Fringe.scala 175:22:@156429.4]
  assign regs_io_argOuts_51_valid = io_argOuts_50_valid; // @[Fringe.scala 176:23:@156433.4]
  assign regs_io_argOuts_51_bits = io_argOuts_50_bits; // @[Fringe.scala 175:22:@156432.4]
  assign regs_io_argOuts_52_valid = io_argOuts_51_valid; // @[Fringe.scala 176:23:@156436.4]
  assign regs_io_argOuts_52_bits = io_argOuts_51_bits; // @[Fringe.scala 175:22:@156435.4]
  assign regs_io_argOuts_53_valid = io_argOuts_52_valid; // @[Fringe.scala 176:23:@156439.4]
  assign regs_io_argOuts_53_bits = io_argOuts_52_bits; // @[Fringe.scala 175:22:@156438.4]
  assign regs_io_argOuts_54_valid = io_argOuts_53_valid; // @[Fringe.scala 176:23:@156442.4]
  assign regs_io_argOuts_54_bits = io_argOuts_53_bits; // @[Fringe.scala 175:22:@156441.4]
  assign regs_io_argOuts_55_valid = io_argOuts_54_valid; // @[Fringe.scala 176:23:@156445.4]
  assign regs_io_argOuts_55_bits = io_argOuts_54_bits; // @[Fringe.scala 175:22:@156444.4]
  assign regs_io_argOuts_56_valid = io_argOuts_55_valid; // @[Fringe.scala 176:23:@156448.4]
  assign regs_io_argOuts_56_bits = io_argOuts_55_bits; // @[Fringe.scala 175:22:@156447.4]
  assign regs_io_argOuts_57_valid = io_argOuts_56_valid; // @[Fringe.scala 176:23:@156451.4]
  assign regs_io_argOuts_57_bits = io_argOuts_56_bits; // @[Fringe.scala 175:22:@156450.4]
  assign regs_io_argOuts_58_valid = io_argOuts_57_valid; // @[Fringe.scala 176:23:@156454.4]
  assign regs_io_argOuts_58_bits = io_argOuts_57_bits; // @[Fringe.scala 175:22:@156453.4]
  assign regs_io_argOuts_59_valid = io_argOuts_58_valid; // @[Fringe.scala 176:23:@156457.4]
  assign regs_io_argOuts_59_bits = io_argOuts_58_bits; // @[Fringe.scala 175:22:@156456.4]
  assign regs_io_argOuts_60_valid = io_argOuts_59_valid; // @[Fringe.scala 176:23:@156460.4]
  assign regs_io_argOuts_60_bits = io_argOuts_59_bits; // @[Fringe.scala 175:22:@156459.4]
  assign regs_io_argOuts_61_bits = {{32'd0}, dramArbs_0_io_debugSignals_0}; // @[Fringe.scala 179:22:@156461.4]
  assign regs_io_argOuts_62_bits = {{32'd0}, dramArbs_0_io_debugSignals_1}; // @[Fringe.scala 179:22:@156463.4]
  assign regs_io_argOuts_63_bits = {{32'd0}, dramArbs_0_io_debugSignals_2}; // @[Fringe.scala 179:22:@156465.4]
  assign regs_io_argOuts_64_bits = {{32'd0}, dramArbs_0_io_debugSignals_3}; // @[Fringe.scala 179:22:@156467.4]
  assign regs_io_argOuts_65_bits = {{32'd0}, dramArbs_0_io_debugSignals_4}; // @[Fringe.scala 179:22:@156469.4]
  assign regs_io_argOuts_66_bits = {{32'd0}, dramArbs_0_io_debugSignals_5}; // @[Fringe.scala 179:22:@156471.4]
  assign regs_io_argOuts_67_bits = {{32'd0}, dramArbs_0_io_debugSignals_6}; // @[Fringe.scala 179:22:@156473.4]
  assign regs_io_argOuts_68_bits = {{32'd0}, dramArbs_0_io_debugSignals_7}; // @[Fringe.scala 179:22:@156475.4]
  assign regs_io_argOuts_69_bits = {{32'd0}, dramArbs_0_io_debugSignals_8}; // @[Fringe.scala 179:22:@156477.4]
  assign regs_io_argOuts_70_bits = {{32'd0}, dramArbs_0_io_debugSignals_9}; // @[Fringe.scala 179:22:@156479.4]
  assign regs_io_argOuts_71_bits = {{32'd0}, dramArbs_0_io_debugSignals_10}; // @[Fringe.scala 179:22:@156481.4]
  assign regs_io_argOuts_72_bits = {{32'd0}, dramArbs_0_io_debugSignals_11}; // @[Fringe.scala 179:22:@156483.4]
  assign regs_io_argOuts_73_bits = {{32'd0}, dramArbs_0_io_debugSignals_12}; // @[Fringe.scala 179:22:@156485.4]
  assign regs_io_argOuts_74_bits = {{32'd0}, dramArbs_0_io_debugSignals_13}; // @[Fringe.scala 179:22:@156487.4]
  assign regs_io_argOuts_75_bits = {{32'd0}, dramArbs_0_io_debugSignals_14}; // @[Fringe.scala 179:22:@156489.4]
  assign regs_io_argOuts_76_bits = {{32'd0}, dramArbs_0_io_debugSignals_15}; // @[Fringe.scala 179:22:@156491.4]
  assign regs_io_argOuts_77_bits = {{32'd0}, dramArbs_0_io_debugSignals_16}; // @[Fringe.scala 179:22:@156493.4]
  assign regs_io_argOuts_78_bits = {{32'd0}, dramArbs_0_io_debugSignals_17}; // @[Fringe.scala 179:22:@156495.4]
  assign regs_io_argOuts_79_bits = {{32'd0}, dramArbs_0_io_debugSignals_18}; // @[Fringe.scala 179:22:@156497.4]
  assign regs_io_argOuts_80_bits = {{32'd0}, dramArbs_0_io_debugSignals_19}; // @[Fringe.scala 179:22:@156499.4]
  assign regs_io_argOuts_81_bits = {{32'd0}, dramArbs_0_io_debugSignals_20}; // @[Fringe.scala 179:22:@156501.4]
  assign regs_io_argOuts_82_bits = {{32'd0}, dramArbs_0_io_debugSignals_21}; // @[Fringe.scala 179:22:@156503.4]
  assign regs_io_argOuts_83_bits = {{32'd0}, dramArbs_0_io_debugSignals_22}; // @[Fringe.scala 179:22:@156505.4]
  assign regs_io_argOuts_84_bits = {{32'd0}, dramArbs_0_io_debugSignals_23}; // @[Fringe.scala 179:22:@156507.4]
  assign regs_io_argOuts_85_bits = {{32'd0}, dramArbs_0_io_debugSignals_24}; // @[Fringe.scala 179:22:@156509.4]
  assign regs_io_argOuts_86_bits = {{32'd0}, dramArbs_0_io_debugSignals_25}; // @[Fringe.scala 179:22:@156511.4]
  assign regs_io_argOuts_87_bits = {{32'd0}, dramArbs_0_io_debugSignals_26}; // @[Fringe.scala 179:22:@156513.4]
  assign regs_io_argOuts_88_bits = {{32'd0}, dramArbs_0_io_debugSignals_27}; // @[Fringe.scala 179:22:@156515.4]
  assign regs_io_argOuts_89_bits = {{32'd0}, dramArbs_0_io_debugSignals_28}; // @[Fringe.scala 179:22:@156517.4]
  assign regs_io_argOuts_90_bits = {{32'd0}, dramArbs_0_io_debugSignals_29}; // @[Fringe.scala 179:22:@156519.4]
  assign regs_io_argOuts_91_bits = {{32'd0}, dramArbs_0_io_debugSignals_30}; // @[Fringe.scala 179:22:@156521.4]
  assign regs_io_argOuts_102_bits = {{32'd0}, dramArbs_0_io_debugSignals_41}; // @[Fringe.scala 179:22:@156543.4]
  assign timeoutCtr_clock = clock; // @[:@156228.4]
  assign timeoutCtr_reset = reset; // @[:@156229.4]
  assign timeoutCtr_io_enable = _T_958 & _T_962; // @[Fringe.scala 149:24:@156243.4]
  assign depulser_clock = clock; // @[:@156247.4]
  assign depulser_reset = reset; // @[:@156248.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@156253.4]
  assign depulser_io_rst = _T_973[0]; // @[Fringe.scala 156:19:@156255.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_949 = _RAND_0[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_980 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1505 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    _T_949 <= regs_io_rdata;
    if (reset) begin
      _T_980 <= 1'h0;
    end else begin
      _T_980 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1505 <= 1'h0;
    end else begin
      _T_1505 <= _T_1502;
    end
  end
endmodule
module SpatialIP( // @[:@157683.2]
  input         clock, // @[:@157684.4]
  input         reset, // @[:@157685.4]
  input  [31:0] io_raddr, // @[:@157686.4]
  input         io_wen, // @[:@157686.4]
  input  [31:0] io_waddr, // @[:@157686.4]
  input  [63:0] io_wdata, // @[:@157686.4]
  output [63:0] io_rdata, // @[:@157686.4]
  input         io_dram_0_cmd_ready, // @[:@157686.4]
  output        io_dram_0_cmd_valid, // @[:@157686.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@157686.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@157686.4]
  output [63:0] io_dram_0_cmd_bits_rawAddr, // @[:@157686.4]
  output        io_dram_0_cmd_bits_isWr, // @[:@157686.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@157686.4]
  input         io_dram_0_wdata_ready, // @[:@157686.4]
  output        io_dram_0_wdata_valid, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_0, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_1, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_2, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_3, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_4, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_5, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_6, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_7, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_8, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_9, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_10, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_11, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_12, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_13, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_14, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_15, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_16, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_17, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_18, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_19, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_20, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_21, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_22, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_23, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_24, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_25, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_26, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_27, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_28, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_29, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_30, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_31, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_32, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_33, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_34, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_35, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_36, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_37, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_38, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_39, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_40, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_41, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_42, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_43, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_44, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_45, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_46, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_47, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_48, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_49, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_50, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_51, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_52, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_53, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_54, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_55, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_56, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_57, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_58, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_59, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_60, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_61, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_62, // @[:@157686.4]
  output [7:0]  io_dram_0_wdata_bits_wdata_63, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_0, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_1, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_2, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_3, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_4, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_5, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_6, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_7, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_8, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_9, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_10, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_11, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_12, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_13, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_14, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_15, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_16, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_17, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_18, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_19, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_20, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_21, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_22, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_23, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_24, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_25, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_26, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_27, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_28, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_29, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_30, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_31, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_32, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_33, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_34, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_35, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_36, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_37, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_38, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_39, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_40, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_41, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_42, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_43, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_44, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_45, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_46, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_47, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_48, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_49, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_50, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_51, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_52, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_53, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_54, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_55, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_56, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_57, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_58, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_59, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_60, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_61, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_62, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wstrb_63, // @[:@157686.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@157686.4]
  output        io_dram_0_rresp_ready, // @[:@157686.4]
  input         io_dram_0_rresp_valid, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_0, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_1, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_2, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_3, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_4, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_5, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_6, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_7, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_8, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_9, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_10, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_11, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_12, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_13, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_14, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_15, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_16, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_17, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_18, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_19, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_20, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_21, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_22, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_23, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_24, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_25, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_26, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_27, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_28, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_29, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_30, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_31, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_32, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_33, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_34, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_35, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_36, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_37, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_38, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_39, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_40, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_41, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_42, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_43, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_44, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_45, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_46, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_47, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_48, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_49, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_50, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_51, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_52, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_53, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_54, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_55, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_56, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_57, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_58, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_59, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_60, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_61, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_62, // @[:@157686.4]
  input  [7:0]  io_dram_0_rresp_bits_rdata_63, // @[:@157686.4]
  input  [31:0] io_dram_0_rresp_bits_tag, // @[:@157686.4]
  output        io_dram_0_wresp_ready, // @[:@157686.4]
  input         io_dram_0_wresp_valid, // @[:@157686.4]
  input  [31:0] io_dram_0_wresp_bits_tag // @[:@157686.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@157688.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@157688.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_16; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_17; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_18; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_19; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_20; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_21; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_22; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_23; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_24; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_25; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_26; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_27; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_28; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_29; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_30; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_31; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_32; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_33; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_34; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_35; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_36; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_37; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_38; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_39; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_40; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_41; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_42; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_43; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_44; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_45; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_46; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_47; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_48; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_49; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_50; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_51; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_52; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_53; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_54; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_55; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_56; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_57; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_58; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_59; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_60; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_61; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_62; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_63; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_16; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_17; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_18; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_19; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_20; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_21; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_22; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_23; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_24; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_25; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_26; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_27; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_28; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_29; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_30; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_31; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_32; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_33; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_34; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_35; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_36; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_37; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_38; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_39; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_40; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_41; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_42; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_43; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_44; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_45; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_46; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_47; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_48; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_49; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_50; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_51; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_52; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_53; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_54; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_55; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_56; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_57; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_58; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_59; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_60; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_61; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_62; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_gathers_0_data_bits_63; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_16; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_17; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_18; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_19; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_20; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_21; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_22; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_23; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_24; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_25; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_26; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_27; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_28; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_29; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_30; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_31; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_32; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_33; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_34; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_35; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_36; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_37; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_38; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_39; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_40; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_41; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_42; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_43; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_44; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_45; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_46; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_47; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_48; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_49; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_50; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_51; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_52; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_53; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_54; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_55; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_56; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_57; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_58; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_59; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_60; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_61; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_62; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_63; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_16; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_17; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_18; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_19; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_20; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_21; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_22; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_23; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_24; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_25; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_26; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_27; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_28; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_29; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_30; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_31; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_32; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_33; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_34; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_35; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_36; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_37; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_38; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_39; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_40; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_41; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_42; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_43; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_44; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_45; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_46; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_47; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_48; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_49; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_50; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_51; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_52; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_53; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_54; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_55; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_56; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_57; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_58; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_59; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_60; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_61; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_62; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_63; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@157688.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@157688.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@157688.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@157688.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@157688.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@157688.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@157688.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@157688.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@157688.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_1_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_1_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_1_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_1_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_2_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_2_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_2_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_2_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_3_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_3_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_3_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_3_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_4_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_4_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_4_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_4_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_5_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_5_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_5_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_5_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_6_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_6_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_6_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_6_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_7_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_7_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_7_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_7_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_8_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_8_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_8_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_8_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_9_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_9_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_9_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_9_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_10_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_10_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_10_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_10_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_11_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_11_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_11_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_11_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_12_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_12_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_12_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_12_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_13_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_13_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_13_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_13_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_14_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_14_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_14_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_14_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_15_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_15_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_15_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_15_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_16_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_16_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_16_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_16_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_17_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_17_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_17_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_17_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_18_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_18_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_18_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_18_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_19_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_19_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_19_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_19_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_20_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_20_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_20_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_20_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_21_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_21_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_21_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_21_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_22_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_22_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_22_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_22_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_23_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_23_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_23_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_23_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_24_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_24_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_24_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_24_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_25_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_25_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_25_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_25_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_26_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_26_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_26_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_26_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_27_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_27_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_27_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_27_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_28_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_28_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_28_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_28_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_29_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_29_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_29_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_29_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_30_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_30_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_30_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_30_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_31_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_31_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_31_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_31_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_32_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_32_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_32_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_32_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_33_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_33_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_33_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_33_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_34_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_34_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_34_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_34_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_35_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_35_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_35_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_35_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_36_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_36_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_36_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_36_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_37_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_37_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_37_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_37_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_38_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_38_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_38_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_38_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_39_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_39_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_39_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_39_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_40_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_40_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_40_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_40_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_41_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_41_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_41_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_41_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_42_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_42_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_42_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_42_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_43_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_43_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_43_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_43_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_44_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_44_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_44_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_44_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_45_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_45_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_45_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_45_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_46_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_46_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_46_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_46_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_47_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_47_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_47_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_47_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_48_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_48_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_48_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_48_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_49_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_49_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_49_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_49_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_50_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_50_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_50_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_50_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_51_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_51_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_51_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_51_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_52_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_52_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_52_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_52_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_53_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_53_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_53_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_53_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_54_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_54_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_54_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_54_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_55_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_55_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_55_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_55_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_56_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_56_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_56_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_56_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_57_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_57_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_57_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_57_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_58_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_58_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_58_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_58_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_59_port_ready; // @[Instantiator.scala 53:44:@157688.4]
  wire  accel_io_argOuts_59_port_valid; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_59_port_bits; // @[Instantiator.scala 53:44:@157688.4]
  wire [63:0] accel_io_argOuts_59_echo; // @[Instantiator.scala 53:44:@157688.4]
  wire  Fringe_clock; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_reset; // @[SimTarget.scala 16:24:@158243.4]
  wire [31:0] Fringe_io_raddr; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_wen; // @[SimTarget.scala 16:24:@158243.4]
  wire [31:0] Fringe_io_waddr; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_wdata; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_rdata; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_enable; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_done; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_reset; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argIns_0; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argIns_1; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_0_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_0_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_1_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_1_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_2_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_2_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_3_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_3_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_4_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_4_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_5_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_5_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_6_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_6_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_7_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_7_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_8_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_8_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_9_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_9_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_10_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_10_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_11_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_11_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_12_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_12_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_13_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_13_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_14_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_14_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_15_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_15_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_16_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_16_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_17_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_17_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_18_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_18_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_19_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_19_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_20_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_20_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_21_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_21_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_22_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_22_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_23_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_23_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_24_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_24_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_25_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_25_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_26_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_26_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_27_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_27_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_28_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_28_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_29_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_29_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_30_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_30_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_31_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_31_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_32_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_32_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_33_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_33_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_34_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_34_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_35_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_35_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_36_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_36_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_37_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_37_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_38_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_38_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_39_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_39_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_40_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_40_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_41_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_41_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_42_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_42_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_43_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_43_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_44_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_44_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_45_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_45_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_46_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_46_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_47_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_47_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_48_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_48_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_49_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_49_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_50_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_50_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_51_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_51_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_52_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_52_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_53_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_53_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_54_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_54_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_55_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_55_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_56_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_56_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_57_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_57_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_58_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_58_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_argOuts_59_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argOuts_59_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_0; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_1; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_2; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_3; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_4; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_5; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_6; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_7; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_8; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_9; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_10; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_11; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_12; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_13; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_14; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_15; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_16; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_17; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_18; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_19; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_20; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_21; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_22; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_23; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_24; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_25; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_26; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_27; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_28; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_29; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_30; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_31; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_32; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_33; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_34; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_35; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_36; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_37; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_38; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_39; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_40; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_41; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_42; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_43; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_44; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_45; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_46; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_47; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_48; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_49; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_50; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_51; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_52; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_53; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_54; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_55; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_56; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_57; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_58; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_argEchos_59; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_memStreams_loads_0_cmd_ready; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_memStreams_loads_0_cmd_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_memStreams_loads_0_cmd_bits_addr; // @[SimTarget.scala 16:24:@158243.4]
  wire [31:0] Fringe_io_memStreams_loads_0_cmd_bits_size; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_memStreams_loads_0_data_ready; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_memStreams_loads_0_data_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [31:0] Fringe_io_memStreams_loads_0_data_bits_rdata_0; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_memStreams_stores_0_cmd_ready; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_memStreams_stores_0_cmd_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_memStreams_stores_0_cmd_bits_addr; // @[SimTarget.scala 16:24:@158243.4]
  wire [31:0] Fringe_io_memStreams_stores_0_cmd_bits_size; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_memStreams_stores_0_data_ready; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_memStreams_stores_0_data_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [31:0] Fringe_io_memStreams_stores_0_data_bits_wdata_0; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_memStreams_stores_0_data_bits_wstrb; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_memStreams_stores_0_wresp_ready; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_memStreams_stores_0_wresp_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_memStreams_stores_0_wresp_bits; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_cmd_ready; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_cmd_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_dram_0_cmd_bits_addr; // @[SimTarget.scala 16:24:@158243.4]
  wire [31:0] Fringe_io_dram_0_cmd_bits_size; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_dram_0_cmd_bits_rawAddr; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_cmd_bits_isWr; // @[SimTarget.scala 16:24:@158243.4]
  wire [31:0] Fringe_io_dram_0_cmd_bits_tag; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_ready; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_0; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_1; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_2; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_3; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_4; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_5; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_6; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_7; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_8; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_9; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_10; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_11; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_12; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_13; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_14; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_15; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_16; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_17; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_18; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_19; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_20; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_21; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_22; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_23; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_24; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_25; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_26; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_27; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_28; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_29; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_30; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_31; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_32; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_33; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_34; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_35; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_36; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_37; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_38; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_39; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_40; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_41; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_42; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_43; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_44; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_45; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_46; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_47; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_48; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_49; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_50; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_51; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_52; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_53; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_54; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_55; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_56; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_57; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_58; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_59; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_60; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_61; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_62; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_wdata_bits_wdata_63; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_0; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_1; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_2; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_3; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_4; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_5; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_6; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_7; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_8; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_9; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_10; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_11; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_12; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_13; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_14; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_15; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_16; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_17; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_18; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_19; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_20; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_21; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_22; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_23; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_24; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_25; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_26; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_27; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_28; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_29; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_30; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_31; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_32; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_33; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_34; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_35; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_36; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_37; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_38; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_39; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_40; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_41; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_42; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_43; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_44; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_45; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_46; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_47; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_48; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_49; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_50; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_51; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_52; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_53; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_54; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_55; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_56; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_57; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_58; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_59; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_60; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_61; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_62; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wstrb_63; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wdata_bits_wlast; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_rresp_ready; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_rresp_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_0; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_1; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_2; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_3; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_4; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_5; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_6; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_7; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_8; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_9; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_10; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_11; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_12; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_13; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_14; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_15; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_16; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_17; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_18; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_19; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_20; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_21; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_22; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_23; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_24; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_25; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_26; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_27; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_28; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_29; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_30; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_31; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_32; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_33; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_34; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_35; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_36; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_37; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_38; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_39; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_40; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_41; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_42; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_43; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_44; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_45; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_46; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_47; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_48; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_49; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_50; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_51; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_52; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_53; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_54; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_55; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_56; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_57; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_58; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_59; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_60; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_61; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_62; // @[SimTarget.scala 16:24:@158243.4]
  wire [7:0] Fringe_io_dram_0_rresp_bits_rdata_63; // @[SimTarget.scala 16:24:@158243.4]
  wire [31:0] Fringe_io_dram_0_rresp_bits_tag; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wresp_ready; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_dram_0_wresp_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire [31:0] Fringe_io_dram_0_wresp_bits_tag; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_heap_0_req_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_heap_0_req_bits_allocDealloc; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_heap_0_req_bits_sizeAddr; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_heap_0_resp_valid; // @[SimTarget.scala 16:24:@158243.4]
  wire  Fringe_io_heap_0_resp_bits_allocDealloc; // @[SimTarget.scala 16:24:@158243.4]
  wire [63:0] Fringe_io_heap_0_resp_bits_sizeAddr; // @[SimTarget.scala 16:24:@158243.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@157688.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_cmd_bits_addr_16(accel_io_memStreams_gathers_0_cmd_bits_addr_16),
    .io_memStreams_gathers_0_cmd_bits_addr_17(accel_io_memStreams_gathers_0_cmd_bits_addr_17),
    .io_memStreams_gathers_0_cmd_bits_addr_18(accel_io_memStreams_gathers_0_cmd_bits_addr_18),
    .io_memStreams_gathers_0_cmd_bits_addr_19(accel_io_memStreams_gathers_0_cmd_bits_addr_19),
    .io_memStreams_gathers_0_cmd_bits_addr_20(accel_io_memStreams_gathers_0_cmd_bits_addr_20),
    .io_memStreams_gathers_0_cmd_bits_addr_21(accel_io_memStreams_gathers_0_cmd_bits_addr_21),
    .io_memStreams_gathers_0_cmd_bits_addr_22(accel_io_memStreams_gathers_0_cmd_bits_addr_22),
    .io_memStreams_gathers_0_cmd_bits_addr_23(accel_io_memStreams_gathers_0_cmd_bits_addr_23),
    .io_memStreams_gathers_0_cmd_bits_addr_24(accel_io_memStreams_gathers_0_cmd_bits_addr_24),
    .io_memStreams_gathers_0_cmd_bits_addr_25(accel_io_memStreams_gathers_0_cmd_bits_addr_25),
    .io_memStreams_gathers_0_cmd_bits_addr_26(accel_io_memStreams_gathers_0_cmd_bits_addr_26),
    .io_memStreams_gathers_0_cmd_bits_addr_27(accel_io_memStreams_gathers_0_cmd_bits_addr_27),
    .io_memStreams_gathers_0_cmd_bits_addr_28(accel_io_memStreams_gathers_0_cmd_bits_addr_28),
    .io_memStreams_gathers_0_cmd_bits_addr_29(accel_io_memStreams_gathers_0_cmd_bits_addr_29),
    .io_memStreams_gathers_0_cmd_bits_addr_30(accel_io_memStreams_gathers_0_cmd_bits_addr_30),
    .io_memStreams_gathers_0_cmd_bits_addr_31(accel_io_memStreams_gathers_0_cmd_bits_addr_31),
    .io_memStreams_gathers_0_cmd_bits_addr_32(accel_io_memStreams_gathers_0_cmd_bits_addr_32),
    .io_memStreams_gathers_0_cmd_bits_addr_33(accel_io_memStreams_gathers_0_cmd_bits_addr_33),
    .io_memStreams_gathers_0_cmd_bits_addr_34(accel_io_memStreams_gathers_0_cmd_bits_addr_34),
    .io_memStreams_gathers_0_cmd_bits_addr_35(accel_io_memStreams_gathers_0_cmd_bits_addr_35),
    .io_memStreams_gathers_0_cmd_bits_addr_36(accel_io_memStreams_gathers_0_cmd_bits_addr_36),
    .io_memStreams_gathers_0_cmd_bits_addr_37(accel_io_memStreams_gathers_0_cmd_bits_addr_37),
    .io_memStreams_gathers_0_cmd_bits_addr_38(accel_io_memStreams_gathers_0_cmd_bits_addr_38),
    .io_memStreams_gathers_0_cmd_bits_addr_39(accel_io_memStreams_gathers_0_cmd_bits_addr_39),
    .io_memStreams_gathers_0_cmd_bits_addr_40(accel_io_memStreams_gathers_0_cmd_bits_addr_40),
    .io_memStreams_gathers_0_cmd_bits_addr_41(accel_io_memStreams_gathers_0_cmd_bits_addr_41),
    .io_memStreams_gathers_0_cmd_bits_addr_42(accel_io_memStreams_gathers_0_cmd_bits_addr_42),
    .io_memStreams_gathers_0_cmd_bits_addr_43(accel_io_memStreams_gathers_0_cmd_bits_addr_43),
    .io_memStreams_gathers_0_cmd_bits_addr_44(accel_io_memStreams_gathers_0_cmd_bits_addr_44),
    .io_memStreams_gathers_0_cmd_bits_addr_45(accel_io_memStreams_gathers_0_cmd_bits_addr_45),
    .io_memStreams_gathers_0_cmd_bits_addr_46(accel_io_memStreams_gathers_0_cmd_bits_addr_46),
    .io_memStreams_gathers_0_cmd_bits_addr_47(accel_io_memStreams_gathers_0_cmd_bits_addr_47),
    .io_memStreams_gathers_0_cmd_bits_addr_48(accel_io_memStreams_gathers_0_cmd_bits_addr_48),
    .io_memStreams_gathers_0_cmd_bits_addr_49(accel_io_memStreams_gathers_0_cmd_bits_addr_49),
    .io_memStreams_gathers_0_cmd_bits_addr_50(accel_io_memStreams_gathers_0_cmd_bits_addr_50),
    .io_memStreams_gathers_0_cmd_bits_addr_51(accel_io_memStreams_gathers_0_cmd_bits_addr_51),
    .io_memStreams_gathers_0_cmd_bits_addr_52(accel_io_memStreams_gathers_0_cmd_bits_addr_52),
    .io_memStreams_gathers_0_cmd_bits_addr_53(accel_io_memStreams_gathers_0_cmd_bits_addr_53),
    .io_memStreams_gathers_0_cmd_bits_addr_54(accel_io_memStreams_gathers_0_cmd_bits_addr_54),
    .io_memStreams_gathers_0_cmd_bits_addr_55(accel_io_memStreams_gathers_0_cmd_bits_addr_55),
    .io_memStreams_gathers_0_cmd_bits_addr_56(accel_io_memStreams_gathers_0_cmd_bits_addr_56),
    .io_memStreams_gathers_0_cmd_bits_addr_57(accel_io_memStreams_gathers_0_cmd_bits_addr_57),
    .io_memStreams_gathers_0_cmd_bits_addr_58(accel_io_memStreams_gathers_0_cmd_bits_addr_58),
    .io_memStreams_gathers_0_cmd_bits_addr_59(accel_io_memStreams_gathers_0_cmd_bits_addr_59),
    .io_memStreams_gathers_0_cmd_bits_addr_60(accel_io_memStreams_gathers_0_cmd_bits_addr_60),
    .io_memStreams_gathers_0_cmd_bits_addr_61(accel_io_memStreams_gathers_0_cmd_bits_addr_61),
    .io_memStreams_gathers_0_cmd_bits_addr_62(accel_io_memStreams_gathers_0_cmd_bits_addr_62),
    .io_memStreams_gathers_0_cmd_bits_addr_63(accel_io_memStreams_gathers_0_cmd_bits_addr_63),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_gathers_0_data_bits_16(accel_io_memStreams_gathers_0_data_bits_16),
    .io_memStreams_gathers_0_data_bits_17(accel_io_memStreams_gathers_0_data_bits_17),
    .io_memStreams_gathers_0_data_bits_18(accel_io_memStreams_gathers_0_data_bits_18),
    .io_memStreams_gathers_0_data_bits_19(accel_io_memStreams_gathers_0_data_bits_19),
    .io_memStreams_gathers_0_data_bits_20(accel_io_memStreams_gathers_0_data_bits_20),
    .io_memStreams_gathers_0_data_bits_21(accel_io_memStreams_gathers_0_data_bits_21),
    .io_memStreams_gathers_0_data_bits_22(accel_io_memStreams_gathers_0_data_bits_22),
    .io_memStreams_gathers_0_data_bits_23(accel_io_memStreams_gathers_0_data_bits_23),
    .io_memStreams_gathers_0_data_bits_24(accel_io_memStreams_gathers_0_data_bits_24),
    .io_memStreams_gathers_0_data_bits_25(accel_io_memStreams_gathers_0_data_bits_25),
    .io_memStreams_gathers_0_data_bits_26(accel_io_memStreams_gathers_0_data_bits_26),
    .io_memStreams_gathers_0_data_bits_27(accel_io_memStreams_gathers_0_data_bits_27),
    .io_memStreams_gathers_0_data_bits_28(accel_io_memStreams_gathers_0_data_bits_28),
    .io_memStreams_gathers_0_data_bits_29(accel_io_memStreams_gathers_0_data_bits_29),
    .io_memStreams_gathers_0_data_bits_30(accel_io_memStreams_gathers_0_data_bits_30),
    .io_memStreams_gathers_0_data_bits_31(accel_io_memStreams_gathers_0_data_bits_31),
    .io_memStreams_gathers_0_data_bits_32(accel_io_memStreams_gathers_0_data_bits_32),
    .io_memStreams_gathers_0_data_bits_33(accel_io_memStreams_gathers_0_data_bits_33),
    .io_memStreams_gathers_0_data_bits_34(accel_io_memStreams_gathers_0_data_bits_34),
    .io_memStreams_gathers_0_data_bits_35(accel_io_memStreams_gathers_0_data_bits_35),
    .io_memStreams_gathers_0_data_bits_36(accel_io_memStreams_gathers_0_data_bits_36),
    .io_memStreams_gathers_0_data_bits_37(accel_io_memStreams_gathers_0_data_bits_37),
    .io_memStreams_gathers_0_data_bits_38(accel_io_memStreams_gathers_0_data_bits_38),
    .io_memStreams_gathers_0_data_bits_39(accel_io_memStreams_gathers_0_data_bits_39),
    .io_memStreams_gathers_0_data_bits_40(accel_io_memStreams_gathers_0_data_bits_40),
    .io_memStreams_gathers_0_data_bits_41(accel_io_memStreams_gathers_0_data_bits_41),
    .io_memStreams_gathers_0_data_bits_42(accel_io_memStreams_gathers_0_data_bits_42),
    .io_memStreams_gathers_0_data_bits_43(accel_io_memStreams_gathers_0_data_bits_43),
    .io_memStreams_gathers_0_data_bits_44(accel_io_memStreams_gathers_0_data_bits_44),
    .io_memStreams_gathers_0_data_bits_45(accel_io_memStreams_gathers_0_data_bits_45),
    .io_memStreams_gathers_0_data_bits_46(accel_io_memStreams_gathers_0_data_bits_46),
    .io_memStreams_gathers_0_data_bits_47(accel_io_memStreams_gathers_0_data_bits_47),
    .io_memStreams_gathers_0_data_bits_48(accel_io_memStreams_gathers_0_data_bits_48),
    .io_memStreams_gathers_0_data_bits_49(accel_io_memStreams_gathers_0_data_bits_49),
    .io_memStreams_gathers_0_data_bits_50(accel_io_memStreams_gathers_0_data_bits_50),
    .io_memStreams_gathers_0_data_bits_51(accel_io_memStreams_gathers_0_data_bits_51),
    .io_memStreams_gathers_0_data_bits_52(accel_io_memStreams_gathers_0_data_bits_52),
    .io_memStreams_gathers_0_data_bits_53(accel_io_memStreams_gathers_0_data_bits_53),
    .io_memStreams_gathers_0_data_bits_54(accel_io_memStreams_gathers_0_data_bits_54),
    .io_memStreams_gathers_0_data_bits_55(accel_io_memStreams_gathers_0_data_bits_55),
    .io_memStreams_gathers_0_data_bits_56(accel_io_memStreams_gathers_0_data_bits_56),
    .io_memStreams_gathers_0_data_bits_57(accel_io_memStreams_gathers_0_data_bits_57),
    .io_memStreams_gathers_0_data_bits_58(accel_io_memStreams_gathers_0_data_bits_58),
    .io_memStreams_gathers_0_data_bits_59(accel_io_memStreams_gathers_0_data_bits_59),
    .io_memStreams_gathers_0_data_bits_60(accel_io_memStreams_gathers_0_data_bits_60),
    .io_memStreams_gathers_0_data_bits_61(accel_io_memStreams_gathers_0_data_bits_61),
    .io_memStreams_gathers_0_data_bits_62(accel_io_memStreams_gathers_0_data_bits_62),
    .io_memStreams_gathers_0_data_bits_63(accel_io_memStreams_gathers_0_data_bits_63),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_16(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_16),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_17(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_17),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_18(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_18),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_19(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_19),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_20(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_20),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_21(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_21),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_22(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_22),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_23(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_23),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_24(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_24),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_25(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_25),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_26(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_26),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_27(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_27),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_28(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_28),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_29(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_29),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_30(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_30),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_31(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_31),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_32(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_32),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_33(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_33),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_34(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_34),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_35(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_35),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_36(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_36),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_37(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_37),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_38(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_38),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_39(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_39),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_40(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_40),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_41(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_41),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_42(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_42),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_43(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_43),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_44(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_44),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_45(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_45),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_46(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_46),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_47(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_47),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_48(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_48),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_49(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_49),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_50(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_50),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_51(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_51),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_52(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_52),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_53(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_53),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_54(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_54),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_55(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_55),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_56(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_56),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_57(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_57),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_58(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_58),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_59(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_59),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_60(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_60),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_61(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_61),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_62(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_62),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_63(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_63),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_16(accel_io_memStreams_scatters_0_cmd_bits_wdata_16),
    .io_memStreams_scatters_0_cmd_bits_wdata_17(accel_io_memStreams_scatters_0_cmd_bits_wdata_17),
    .io_memStreams_scatters_0_cmd_bits_wdata_18(accel_io_memStreams_scatters_0_cmd_bits_wdata_18),
    .io_memStreams_scatters_0_cmd_bits_wdata_19(accel_io_memStreams_scatters_0_cmd_bits_wdata_19),
    .io_memStreams_scatters_0_cmd_bits_wdata_20(accel_io_memStreams_scatters_0_cmd_bits_wdata_20),
    .io_memStreams_scatters_0_cmd_bits_wdata_21(accel_io_memStreams_scatters_0_cmd_bits_wdata_21),
    .io_memStreams_scatters_0_cmd_bits_wdata_22(accel_io_memStreams_scatters_0_cmd_bits_wdata_22),
    .io_memStreams_scatters_0_cmd_bits_wdata_23(accel_io_memStreams_scatters_0_cmd_bits_wdata_23),
    .io_memStreams_scatters_0_cmd_bits_wdata_24(accel_io_memStreams_scatters_0_cmd_bits_wdata_24),
    .io_memStreams_scatters_0_cmd_bits_wdata_25(accel_io_memStreams_scatters_0_cmd_bits_wdata_25),
    .io_memStreams_scatters_0_cmd_bits_wdata_26(accel_io_memStreams_scatters_0_cmd_bits_wdata_26),
    .io_memStreams_scatters_0_cmd_bits_wdata_27(accel_io_memStreams_scatters_0_cmd_bits_wdata_27),
    .io_memStreams_scatters_0_cmd_bits_wdata_28(accel_io_memStreams_scatters_0_cmd_bits_wdata_28),
    .io_memStreams_scatters_0_cmd_bits_wdata_29(accel_io_memStreams_scatters_0_cmd_bits_wdata_29),
    .io_memStreams_scatters_0_cmd_bits_wdata_30(accel_io_memStreams_scatters_0_cmd_bits_wdata_30),
    .io_memStreams_scatters_0_cmd_bits_wdata_31(accel_io_memStreams_scatters_0_cmd_bits_wdata_31),
    .io_memStreams_scatters_0_cmd_bits_wdata_32(accel_io_memStreams_scatters_0_cmd_bits_wdata_32),
    .io_memStreams_scatters_0_cmd_bits_wdata_33(accel_io_memStreams_scatters_0_cmd_bits_wdata_33),
    .io_memStreams_scatters_0_cmd_bits_wdata_34(accel_io_memStreams_scatters_0_cmd_bits_wdata_34),
    .io_memStreams_scatters_0_cmd_bits_wdata_35(accel_io_memStreams_scatters_0_cmd_bits_wdata_35),
    .io_memStreams_scatters_0_cmd_bits_wdata_36(accel_io_memStreams_scatters_0_cmd_bits_wdata_36),
    .io_memStreams_scatters_0_cmd_bits_wdata_37(accel_io_memStreams_scatters_0_cmd_bits_wdata_37),
    .io_memStreams_scatters_0_cmd_bits_wdata_38(accel_io_memStreams_scatters_0_cmd_bits_wdata_38),
    .io_memStreams_scatters_0_cmd_bits_wdata_39(accel_io_memStreams_scatters_0_cmd_bits_wdata_39),
    .io_memStreams_scatters_0_cmd_bits_wdata_40(accel_io_memStreams_scatters_0_cmd_bits_wdata_40),
    .io_memStreams_scatters_0_cmd_bits_wdata_41(accel_io_memStreams_scatters_0_cmd_bits_wdata_41),
    .io_memStreams_scatters_0_cmd_bits_wdata_42(accel_io_memStreams_scatters_0_cmd_bits_wdata_42),
    .io_memStreams_scatters_0_cmd_bits_wdata_43(accel_io_memStreams_scatters_0_cmd_bits_wdata_43),
    .io_memStreams_scatters_0_cmd_bits_wdata_44(accel_io_memStreams_scatters_0_cmd_bits_wdata_44),
    .io_memStreams_scatters_0_cmd_bits_wdata_45(accel_io_memStreams_scatters_0_cmd_bits_wdata_45),
    .io_memStreams_scatters_0_cmd_bits_wdata_46(accel_io_memStreams_scatters_0_cmd_bits_wdata_46),
    .io_memStreams_scatters_0_cmd_bits_wdata_47(accel_io_memStreams_scatters_0_cmd_bits_wdata_47),
    .io_memStreams_scatters_0_cmd_bits_wdata_48(accel_io_memStreams_scatters_0_cmd_bits_wdata_48),
    .io_memStreams_scatters_0_cmd_bits_wdata_49(accel_io_memStreams_scatters_0_cmd_bits_wdata_49),
    .io_memStreams_scatters_0_cmd_bits_wdata_50(accel_io_memStreams_scatters_0_cmd_bits_wdata_50),
    .io_memStreams_scatters_0_cmd_bits_wdata_51(accel_io_memStreams_scatters_0_cmd_bits_wdata_51),
    .io_memStreams_scatters_0_cmd_bits_wdata_52(accel_io_memStreams_scatters_0_cmd_bits_wdata_52),
    .io_memStreams_scatters_0_cmd_bits_wdata_53(accel_io_memStreams_scatters_0_cmd_bits_wdata_53),
    .io_memStreams_scatters_0_cmd_bits_wdata_54(accel_io_memStreams_scatters_0_cmd_bits_wdata_54),
    .io_memStreams_scatters_0_cmd_bits_wdata_55(accel_io_memStreams_scatters_0_cmd_bits_wdata_55),
    .io_memStreams_scatters_0_cmd_bits_wdata_56(accel_io_memStreams_scatters_0_cmd_bits_wdata_56),
    .io_memStreams_scatters_0_cmd_bits_wdata_57(accel_io_memStreams_scatters_0_cmd_bits_wdata_57),
    .io_memStreams_scatters_0_cmd_bits_wdata_58(accel_io_memStreams_scatters_0_cmd_bits_wdata_58),
    .io_memStreams_scatters_0_cmd_bits_wdata_59(accel_io_memStreams_scatters_0_cmd_bits_wdata_59),
    .io_memStreams_scatters_0_cmd_bits_wdata_60(accel_io_memStreams_scatters_0_cmd_bits_wdata_60),
    .io_memStreams_scatters_0_cmd_bits_wdata_61(accel_io_memStreams_scatters_0_cmd_bits_wdata_61),
    .io_memStreams_scatters_0_cmd_bits_wdata_62(accel_io_memStreams_scatters_0_cmd_bits_wdata_62),
    .io_memStreams_scatters_0_cmd_bits_wdata_63(accel_io_memStreams_scatters_0_cmd_bits_wdata_63),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo),
    .io_argOuts_1_port_ready(accel_io_argOuts_1_port_ready),
    .io_argOuts_1_port_valid(accel_io_argOuts_1_port_valid),
    .io_argOuts_1_port_bits(accel_io_argOuts_1_port_bits),
    .io_argOuts_1_echo(accel_io_argOuts_1_echo),
    .io_argOuts_2_port_ready(accel_io_argOuts_2_port_ready),
    .io_argOuts_2_port_valid(accel_io_argOuts_2_port_valid),
    .io_argOuts_2_port_bits(accel_io_argOuts_2_port_bits),
    .io_argOuts_2_echo(accel_io_argOuts_2_echo),
    .io_argOuts_3_port_ready(accel_io_argOuts_3_port_ready),
    .io_argOuts_3_port_valid(accel_io_argOuts_3_port_valid),
    .io_argOuts_3_port_bits(accel_io_argOuts_3_port_bits),
    .io_argOuts_3_echo(accel_io_argOuts_3_echo),
    .io_argOuts_4_port_ready(accel_io_argOuts_4_port_ready),
    .io_argOuts_4_port_valid(accel_io_argOuts_4_port_valid),
    .io_argOuts_4_port_bits(accel_io_argOuts_4_port_bits),
    .io_argOuts_4_echo(accel_io_argOuts_4_echo),
    .io_argOuts_5_port_ready(accel_io_argOuts_5_port_ready),
    .io_argOuts_5_port_valid(accel_io_argOuts_5_port_valid),
    .io_argOuts_5_port_bits(accel_io_argOuts_5_port_bits),
    .io_argOuts_5_echo(accel_io_argOuts_5_echo),
    .io_argOuts_6_port_ready(accel_io_argOuts_6_port_ready),
    .io_argOuts_6_port_valid(accel_io_argOuts_6_port_valid),
    .io_argOuts_6_port_bits(accel_io_argOuts_6_port_bits),
    .io_argOuts_6_echo(accel_io_argOuts_6_echo),
    .io_argOuts_7_port_ready(accel_io_argOuts_7_port_ready),
    .io_argOuts_7_port_valid(accel_io_argOuts_7_port_valid),
    .io_argOuts_7_port_bits(accel_io_argOuts_7_port_bits),
    .io_argOuts_7_echo(accel_io_argOuts_7_echo),
    .io_argOuts_8_port_ready(accel_io_argOuts_8_port_ready),
    .io_argOuts_8_port_valid(accel_io_argOuts_8_port_valid),
    .io_argOuts_8_port_bits(accel_io_argOuts_8_port_bits),
    .io_argOuts_8_echo(accel_io_argOuts_8_echo),
    .io_argOuts_9_port_ready(accel_io_argOuts_9_port_ready),
    .io_argOuts_9_port_valid(accel_io_argOuts_9_port_valid),
    .io_argOuts_9_port_bits(accel_io_argOuts_9_port_bits),
    .io_argOuts_9_echo(accel_io_argOuts_9_echo),
    .io_argOuts_10_port_ready(accel_io_argOuts_10_port_ready),
    .io_argOuts_10_port_valid(accel_io_argOuts_10_port_valid),
    .io_argOuts_10_port_bits(accel_io_argOuts_10_port_bits),
    .io_argOuts_10_echo(accel_io_argOuts_10_echo),
    .io_argOuts_11_port_ready(accel_io_argOuts_11_port_ready),
    .io_argOuts_11_port_valid(accel_io_argOuts_11_port_valid),
    .io_argOuts_11_port_bits(accel_io_argOuts_11_port_bits),
    .io_argOuts_11_echo(accel_io_argOuts_11_echo),
    .io_argOuts_12_port_ready(accel_io_argOuts_12_port_ready),
    .io_argOuts_12_port_valid(accel_io_argOuts_12_port_valid),
    .io_argOuts_12_port_bits(accel_io_argOuts_12_port_bits),
    .io_argOuts_12_echo(accel_io_argOuts_12_echo),
    .io_argOuts_13_port_ready(accel_io_argOuts_13_port_ready),
    .io_argOuts_13_port_valid(accel_io_argOuts_13_port_valid),
    .io_argOuts_13_port_bits(accel_io_argOuts_13_port_bits),
    .io_argOuts_13_echo(accel_io_argOuts_13_echo),
    .io_argOuts_14_port_ready(accel_io_argOuts_14_port_ready),
    .io_argOuts_14_port_valid(accel_io_argOuts_14_port_valid),
    .io_argOuts_14_port_bits(accel_io_argOuts_14_port_bits),
    .io_argOuts_14_echo(accel_io_argOuts_14_echo),
    .io_argOuts_15_port_ready(accel_io_argOuts_15_port_ready),
    .io_argOuts_15_port_valid(accel_io_argOuts_15_port_valid),
    .io_argOuts_15_port_bits(accel_io_argOuts_15_port_bits),
    .io_argOuts_15_echo(accel_io_argOuts_15_echo),
    .io_argOuts_16_port_ready(accel_io_argOuts_16_port_ready),
    .io_argOuts_16_port_valid(accel_io_argOuts_16_port_valid),
    .io_argOuts_16_port_bits(accel_io_argOuts_16_port_bits),
    .io_argOuts_16_echo(accel_io_argOuts_16_echo),
    .io_argOuts_17_port_ready(accel_io_argOuts_17_port_ready),
    .io_argOuts_17_port_valid(accel_io_argOuts_17_port_valid),
    .io_argOuts_17_port_bits(accel_io_argOuts_17_port_bits),
    .io_argOuts_17_echo(accel_io_argOuts_17_echo),
    .io_argOuts_18_port_ready(accel_io_argOuts_18_port_ready),
    .io_argOuts_18_port_valid(accel_io_argOuts_18_port_valid),
    .io_argOuts_18_port_bits(accel_io_argOuts_18_port_bits),
    .io_argOuts_18_echo(accel_io_argOuts_18_echo),
    .io_argOuts_19_port_ready(accel_io_argOuts_19_port_ready),
    .io_argOuts_19_port_valid(accel_io_argOuts_19_port_valid),
    .io_argOuts_19_port_bits(accel_io_argOuts_19_port_bits),
    .io_argOuts_19_echo(accel_io_argOuts_19_echo),
    .io_argOuts_20_port_ready(accel_io_argOuts_20_port_ready),
    .io_argOuts_20_port_valid(accel_io_argOuts_20_port_valid),
    .io_argOuts_20_port_bits(accel_io_argOuts_20_port_bits),
    .io_argOuts_20_echo(accel_io_argOuts_20_echo),
    .io_argOuts_21_port_ready(accel_io_argOuts_21_port_ready),
    .io_argOuts_21_port_valid(accel_io_argOuts_21_port_valid),
    .io_argOuts_21_port_bits(accel_io_argOuts_21_port_bits),
    .io_argOuts_21_echo(accel_io_argOuts_21_echo),
    .io_argOuts_22_port_ready(accel_io_argOuts_22_port_ready),
    .io_argOuts_22_port_valid(accel_io_argOuts_22_port_valid),
    .io_argOuts_22_port_bits(accel_io_argOuts_22_port_bits),
    .io_argOuts_22_echo(accel_io_argOuts_22_echo),
    .io_argOuts_23_port_ready(accel_io_argOuts_23_port_ready),
    .io_argOuts_23_port_valid(accel_io_argOuts_23_port_valid),
    .io_argOuts_23_port_bits(accel_io_argOuts_23_port_bits),
    .io_argOuts_23_echo(accel_io_argOuts_23_echo),
    .io_argOuts_24_port_ready(accel_io_argOuts_24_port_ready),
    .io_argOuts_24_port_valid(accel_io_argOuts_24_port_valid),
    .io_argOuts_24_port_bits(accel_io_argOuts_24_port_bits),
    .io_argOuts_24_echo(accel_io_argOuts_24_echo),
    .io_argOuts_25_port_ready(accel_io_argOuts_25_port_ready),
    .io_argOuts_25_port_valid(accel_io_argOuts_25_port_valid),
    .io_argOuts_25_port_bits(accel_io_argOuts_25_port_bits),
    .io_argOuts_25_echo(accel_io_argOuts_25_echo),
    .io_argOuts_26_port_ready(accel_io_argOuts_26_port_ready),
    .io_argOuts_26_port_valid(accel_io_argOuts_26_port_valid),
    .io_argOuts_26_port_bits(accel_io_argOuts_26_port_bits),
    .io_argOuts_26_echo(accel_io_argOuts_26_echo),
    .io_argOuts_27_port_ready(accel_io_argOuts_27_port_ready),
    .io_argOuts_27_port_valid(accel_io_argOuts_27_port_valid),
    .io_argOuts_27_port_bits(accel_io_argOuts_27_port_bits),
    .io_argOuts_27_echo(accel_io_argOuts_27_echo),
    .io_argOuts_28_port_ready(accel_io_argOuts_28_port_ready),
    .io_argOuts_28_port_valid(accel_io_argOuts_28_port_valid),
    .io_argOuts_28_port_bits(accel_io_argOuts_28_port_bits),
    .io_argOuts_28_echo(accel_io_argOuts_28_echo),
    .io_argOuts_29_port_ready(accel_io_argOuts_29_port_ready),
    .io_argOuts_29_port_valid(accel_io_argOuts_29_port_valid),
    .io_argOuts_29_port_bits(accel_io_argOuts_29_port_bits),
    .io_argOuts_29_echo(accel_io_argOuts_29_echo),
    .io_argOuts_30_port_ready(accel_io_argOuts_30_port_ready),
    .io_argOuts_30_port_valid(accel_io_argOuts_30_port_valid),
    .io_argOuts_30_port_bits(accel_io_argOuts_30_port_bits),
    .io_argOuts_30_echo(accel_io_argOuts_30_echo),
    .io_argOuts_31_port_ready(accel_io_argOuts_31_port_ready),
    .io_argOuts_31_port_valid(accel_io_argOuts_31_port_valid),
    .io_argOuts_31_port_bits(accel_io_argOuts_31_port_bits),
    .io_argOuts_31_echo(accel_io_argOuts_31_echo),
    .io_argOuts_32_port_ready(accel_io_argOuts_32_port_ready),
    .io_argOuts_32_port_valid(accel_io_argOuts_32_port_valid),
    .io_argOuts_32_port_bits(accel_io_argOuts_32_port_bits),
    .io_argOuts_32_echo(accel_io_argOuts_32_echo),
    .io_argOuts_33_port_ready(accel_io_argOuts_33_port_ready),
    .io_argOuts_33_port_valid(accel_io_argOuts_33_port_valid),
    .io_argOuts_33_port_bits(accel_io_argOuts_33_port_bits),
    .io_argOuts_33_echo(accel_io_argOuts_33_echo),
    .io_argOuts_34_port_ready(accel_io_argOuts_34_port_ready),
    .io_argOuts_34_port_valid(accel_io_argOuts_34_port_valid),
    .io_argOuts_34_port_bits(accel_io_argOuts_34_port_bits),
    .io_argOuts_34_echo(accel_io_argOuts_34_echo),
    .io_argOuts_35_port_ready(accel_io_argOuts_35_port_ready),
    .io_argOuts_35_port_valid(accel_io_argOuts_35_port_valid),
    .io_argOuts_35_port_bits(accel_io_argOuts_35_port_bits),
    .io_argOuts_35_echo(accel_io_argOuts_35_echo),
    .io_argOuts_36_port_ready(accel_io_argOuts_36_port_ready),
    .io_argOuts_36_port_valid(accel_io_argOuts_36_port_valid),
    .io_argOuts_36_port_bits(accel_io_argOuts_36_port_bits),
    .io_argOuts_36_echo(accel_io_argOuts_36_echo),
    .io_argOuts_37_port_ready(accel_io_argOuts_37_port_ready),
    .io_argOuts_37_port_valid(accel_io_argOuts_37_port_valid),
    .io_argOuts_37_port_bits(accel_io_argOuts_37_port_bits),
    .io_argOuts_37_echo(accel_io_argOuts_37_echo),
    .io_argOuts_38_port_ready(accel_io_argOuts_38_port_ready),
    .io_argOuts_38_port_valid(accel_io_argOuts_38_port_valid),
    .io_argOuts_38_port_bits(accel_io_argOuts_38_port_bits),
    .io_argOuts_38_echo(accel_io_argOuts_38_echo),
    .io_argOuts_39_port_ready(accel_io_argOuts_39_port_ready),
    .io_argOuts_39_port_valid(accel_io_argOuts_39_port_valid),
    .io_argOuts_39_port_bits(accel_io_argOuts_39_port_bits),
    .io_argOuts_39_echo(accel_io_argOuts_39_echo),
    .io_argOuts_40_port_ready(accel_io_argOuts_40_port_ready),
    .io_argOuts_40_port_valid(accel_io_argOuts_40_port_valid),
    .io_argOuts_40_port_bits(accel_io_argOuts_40_port_bits),
    .io_argOuts_40_echo(accel_io_argOuts_40_echo),
    .io_argOuts_41_port_ready(accel_io_argOuts_41_port_ready),
    .io_argOuts_41_port_valid(accel_io_argOuts_41_port_valid),
    .io_argOuts_41_port_bits(accel_io_argOuts_41_port_bits),
    .io_argOuts_41_echo(accel_io_argOuts_41_echo),
    .io_argOuts_42_port_ready(accel_io_argOuts_42_port_ready),
    .io_argOuts_42_port_valid(accel_io_argOuts_42_port_valid),
    .io_argOuts_42_port_bits(accel_io_argOuts_42_port_bits),
    .io_argOuts_42_echo(accel_io_argOuts_42_echo),
    .io_argOuts_43_port_ready(accel_io_argOuts_43_port_ready),
    .io_argOuts_43_port_valid(accel_io_argOuts_43_port_valid),
    .io_argOuts_43_port_bits(accel_io_argOuts_43_port_bits),
    .io_argOuts_43_echo(accel_io_argOuts_43_echo),
    .io_argOuts_44_port_ready(accel_io_argOuts_44_port_ready),
    .io_argOuts_44_port_valid(accel_io_argOuts_44_port_valid),
    .io_argOuts_44_port_bits(accel_io_argOuts_44_port_bits),
    .io_argOuts_44_echo(accel_io_argOuts_44_echo),
    .io_argOuts_45_port_ready(accel_io_argOuts_45_port_ready),
    .io_argOuts_45_port_valid(accel_io_argOuts_45_port_valid),
    .io_argOuts_45_port_bits(accel_io_argOuts_45_port_bits),
    .io_argOuts_45_echo(accel_io_argOuts_45_echo),
    .io_argOuts_46_port_ready(accel_io_argOuts_46_port_ready),
    .io_argOuts_46_port_valid(accel_io_argOuts_46_port_valid),
    .io_argOuts_46_port_bits(accel_io_argOuts_46_port_bits),
    .io_argOuts_46_echo(accel_io_argOuts_46_echo),
    .io_argOuts_47_port_ready(accel_io_argOuts_47_port_ready),
    .io_argOuts_47_port_valid(accel_io_argOuts_47_port_valid),
    .io_argOuts_47_port_bits(accel_io_argOuts_47_port_bits),
    .io_argOuts_47_echo(accel_io_argOuts_47_echo),
    .io_argOuts_48_port_ready(accel_io_argOuts_48_port_ready),
    .io_argOuts_48_port_valid(accel_io_argOuts_48_port_valid),
    .io_argOuts_48_port_bits(accel_io_argOuts_48_port_bits),
    .io_argOuts_48_echo(accel_io_argOuts_48_echo),
    .io_argOuts_49_port_ready(accel_io_argOuts_49_port_ready),
    .io_argOuts_49_port_valid(accel_io_argOuts_49_port_valid),
    .io_argOuts_49_port_bits(accel_io_argOuts_49_port_bits),
    .io_argOuts_49_echo(accel_io_argOuts_49_echo),
    .io_argOuts_50_port_ready(accel_io_argOuts_50_port_ready),
    .io_argOuts_50_port_valid(accel_io_argOuts_50_port_valid),
    .io_argOuts_50_port_bits(accel_io_argOuts_50_port_bits),
    .io_argOuts_50_echo(accel_io_argOuts_50_echo),
    .io_argOuts_51_port_ready(accel_io_argOuts_51_port_ready),
    .io_argOuts_51_port_valid(accel_io_argOuts_51_port_valid),
    .io_argOuts_51_port_bits(accel_io_argOuts_51_port_bits),
    .io_argOuts_51_echo(accel_io_argOuts_51_echo),
    .io_argOuts_52_port_ready(accel_io_argOuts_52_port_ready),
    .io_argOuts_52_port_valid(accel_io_argOuts_52_port_valid),
    .io_argOuts_52_port_bits(accel_io_argOuts_52_port_bits),
    .io_argOuts_52_echo(accel_io_argOuts_52_echo),
    .io_argOuts_53_port_ready(accel_io_argOuts_53_port_ready),
    .io_argOuts_53_port_valid(accel_io_argOuts_53_port_valid),
    .io_argOuts_53_port_bits(accel_io_argOuts_53_port_bits),
    .io_argOuts_53_echo(accel_io_argOuts_53_echo),
    .io_argOuts_54_port_ready(accel_io_argOuts_54_port_ready),
    .io_argOuts_54_port_valid(accel_io_argOuts_54_port_valid),
    .io_argOuts_54_port_bits(accel_io_argOuts_54_port_bits),
    .io_argOuts_54_echo(accel_io_argOuts_54_echo),
    .io_argOuts_55_port_ready(accel_io_argOuts_55_port_ready),
    .io_argOuts_55_port_valid(accel_io_argOuts_55_port_valid),
    .io_argOuts_55_port_bits(accel_io_argOuts_55_port_bits),
    .io_argOuts_55_echo(accel_io_argOuts_55_echo),
    .io_argOuts_56_port_ready(accel_io_argOuts_56_port_ready),
    .io_argOuts_56_port_valid(accel_io_argOuts_56_port_valid),
    .io_argOuts_56_port_bits(accel_io_argOuts_56_port_bits),
    .io_argOuts_56_echo(accel_io_argOuts_56_echo),
    .io_argOuts_57_port_ready(accel_io_argOuts_57_port_ready),
    .io_argOuts_57_port_valid(accel_io_argOuts_57_port_valid),
    .io_argOuts_57_port_bits(accel_io_argOuts_57_port_bits),
    .io_argOuts_57_echo(accel_io_argOuts_57_echo),
    .io_argOuts_58_port_ready(accel_io_argOuts_58_port_ready),
    .io_argOuts_58_port_valid(accel_io_argOuts_58_port_valid),
    .io_argOuts_58_port_bits(accel_io_argOuts_58_port_bits),
    .io_argOuts_58_echo(accel_io_argOuts_58_echo),
    .io_argOuts_59_port_ready(accel_io_argOuts_59_port_ready),
    .io_argOuts_59_port_valid(accel_io_argOuts_59_port_valid),
    .io_argOuts_59_port_bits(accel_io_argOuts_59_port_bits),
    .io_argOuts_59_echo(accel_io_argOuts_59_echo)
  );
  Fringe Fringe ( // @[SimTarget.scala 16:24:@158243.4]
    .clock(Fringe_clock),
    .reset(Fringe_reset),
    .io_raddr(Fringe_io_raddr),
    .io_wen(Fringe_io_wen),
    .io_waddr(Fringe_io_waddr),
    .io_wdata(Fringe_io_wdata),
    .io_rdata(Fringe_io_rdata),
    .io_enable(Fringe_io_enable),
    .io_done(Fringe_io_done),
    .io_reset(Fringe_io_reset),
    .io_argIns_0(Fringe_io_argIns_0),
    .io_argIns_1(Fringe_io_argIns_1),
    .io_argOuts_0_valid(Fringe_io_argOuts_0_valid),
    .io_argOuts_0_bits(Fringe_io_argOuts_0_bits),
    .io_argOuts_1_valid(Fringe_io_argOuts_1_valid),
    .io_argOuts_1_bits(Fringe_io_argOuts_1_bits),
    .io_argOuts_2_valid(Fringe_io_argOuts_2_valid),
    .io_argOuts_2_bits(Fringe_io_argOuts_2_bits),
    .io_argOuts_3_valid(Fringe_io_argOuts_3_valid),
    .io_argOuts_3_bits(Fringe_io_argOuts_3_bits),
    .io_argOuts_4_valid(Fringe_io_argOuts_4_valid),
    .io_argOuts_4_bits(Fringe_io_argOuts_4_bits),
    .io_argOuts_5_valid(Fringe_io_argOuts_5_valid),
    .io_argOuts_5_bits(Fringe_io_argOuts_5_bits),
    .io_argOuts_6_valid(Fringe_io_argOuts_6_valid),
    .io_argOuts_6_bits(Fringe_io_argOuts_6_bits),
    .io_argOuts_7_valid(Fringe_io_argOuts_7_valid),
    .io_argOuts_7_bits(Fringe_io_argOuts_7_bits),
    .io_argOuts_8_valid(Fringe_io_argOuts_8_valid),
    .io_argOuts_8_bits(Fringe_io_argOuts_8_bits),
    .io_argOuts_9_valid(Fringe_io_argOuts_9_valid),
    .io_argOuts_9_bits(Fringe_io_argOuts_9_bits),
    .io_argOuts_10_valid(Fringe_io_argOuts_10_valid),
    .io_argOuts_10_bits(Fringe_io_argOuts_10_bits),
    .io_argOuts_11_valid(Fringe_io_argOuts_11_valid),
    .io_argOuts_11_bits(Fringe_io_argOuts_11_bits),
    .io_argOuts_12_valid(Fringe_io_argOuts_12_valid),
    .io_argOuts_12_bits(Fringe_io_argOuts_12_bits),
    .io_argOuts_13_valid(Fringe_io_argOuts_13_valid),
    .io_argOuts_13_bits(Fringe_io_argOuts_13_bits),
    .io_argOuts_14_valid(Fringe_io_argOuts_14_valid),
    .io_argOuts_14_bits(Fringe_io_argOuts_14_bits),
    .io_argOuts_15_valid(Fringe_io_argOuts_15_valid),
    .io_argOuts_15_bits(Fringe_io_argOuts_15_bits),
    .io_argOuts_16_valid(Fringe_io_argOuts_16_valid),
    .io_argOuts_16_bits(Fringe_io_argOuts_16_bits),
    .io_argOuts_17_valid(Fringe_io_argOuts_17_valid),
    .io_argOuts_17_bits(Fringe_io_argOuts_17_bits),
    .io_argOuts_18_valid(Fringe_io_argOuts_18_valid),
    .io_argOuts_18_bits(Fringe_io_argOuts_18_bits),
    .io_argOuts_19_valid(Fringe_io_argOuts_19_valid),
    .io_argOuts_19_bits(Fringe_io_argOuts_19_bits),
    .io_argOuts_20_valid(Fringe_io_argOuts_20_valid),
    .io_argOuts_20_bits(Fringe_io_argOuts_20_bits),
    .io_argOuts_21_valid(Fringe_io_argOuts_21_valid),
    .io_argOuts_21_bits(Fringe_io_argOuts_21_bits),
    .io_argOuts_22_valid(Fringe_io_argOuts_22_valid),
    .io_argOuts_22_bits(Fringe_io_argOuts_22_bits),
    .io_argOuts_23_valid(Fringe_io_argOuts_23_valid),
    .io_argOuts_23_bits(Fringe_io_argOuts_23_bits),
    .io_argOuts_24_valid(Fringe_io_argOuts_24_valid),
    .io_argOuts_24_bits(Fringe_io_argOuts_24_bits),
    .io_argOuts_25_valid(Fringe_io_argOuts_25_valid),
    .io_argOuts_25_bits(Fringe_io_argOuts_25_bits),
    .io_argOuts_26_valid(Fringe_io_argOuts_26_valid),
    .io_argOuts_26_bits(Fringe_io_argOuts_26_bits),
    .io_argOuts_27_valid(Fringe_io_argOuts_27_valid),
    .io_argOuts_27_bits(Fringe_io_argOuts_27_bits),
    .io_argOuts_28_valid(Fringe_io_argOuts_28_valid),
    .io_argOuts_28_bits(Fringe_io_argOuts_28_bits),
    .io_argOuts_29_valid(Fringe_io_argOuts_29_valid),
    .io_argOuts_29_bits(Fringe_io_argOuts_29_bits),
    .io_argOuts_30_valid(Fringe_io_argOuts_30_valid),
    .io_argOuts_30_bits(Fringe_io_argOuts_30_bits),
    .io_argOuts_31_valid(Fringe_io_argOuts_31_valid),
    .io_argOuts_31_bits(Fringe_io_argOuts_31_bits),
    .io_argOuts_32_valid(Fringe_io_argOuts_32_valid),
    .io_argOuts_32_bits(Fringe_io_argOuts_32_bits),
    .io_argOuts_33_valid(Fringe_io_argOuts_33_valid),
    .io_argOuts_33_bits(Fringe_io_argOuts_33_bits),
    .io_argOuts_34_valid(Fringe_io_argOuts_34_valid),
    .io_argOuts_34_bits(Fringe_io_argOuts_34_bits),
    .io_argOuts_35_valid(Fringe_io_argOuts_35_valid),
    .io_argOuts_35_bits(Fringe_io_argOuts_35_bits),
    .io_argOuts_36_valid(Fringe_io_argOuts_36_valid),
    .io_argOuts_36_bits(Fringe_io_argOuts_36_bits),
    .io_argOuts_37_valid(Fringe_io_argOuts_37_valid),
    .io_argOuts_37_bits(Fringe_io_argOuts_37_bits),
    .io_argOuts_38_valid(Fringe_io_argOuts_38_valid),
    .io_argOuts_38_bits(Fringe_io_argOuts_38_bits),
    .io_argOuts_39_valid(Fringe_io_argOuts_39_valid),
    .io_argOuts_39_bits(Fringe_io_argOuts_39_bits),
    .io_argOuts_40_valid(Fringe_io_argOuts_40_valid),
    .io_argOuts_40_bits(Fringe_io_argOuts_40_bits),
    .io_argOuts_41_valid(Fringe_io_argOuts_41_valid),
    .io_argOuts_41_bits(Fringe_io_argOuts_41_bits),
    .io_argOuts_42_valid(Fringe_io_argOuts_42_valid),
    .io_argOuts_42_bits(Fringe_io_argOuts_42_bits),
    .io_argOuts_43_valid(Fringe_io_argOuts_43_valid),
    .io_argOuts_43_bits(Fringe_io_argOuts_43_bits),
    .io_argOuts_44_valid(Fringe_io_argOuts_44_valid),
    .io_argOuts_44_bits(Fringe_io_argOuts_44_bits),
    .io_argOuts_45_valid(Fringe_io_argOuts_45_valid),
    .io_argOuts_45_bits(Fringe_io_argOuts_45_bits),
    .io_argOuts_46_valid(Fringe_io_argOuts_46_valid),
    .io_argOuts_46_bits(Fringe_io_argOuts_46_bits),
    .io_argOuts_47_valid(Fringe_io_argOuts_47_valid),
    .io_argOuts_47_bits(Fringe_io_argOuts_47_bits),
    .io_argOuts_48_valid(Fringe_io_argOuts_48_valid),
    .io_argOuts_48_bits(Fringe_io_argOuts_48_bits),
    .io_argOuts_49_valid(Fringe_io_argOuts_49_valid),
    .io_argOuts_49_bits(Fringe_io_argOuts_49_bits),
    .io_argOuts_50_valid(Fringe_io_argOuts_50_valid),
    .io_argOuts_50_bits(Fringe_io_argOuts_50_bits),
    .io_argOuts_51_valid(Fringe_io_argOuts_51_valid),
    .io_argOuts_51_bits(Fringe_io_argOuts_51_bits),
    .io_argOuts_52_valid(Fringe_io_argOuts_52_valid),
    .io_argOuts_52_bits(Fringe_io_argOuts_52_bits),
    .io_argOuts_53_valid(Fringe_io_argOuts_53_valid),
    .io_argOuts_53_bits(Fringe_io_argOuts_53_bits),
    .io_argOuts_54_valid(Fringe_io_argOuts_54_valid),
    .io_argOuts_54_bits(Fringe_io_argOuts_54_bits),
    .io_argOuts_55_valid(Fringe_io_argOuts_55_valid),
    .io_argOuts_55_bits(Fringe_io_argOuts_55_bits),
    .io_argOuts_56_valid(Fringe_io_argOuts_56_valid),
    .io_argOuts_56_bits(Fringe_io_argOuts_56_bits),
    .io_argOuts_57_valid(Fringe_io_argOuts_57_valid),
    .io_argOuts_57_bits(Fringe_io_argOuts_57_bits),
    .io_argOuts_58_valid(Fringe_io_argOuts_58_valid),
    .io_argOuts_58_bits(Fringe_io_argOuts_58_bits),
    .io_argOuts_59_valid(Fringe_io_argOuts_59_valid),
    .io_argOuts_59_bits(Fringe_io_argOuts_59_bits),
    .io_argEchos_0(Fringe_io_argEchos_0),
    .io_argEchos_1(Fringe_io_argEchos_1),
    .io_argEchos_2(Fringe_io_argEchos_2),
    .io_argEchos_3(Fringe_io_argEchos_3),
    .io_argEchos_4(Fringe_io_argEchos_4),
    .io_argEchos_5(Fringe_io_argEchos_5),
    .io_argEchos_6(Fringe_io_argEchos_6),
    .io_argEchos_7(Fringe_io_argEchos_7),
    .io_argEchos_8(Fringe_io_argEchos_8),
    .io_argEchos_9(Fringe_io_argEchos_9),
    .io_argEchos_10(Fringe_io_argEchos_10),
    .io_argEchos_11(Fringe_io_argEchos_11),
    .io_argEchos_12(Fringe_io_argEchos_12),
    .io_argEchos_13(Fringe_io_argEchos_13),
    .io_argEchos_14(Fringe_io_argEchos_14),
    .io_argEchos_15(Fringe_io_argEchos_15),
    .io_argEchos_16(Fringe_io_argEchos_16),
    .io_argEchos_17(Fringe_io_argEchos_17),
    .io_argEchos_18(Fringe_io_argEchos_18),
    .io_argEchos_19(Fringe_io_argEchos_19),
    .io_argEchos_20(Fringe_io_argEchos_20),
    .io_argEchos_21(Fringe_io_argEchos_21),
    .io_argEchos_22(Fringe_io_argEchos_22),
    .io_argEchos_23(Fringe_io_argEchos_23),
    .io_argEchos_24(Fringe_io_argEchos_24),
    .io_argEchos_25(Fringe_io_argEchos_25),
    .io_argEchos_26(Fringe_io_argEchos_26),
    .io_argEchos_27(Fringe_io_argEchos_27),
    .io_argEchos_28(Fringe_io_argEchos_28),
    .io_argEchos_29(Fringe_io_argEchos_29),
    .io_argEchos_30(Fringe_io_argEchos_30),
    .io_argEchos_31(Fringe_io_argEchos_31),
    .io_argEchos_32(Fringe_io_argEchos_32),
    .io_argEchos_33(Fringe_io_argEchos_33),
    .io_argEchos_34(Fringe_io_argEchos_34),
    .io_argEchos_35(Fringe_io_argEchos_35),
    .io_argEchos_36(Fringe_io_argEchos_36),
    .io_argEchos_37(Fringe_io_argEchos_37),
    .io_argEchos_38(Fringe_io_argEchos_38),
    .io_argEchos_39(Fringe_io_argEchos_39),
    .io_argEchos_40(Fringe_io_argEchos_40),
    .io_argEchos_41(Fringe_io_argEchos_41),
    .io_argEchos_42(Fringe_io_argEchos_42),
    .io_argEchos_43(Fringe_io_argEchos_43),
    .io_argEchos_44(Fringe_io_argEchos_44),
    .io_argEchos_45(Fringe_io_argEchos_45),
    .io_argEchos_46(Fringe_io_argEchos_46),
    .io_argEchos_47(Fringe_io_argEchos_47),
    .io_argEchos_48(Fringe_io_argEchos_48),
    .io_argEchos_49(Fringe_io_argEchos_49),
    .io_argEchos_50(Fringe_io_argEchos_50),
    .io_argEchos_51(Fringe_io_argEchos_51),
    .io_argEchos_52(Fringe_io_argEchos_52),
    .io_argEchos_53(Fringe_io_argEchos_53),
    .io_argEchos_54(Fringe_io_argEchos_54),
    .io_argEchos_55(Fringe_io_argEchos_55),
    .io_argEchos_56(Fringe_io_argEchos_56),
    .io_argEchos_57(Fringe_io_argEchos_57),
    .io_argEchos_58(Fringe_io_argEchos_58),
    .io_argEchos_59(Fringe_io_argEchos_59),
    .io_memStreams_loads_0_cmd_ready(Fringe_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(Fringe_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(Fringe_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(Fringe_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(Fringe_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(Fringe_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(Fringe_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_stores_0_cmd_ready(Fringe_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(Fringe_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(Fringe_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(Fringe_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(Fringe_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(Fringe_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(Fringe_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(Fringe_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(Fringe_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(Fringe_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(Fringe_io_memStreams_stores_0_wresp_bits),
    .io_dram_0_cmd_ready(Fringe_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(Fringe_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(Fringe_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(Fringe_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_rawAddr(Fringe_io_dram_0_cmd_bits_rawAddr),
    .io_dram_0_cmd_bits_isWr(Fringe_io_dram_0_cmd_bits_isWr),
    .io_dram_0_cmd_bits_tag(Fringe_io_dram_0_cmd_bits_tag),
    .io_dram_0_wdata_ready(Fringe_io_dram_0_wdata_ready),
    .io_dram_0_wdata_valid(Fringe_io_dram_0_wdata_valid),
    .io_dram_0_wdata_bits_wdata_0(Fringe_io_dram_0_wdata_bits_wdata_0),
    .io_dram_0_wdata_bits_wdata_1(Fringe_io_dram_0_wdata_bits_wdata_1),
    .io_dram_0_wdata_bits_wdata_2(Fringe_io_dram_0_wdata_bits_wdata_2),
    .io_dram_0_wdata_bits_wdata_3(Fringe_io_dram_0_wdata_bits_wdata_3),
    .io_dram_0_wdata_bits_wdata_4(Fringe_io_dram_0_wdata_bits_wdata_4),
    .io_dram_0_wdata_bits_wdata_5(Fringe_io_dram_0_wdata_bits_wdata_5),
    .io_dram_0_wdata_bits_wdata_6(Fringe_io_dram_0_wdata_bits_wdata_6),
    .io_dram_0_wdata_bits_wdata_7(Fringe_io_dram_0_wdata_bits_wdata_7),
    .io_dram_0_wdata_bits_wdata_8(Fringe_io_dram_0_wdata_bits_wdata_8),
    .io_dram_0_wdata_bits_wdata_9(Fringe_io_dram_0_wdata_bits_wdata_9),
    .io_dram_0_wdata_bits_wdata_10(Fringe_io_dram_0_wdata_bits_wdata_10),
    .io_dram_0_wdata_bits_wdata_11(Fringe_io_dram_0_wdata_bits_wdata_11),
    .io_dram_0_wdata_bits_wdata_12(Fringe_io_dram_0_wdata_bits_wdata_12),
    .io_dram_0_wdata_bits_wdata_13(Fringe_io_dram_0_wdata_bits_wdata_13),
    .io_dram_0_wdata_bits_wdata_14(Fringe_io_dram_0_wdata_bits_wdata_14),
    .io_dram_0_wdata_bits_wdata_15(Fringe_io_dram_0_wdata_bits_wdata_15),
    .io_dram_0_wdata_bits_wdata_16(Fringe_io_dram_0_wdata_bits_wdata_16),
    .io_dram_0_wdata_bits_wdata_17(Fringe_io_dram_0_wdata_bits_wdata_17),
    .io_dram_0_wdata_bits_wdata_18(Fringe_io_dram_0_wdata_bits_wdata_18),
    .io_dram_0_wdata_bits_wdata_19(Fringe_io_dram_0_wdata_bits_wdata_19),
    .io_dram_0_wdata_bits_wdata_20(Fringe_io_dram_0_wdata_bits_wdata_20),
    .io_dram_0_wdata_bits_wdata_21(Fringe_io_dram_0_wdata_bits_wdata_21),
    .io_dram_0_wdata_bits_wdata_22(Fringe_io_dram_0_wdata_bits_wdata_22),
    .io_dram_0_wdata_bits_wdata_23(Fringe_io_dram_0_wdata_bits_wdata_23),
    .io_dram_0_wdata_bits_wdata_24(Fringe_io_dram_0_wdata_bits_wdata_24),
    .io_dram_0_wdata_bits_wdata_25(Fringe_io_dram_0_wdata_bits_wdata_25),
    .io_dram_0_wdata_bits_wdata_26(Fringe_io_dram_0_wdata_bits_wdata_26),
    .io_dram_0_wdata_bits_wdata_27(Fringe_io_dram_0_wdata_bits_wdata_27),
    .io_dram_0_wdata_bits_wdata_28(Fringe_io_dram_0_wdata_bits_wdata_28),
    .io_dram_0_wdata_bits_wdata_29(Fringe_io_dram_0_wdata_bits_wdata_29),
    .io_dram_0_wdata_bits_wdata_30(Fringe_io_dram_0_wdata_bits_wdata_30),
    .io_dram_0_wdata_bits_wdata_31(Fringe_io_dram_0_wdata_bits_wdata_31),
    .io_dram_0_wdata_bits_wdata_32(Fringe_io_dram_0_wdata_bits_wdata_32),
    .io_dram_0_wdata_bits_wdata_33(Fringe_io_dram_0_wdata_bits_wdata_33),
    .io_dram_0_wdata_bits_wdata_34(Fringe_io_dram_0_wdata_bits_wdata_34),
    .io_dram_0_wdata_bits_wdata_35(Fringe_io_dram_0_wdata_bits_wdata_35),
    .io_dram_0_wdata_bits_wdata_36(Fringe_io_dram_0_wdata_bits_wdata_36),
    .io_dram_0_wdata_bits_wdata_37(Fringe_io_dram_0_wdata_bits_wdata_37),
    .io_dram_0_wdata_bits_wdata_38(Fringe_io_dram_0_wdata_bits_wdata_38),
    .io_dram_0_wdata_bits_wdata_39(Fringe_io_dram_0_wdata_bits_wdata_39),
    .io_dram_0_wdata_bits_wdata_40(Fringe_io_dram_0_wdata_bits_wdata_40),
    .io_dram_0_wdata_bits_wdata_41(Fringe_io_dram_0_wdata_bits_wdata_41),
    .io_dram_0_wdata_bits_wdata_42(Fringe_io_dram_0_wdata_bits_wdata_42),
    .io_dram_0_wdata_bits_wdata_43(Fringe_io_dram_0_wdata_bits_wdata_43),
    .io_dram_0_wdata_bits_wdata_44(Fringe_io_dram_0_wdata_bits_wdata_44),
    .io_dram_0_wdata_bits_wdata_45(Fringe_io_dram_0_wdata_bits_wdata_45),
    .io_dram_0_wdata_bits_wdata_46(Fringe_io_dram_0_wdata_bits_wdata_46),
    .io_dram_0_wdata_bits_wdata_47(Fringe_io_dram_0_wdata_bits_wdata_47),
    .io_dram_0_wdata_bits_wdata_48(Fringe_io_dram_0_wdata_bits_wdata_48),
    .io_dram_0_wdata_bits_wdata_49(Fringe_io_dram_0_wdata_bits_wdata_49),
    .io_dram_0_wdata_bits_wdata_50(Fringe_io_dram_0_wdata_bits_wdata_50),
    .io_dram_0_wdata_bits_wdata_51(Fringe_io_dram_0_wdata_bits_wdata_51),
    .io_dram_0_wdata_bits_wdata_52(Fringe_io_dram_0_wdata_bits_wdata_52),
    .io_dram_0_wdata_bits_wdata_53(Fringe_io_dram_0_wdata_bits_wdata_53),
    .io_dram_0_wdata_bits_wdata_54(Fringe_io_dram_0_wdata_bits_wdata_54),
    .io_dram_0_wdata_bits_wdata_55(Fringe_io_dram_0_wdata_bits_wdata_55),
    .io_dram_0_wdata_bits_wdata_56(Fringe_io_dram_0_wdata_bits_wdata_56),
    .io_dram_0_wdata_bits_wdata_57(Fringe_io_dram_0_wdata_bits_wdata_57),
    .io_dram_0_wdata_bits_wdata_58(Fringe_io_dram_0_wdata_bits_wdata_58),
    .io_dram_0_wdata_bits_wdata_59(Fringe_io_dram_0_wdata_bits_wdata_59),
    .io_dram_0_wdata_bits_wdata_60(Fringe_io_dram_0_wdata_bits_wdata_60),
    .io_dram_0_wdata_bits_wdata_61(Fringe_io_dram_0_wdata_bits_wdata_61),
    .io_dram_0_wdata_bits_wdata_62(Fringe_io_dram_0_wdata_bits_wdata_62),
    .io_dram_0_wdata_bits_wdata_63(Fringe_io_dram_0_wdata_bits_wdata_63),
    .io_dram_0_wdata_bits_wstrb_0(Fringe_io_dram_0_wdata_bits_wstrb_0),
    .io_dram_0_wdata_bits_wstrb_1(Fringe_io_dram_0_wdata_bits_wstrb_1),
    .io_dram_0_wdata_bits_wstrb_2(Fringe_io_dram_0_wdata_bits_wstrb_2),
    .io_dram_0_wdata_bits_wstrb_3(Fringe_io_dram_0_wdata_bits_wstrb_3),
    .io_dram_0_wdata_bits_wstrb_4(Fringe_io_dram_0_wdata_bits_wstrb_4),
    .io_dram_0_wdata_bits_wstrb_5(Fringe_io_dram_0_wdata_bits_wstrb_5),
    .io_dram_0_wdata_bits_wstrb_6(Fringe_io_dram_0_wdata_bits_wstrb_6),
    .io_dram_0_wdata_bits_wstrb_7(Fringe_io_dram_0_wdata_bits_wstrb_7),
    .io_dram_0_wdata_bits_wstrb_8(Fringe_io_dram_0_wdata_bits_wstrb_8),
    .io_dram_0_wdata_bits_wstrb_9(Fringe_io_dram_0_wdata_bits_wstrb_9),
    .io_dram_0_wdata_bits_wstrb_10(Fringe_io_dram_0_wdata_bits_wstrb_10),
    .io_dram_0_wdata_bits_wstrb_11(Fringe_io_dram_0_wdata_bits_wstrb_11),
    .io_dram_0_wdata_bits_wstrb_12(Fringe_io_dram_0_wdata_bits_wstrb_12),
    .io_dram_0_wdata_bits_wstrb_13(Fringe_io_dram_0_wdata_bits_wstrb_13),
    .io_dram_0_wdata_bits_wstrb_14(Fringe_io_dram_0_wdata_bits_wstrb_14),
    .io_dram_0_wdata_bits_wstrb_15(Fringe_io_dram_0_wdata_bits_wstrb_15),
    .io_dram_0_wdata_bits_wstrb_16(Fringe_io_dram_0_wdata_bits_wstrb_16),
    .io_dram_0_wdata_bits_wstrb_17(Fringe_io_dram_0_wdata_bits_wstrb_17),
    .io_dram_0_wdata_bits_wstrb_18(Fringe_io_dram_0_wdata_bits_wstrb_18),
    .io_dram_0_wdata_bits_wstrb_19(Fringe_io_dram_0_wdata_bits_wstrb_19),
    .io_dram_0_wdata_bits_wstrb_20(Fringe_io_dram_0_wdata_bits_wstrb_20),
    .io_dram_0_wdata_bits_wstrb_21(Fringe_io_dram_0_wdata_bits_wstrb_21),
    .io_dram_0_wdata_bits_wstrb_22(Fringe_io_dram_0_wdata_bits_wstrb_22),
    .io_dram_0_wdata_bits_wstrb_23(Fringe_io_dram_0_wdata_bits_wstrb_23),
    .io_dram_0_wdata_bits_wstrb_24(Fringe_io_dram_0_wdata_bits_wstrb_24),
    .io_dram_0_wdata_bits_wstrb_25(Fringe_io_dram_0_wdata_bits_wstrb_25),
    .io_dram_0_wdata_bits_wstrb_26(Fringe_io_dram_0_wdata_bits_wstrb_26),
    .io_dram_0_wdata_bits_wstrb_27(Fringe_io_dram_0_wdata_bits_wstrb_27),
    .io_dram_0_wdata_bits_wstrb_28(Fringe_io_dram_0_wdata_bits_wstrb_28),
    .io_dram_0_wdata_bits_wstrb_29(Fringe_io_dram_0_wdata_bits_wstrb_29),
    .io_dram_0_wdata_bits_wstrb_30(Fringe_io_dram_0_wdata_bits_wstrb_30),
    .io_dram_0_wdata_bits_wstrb_31(Fringe_io_dram_0_wdata_bits_wstrb_31),
    .io_dram_0_wdata_bits_wstrb_32(Fringe_io_dram_0_wdata_bits_wstrb_32),
    .io_dram_0_wdata_bits_wstrb_33(Fringe_io_dram_0_wdata_bits_wstrb_33),
    .io_dram_0_wdata_bits_wstrb_34(Fringe_io_dram_0_wdata_bits_wstrb_34),
    .io_dram_0_wdata_bits_wstrb_35(Fringe_io_dram_0_wdata_bits_wstrb_35),
    .io_dram_0_wdata_bits_wstrb_36(Fringe_io_dram_0_wdata_bits_wstrb_36),
    .io_dram_0_wdata_bits_wstrb_37(Fringe_io_dram_0_wdata_bits_wstrb_37),
    .io_dram_0_wdata_bits_wstrb_38(Fringe_io_dram_0_wdata_bits_wstrb_38),
    .io_dram_0_wdata_bits_wstrb_39(Fringe_io_dram_0_wdata_bits_wstrb_39),
    .io_dram_0_wdata_bits_wstrb_40(Fringe_io_dram_0_wdata_bits_wstrb_40),
    .io_dram_0_wdata_bits_wstrb_41(Fringe_io_dram_0_wdata_bits_wstrb_41),
    .io_dram_0_wdata_bits_wstrb_42(Fringe_io_dram_0_wdata_bits_wstrb_42),
    .io_dram_0_wdata_bits_wstrb_43(Fringe_io_dram_0_wdata_bits_wstrb_43),
    .io_dram_0_wdata_bits_wstrb_44(Fringe_io_dram_0_wdata_bits_wstrb_44),
    .io_dram_0_wdata_bits_wstrb_45(Fringe_io_dram_0_wdata_bits_wstrb_45),
    .io_dram_0_wdata_bits_wstrb_46(Fringe_io_dram_0_wdata_bits_wstrb_46),
    .io_dram_0_wdata_bits_wstrb_47(Fringe_io_dram_0_wdata_bits_wstrb_47),
    .io_dram_0_wdata_bits_wstrb_48(Fringe_io_dram_0_wdata_bits_wstrb_48),
    .io_dram_0_wdata_bits_wstrb_49(Fringe_io_dram_0_wdata_bits_wstrb_49),
    .io_dram_0_wdata_bits_wstrb_50(Fringe_io_dram_0_wdata_bits_wstrb_50),
    .io_dram_0_wdata_bits_wstrb_51(Fringe_io_dram_0_wdata_bits_wstrb_51),
    .io_dram_0_wdata_bits_wstrb_52(Fringe_io_dram_0_wdata_bits_wstrb_52),
    .io_dram_0_wdata_bits_wstrb_53(Fringe_io_dram_0_wdata_bits_wstrb_53),
    .io_dram_0_wdata_bits_wstrb_54(Fringe_io_dram_0_wdata_bits_wstrb_54),
    .io_dram_0_wdata_bits_wstrb_55(Fringe_io_dram_0_wdata_bits_wstrb_55),
    .io_dram_0_wdata_bits_wstrb_56(Fringe_io_dram_0_wdata_bits_wstrb_56),
    .io_dram_0_wdata_bits_wstrb_57(Fringe_io_dram_0_wdata_bits_wstrb_57),
    .io_dram_0_wdata_bits_wstrb_58(Fringe_io_dram_0_wdata_bits_wstrb_58),
    .io_dram_0_wdata_bits_wstrb_59(Fringe_io_dram_0_wdata_bits_wstrb_59),
    .io_dram_0_wdata_bits_wstrb_60(Fringe_io_dram_0_wdata_bits_wstrb_60),
    .io_dram_0_wdata_bits_wstrb_61(Fringe_io_dram_0_wdata_bits_wstrb_61),
    .io_dram_0_wdata_bits_wstrb_62(Fringe_io_dram_0_wdata_bits_wstrb_62),
    .io_dram_0_wdata_bits_wstrb_63(Fringe_io_dram_0_wdata_bits_wstrb_63),
    .io_dram_0_wdata_bits_wlast(Fringe_io_dram_0_wdata_bits_wlast),
    .io_dram_0_rresp_ready(Fringe_io_dram_0_rresp_ready),
    .io_dram_0_rresp_valid(Fringe_io_dram_0_rresp_valid),
    .io_dram_0_rresp_bits_rdata_0(Fringe_io_dram_0_rresp_bits_rdata_0),
    .io_dram_0_rresp_bits_rdata_1(Fringe_io_dram_0_rresp_bits_rdata_1),
    .io_dram_0_rresp_bits_rdata_2(Fringe_io_dram_0_rresp_bits_rdata_2),
    .io_dram_0_rresp_bits_rdata_3(Fringe_io_dram_0_rresp_bits_rdata_3),
    .io_dram_0_rresp_bits_rdata_4(Fringe_io_dram_0_rresp_bits_rdata_4),
    .io_dram_0_rresp_bits_rdata_5(Fringe_io_dram_0_rresp_bits_rdata_5),
    .io_dram_0_rresp_bits_rdata_6(Fringe_io_dram_0_rresp_bits_rdata_6),
    .io_dram_0_rresp_bits_rdata_7(Fringe_io_dram_0_rresp_bits_rdata_7),
    .io_dram_0_rresp_bits_rdata_8(Fringe_io_dram_0_rresp_bits_rdata_8),
    .io_dram_0_rresp_bits_rdata_9(Fringe_io_dram_0_rresp_bits_rdata_9),
    .io_dram_0_rresp_bits_rdata_10(Fringe_io_dram_0_rresp_bits_rdata_10),
    .io_dram_0_rresp_bits_rdata_11(Fringe_io_dram_0_rresp_bits_rdata_11),
    .io_dram_0_rresp_bits_rdata_12(Fringe_io_dram_0_rresp_bits_rdata_12),
    .io_dram_0_rresp_bits_rdata_13(Fringe_io_dram_0_rresp_bits_rdata_13),
    .io_dram_0_rresp_bits_rdata_14(Fringe_io_dram_0_rresp_bits_rdata_14),
    .io_dram_0_rresp_bits_rdata_15(Fringe_io_dram_0_rresp_bits_rdata_15),
    .io_dram_0_rresp_bits_rdata_16(Fringe_io_dram_0_rresp_bits_rdata_16),
    .io_dram_0_rresp_bits_rdata_17(Fringe_io_dram_0_rresp_bits_rdata_17),
    .io_dram_0_rresp_bits_rdata_18(Fringe_io_dram_0_rresp_bits_rdata_18),
    .io_dram_0_rresp_bits_rdata_19(Fringe_io_dram_0_rresp_bits_rdata_19),
    .io_dram_0_rresp_bits_rdata_20(Fringe_io_dram_0_rresp_bits_rdata_20),
    .io_dram_0_rresp_bits_rdata_21(Fringe_io_dram_0_rresp_bits_rdata_21),
    .io_dram_0_rresp_bits_rdata_22(Fringe_io_dram_0_rresp_bits_rdata_22),
    .io_dram_0_rresp_bits_rdata_23(Fringe_io_dram_0_rresp_bits_rdata_23),
    .io_dram_0_rresp_bits_rdata_24(Fringe_io_dram_0_rresp_bits_rdata_24),
    .io_dram_0_rresp_bits_rdata_25(Fringe_io_dram_0_rresp_bits_rdata_25),
    .io_dram_0_rresp_bits_rdata_26(Fringe_io_dram_0_rresp_bits_rdata_26),
    .io_dram_0_rresp_bits_rdata_27(Fringe_io_dram_0_rresp_bits_rdata_27),
    .io_dram_0_rresp_bits_rdata_28(Fringe_io_dram_0_rresp_bits_rdata_28),
    .io_dram_0_rresp_bits_rdata_29(Fringe_io_dram_0_rresp_bits_rdata_29),
    .io_dram_0_rresp_bits_rdata_30(Fringe_io_dram_0_rresp_bits_rdata_30),
    .io_dram_0_rresp_bits_rdata_31(Fringe_io_dram_0_rresp_bits_rdata_31),
    .io_dram_0_rresp_bits_rdata_32(Fringe_io_dram_0_rresp_bits_rdata_32),
    .io_dram_0_rresp_bits_rdata_33(Fringe_io_dram_0_rresp_bits_rdata_33),
    .io_dram_0_rresp_bits_rdata_34(Fringe_io_dram_0_rresp_bits_rdata_34),
    .io_dram_0_rresp_bits_rdata_35(Fringe_io_dram_0_rresp_bits_rdata_35),
    .io_dram_0_rresp_bits_rdata_36(Fringe_io_dram_0_rresp_bits_rdata_36),
    .io_dram_0_rresp_bits_rdata_37(Fringe_io_dram_0_rresp_bits_rdata_37),
    .io_dram_0_rresp_bits_rdata_38(Fringe_io_dram_0_rresp_bits_rdata_38),
    .io_dram_0_rresp_bits_rdata_39(Fringe_io_dram_0_rresp_bits_rdata_39),
    .io_dram_0_rresp_bits_rdata_40(Fringe_io_dram_0_rresp_bits_rdata_40),
    .io_dram_0_rresp_bits_rdata_41(Fringe_io_dram_0_rresp_bits_rdata_41),
    .io_dram_0_rresp_bits_rdata_42(Fringe_io_dram_0_rresp_bits_rdata_42),
    .io_dram_0_rresp_bits_rdata_43(Fringe_io_dram_0_rresp_bits_rdata_43),
    .io_dram_0_rresp_bits_rdata_44(Fringe_io_dram_0_rresp_bits_rdata_44),
    .io_dram_0_rresp_bits_rdata_45(Fringe_io_dram_0_rresp_bits_rdata_45),
    .io_dram_0_rresp_bits_rdata_46(Fringe_io_dram_0_rresp_bits_rdata_46),
    .io_dram_0_rresp_bits_rdata_47(Fringe_io_dram_0_rresp_bits_rdata_47),
    .io_dram_0_rresp_bits_rdata_48(Fringe_io_dram_0_rresp_bits_rdata_48),
    .io_dram_0_rresp_bits_rdata_49(Fringe_io_dram_0_rresp_bits_rdata_49),
    .io_dram_0_rresp_bits_rdata_50(Fringe_io_dram_0_rresp_bits_rdata_50),
    .io_dram_0_rresp_bits_rdata_51(Fringe_io_dram_0_rresp_bits_rdata_51),
    .io_dram_0_rresp_bits_rdata_52(Fringe_io_dram_0_rresp_bits_rdata_52),
    .io_dram_0_rresp_bits_rdata_53(Fringe_io_dram_0_rresp_bits_rdata_53),
    .io_dram_0_rresp_bits_rdata_54(Fringe_io_dram_0_rresp_bits_rdata_54),
    .io_dram_0_rresp_bits_rdata_55(Fringe_io_dram_0_rresp_bits_rdata_55),
    .io_dram_0_rresp_bits_rdata_56(Fringe_io_dram_0_rresp_bits_rdata_56),
    .io_dram_0_rresp_bits_rdata_57(Fringe_io_dram_0_rresp_bits_rdata_57),
    .io_dram_0_rresp_bits_rdata_58(Fringe_io_dram_0_rresp_bits_rdata_58),
    .io_dram_0_rresp_bits_rdata_59(Fringe_io_dram_0_rresp_bits_rdata_59),
    .io_dram_0_rresp_bits_rdata_60(Fringe_io_dram_0_rresp_bits_rdata_60),
    .io_dram_0_rresp_bits_rdata_61(Fringe_io_dram_0_rresp_bits_rdata_61),
    .io_dram_0_rresp_bits_rdata_62(Fringe_io_dram_0_rresp_bits_rdata_62),
    .io_dram_0_rresp_bits_rdata_63(Fringe_io_dram_0_rresp_bits_rdata_63),
    .io_dram_0_rresp_bits_tag(Fringe_io_dram_0_rresp_bits_tag),
    .io_dram_0_wresp_ready(Fringe_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(Fringe_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag(Fringe_io_dram_0_wresp_bits_tag),
    .io_heap_0_req_valid(Fringe_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(Fringe_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(Fringe_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(Fringe_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(Fringe_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(Fringe_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = Fringe_io_rdata; // @[SimTarget.scala 24:14:@158998.4]
  assign io_dram_0_cmd_valid = Fringe_io_dram_0_cmd_valid; // @[SimTarget.scala 27:13:@159205.4]
  assign io_dram_0_cmd_bits_addr = Fringe_io_dram_0_cmd_bits_addr; // @[SimTarget.scala 27:13:@159204.4]
  assign io_dram_0_cmd_bits_size = Fringe_io_dram_0_cmd_bits_size; // @[SimTarget.scala 27:13:@159203.4]
  assign io_dram_0_cmd_bits_rawAddr = Fringe_io_dram_0_cmd_bits_rawAddr; // @[SimTarget.scala 27:13:@159202.4]
  assign io_dram_0_cmd_bits_isWr = Fringe_io_dram_0_cmd_bits_isWr; // @[SimTarget.scala 27:13:@159201.4]
  assign io_dram_0_cmd_bits_tag = Fringe_io_dram_0_cmd_bits_tag; // @[SimTarget.scala 27:13:@159200.4]
  assign io_dram_0_wdata_valid = Fringe_io_dram_0_wdata_valid; // @[SimTarget.scala 27:13:@159198.4]
  assign io_dram_0_wdata_bits_wdata_0 = Fringe_io_dram_0_wdata_bits_wdata_0; // @[SimTarget.scala 27:13:@159134.4]
  assign io_dram_0_wdata_bits_wdata_1 = Fringe_io_dram_0_wdata_bits_wdata_1; // @[SimTarget.scala 27:13:@159135.4]
  assign io_dram_0_wdata_bits_wdata_2 = Fringe_io_dram_0_wdata_bits_wdata_2; // @[SimTarget.scala 27:13:@159136.4]
  assign io_dram_0_wdata_bits_wdata_3 = Fringe_io_dram_0_wdata_bits_wdata_3; // @[SimTarget.scala 27:13:@159137.4]
  assign io_dram_0_wdata_bits_wdata_4 = Fringe_io_dram_0_wdata_bits_wdata_4; // @[SimTarget.scala 27:13:@159138.4]
  assign io_dram_0_wdata_bits_wdata_5 = Fringe_io_dram_0_wdata_bits_wdata_5; // @[SimTarget.scala 27:13:@159139.4]
  assign io_dram_0_wdata_bits_wdata_6 = Fringe_io_dram_0_wdata_bits_wdata_6; // @[SimTarget.scala 27:13:@159140.4]
  assign io_dram_0_wdata_bits_wdata_7 = Fringe_io_dram_0_wdata_bits_wdata_7; // @[SimTarget.scala 27:13:@159141.4]
  assign io_dram_0_wdata_bits_wdata_8 = Fringe_io_dram_0_wdata_bits_wdata_8; // @[SimTarget.scala 27:13:@159142.4]
  assign io_dram_0_wdata_bits_wdata_9 = Fringe_io_dram_0_wdata_bits_wdata_9; // @[SimTarget.scala 27:13:@159143.4]
  assign io_dram_0_wdata_bits_wdata_10 = Fringe_io_dram_0_wdata_bits_wdata_10; // @[SimTarget.scala 27:13:@159144.4]
  assign io_dram_0_wdata_bits_wdata_11 = Fringe_io_dram_0_wdata_bits_wdata_11; // @[SimTarget.scala 27:13:@159145.4]
  assign io_dram_0_wdata_bits_wdata_12 = Fringe_io_dram_0_wdata_bits_wdata_12; // @[SimTarget.scala 27:13:@159146.4]
  assign io_dram_0_wdata_bits_wdata_13 = Fringe_io_dram_0_wdata_bits_wdata_13; // @[SimTarget.scala 27:13:@159147.4]
  assign io_dram_0_wdata_bits_wdata_14 = Fringe_io_dram_0_wdata_bits_wdata_14; // @[SimTarget.scala 27:13:@159148.4]
  assign io_dram_0_wdata_bits_wdata_15 = Fringe_io_dram_0_wdata_bits_wdata_15; // @[SimTarget.scala 27:13:@159149.4]
  assign io_dram_0_wdata_bits_wdata_16 = Fringe_io_dram_0_wdata_bits_wdata_16; // @[SimTarget.scala 27:13:@159150.4]
  assign io_dram_0_wdata_bits_wdata_17 = Fringe_io_dram_0_wdata_bits_wdata_17; // @[SimTarget.scala 27:13:@159151.4]
  assign io_dram_0_wdata_bits_wdata_18 = Fringe_io_dram_0_wdata_bits_wdata_18; // @[SimTarget.scala 27:13:@159152.4]
  assign io_dram_0_wdata_bits_wdata_19 = Fringe_io_dram_0_wdata_bits_wdata_19; // @[SimTarget.scala 27:13:@159153.4]
  assign io_dram_0_wdata_bits_wdata_20 = Fringe_io_dram_0_wdata_bits_wdata_20; // @[SimTarget.scala 27:13:@159154.4]
  assign io_dram_0_wdata_bits_wdata_21 = Fringe_io_dram_0_wdata_bits_wdata_21; // @[SimTarget.scala 27:13:@159155.4]
  assign io_dram_0_wdata_bits_wdata_22 = Fringe_io_dram_0_wdata_bits_wdata_22; // @[SimTarget.scala 27:13:@159156.4]
  assign io_dram_0_wdata_bits_wdata_23 = Fringe_io_dram_0_wdata_bits_wdata_23; // @[SimTarget.scala 27:13:@159157.4]
  assign io_dram_0_wdata_bits_wdata_24 = Fringe_io_dram_0_wdata_bits_wdata_24; // @[SimTarget.scala 27:13:@159158.4]
  assign io_dram_0_wdata_bits_wdata_25 = Fringe_io_dram_0_wdata_bits_wdata_25; // @[SimTarget.scala 27:13:@159159.4]
  assign io_dram_0_wdata_bits_wdata_26 = Fringe_io_dram_0_wdata_bits_wdata_26; // @[SimTarget.scala 27:13:@159160.4]
  assign io_dram_0_wdata_bits_wdata_27 = Fringe_io_dram_0_wdata_bits_wdata_27; // @[SimTarget.scala 27:13:@159161.4]
  assign io_dram_0_wdata_bits_wdata_28 = Fringe_io_dram_0_wdata_bits_wdata_28; // @[SimTarget.scala 27:13:@159162.4]
  assign io_dram_0_wdata_bits_wdata_29 = Fringe_io_dram_0_wdata_bits_wdata_29; // @[SimTarget.scala 27:13:@159163.4]
  assign io_dram_0_wdata_bits_wdata_30 = Fringe_io_dram_0_wdata_bits_wdata_30; // @[SimTarget.scala 27:13:@159164.4]
  assign io_dram_0_wdata_bits_wdata_31 = Fringe_io_dram_0_wdata_bits_wdata_31; // @[SimTarget.scala 27:13:@159165.4]
  assign io_dram_0_wdata_bits_wdata_32 = Fringe_io_dram_0_wdata_bits_wdata_32; // @[SimTarget.scala 27:13:@159166.4]
  assign io_dram_0_wdata_bits_wdata_33 = Fringe_io_dram_0_wdata_bits_wdata_33; // @[SimTarget.scala 27:13:@159167.4]
  assign io_dram_0_wdata_bits_wdata_34 = Fringe_io_dram_0_wdata_bits_wdata_34; // @[SimTarget.scala 27:13:@159168.4]
  assign io_dram_0_wdata_bits_wdata_35 = Fringe_io_dram_0_wdata_bits_wdata_35; // @[SimTarget.scala 27:13:@159169.4]
  assign io_dram_0_wdata_bits_wdata_36 = Fringe_io_dram_0_wdata_bits_wdata_36; // @[SimTarget.scala 27:13:@159170.4]
  assign io_dram_0_wdata_bits_wdata_37 = Fringe_io_dram_0_wdata_bits_wdata_37; // @[SimTarget.scala 27:13:@159171.4]
  assign io_dram_0_wdata_bits_wdata_38 = Fringe_io_dram_0_wdata_bits_wdata_38; // @[SimTarget.scala 27:13:@159172.4]
  assign io_dram_0_wdata_bits_wdata_39 = Fringe_io_dram_0_wdata_bits_wdata_39; // @[SimTarget.scala 27:13:@159173.4]
  assign io_dram_0_wdata_bits_wdata_40 = Fringe_io_dram_0_wdata_bits_wdata_40; // @[SimTarget.scala 27:13:@159174.4]
  assign io_dram_0_wdata_bits_wdata_41 = Fringe_io_dram_0_wdata_bits_wdata_41; // @[SimTarget.scala 27:13:@159175.4]
  assign io_dram_0_wdata_bits_wdata_42 = Fringe_io_dram_0_wdata_bits_wdata_42; // @[SimTarget.scala 27:13:@159176.4]
  assign io_dram_0_wdata_bits_wdata_43 = Fringe_io_dram_0_wdata_bits_wdata_43; // @[SimTarget.scala 27:13:@159177.4]
  assign io_dram_0_wdata_bits_wdata_44 = Fringe_io_dram_0_wdata_bits_wdata_44; // @[SimTarget.scala 27:13:@159178.4]
  assign io_dram_0_wdata_bits_wdata_45 = Fringe_io_dram_0_wdata_bits_wdata_45; // @[SimTarget.scala 27:13:@159179.4]
  assign io_dram_0_wdata_bits_wdata_46 = Fringe_io_dram_0_wdata_bits_wdata_46; // @[SimTarget.scala 27:13:@159180.4]
  assign io_dram_0_wdata_bits_wdata_47 = Fringe_io_dram_0_wdata_bits_wdata_47; // @[SimTarget.scala 27:13:@159181.4]
  assign io_dram_0_wdata_bits_wdata_48 = Fringe_io_dram_0_wdata_bits_wdata_48; // @[SimTarget.scala 27:13:@159182.4]
  assign io_dram_0_wdata_bits_wdata_49 = Fringe_io_dram_0_wdata_bits_wdata_49; // @[SimTarget.scala 27:13:@159183.4]
  assign io_dram_0_wdata_bits_wdata_50 = Fringe_io_dram_0_wdata_bits_wdata_50; // @[SimTarget.scala 27:13:@159184.4]
  assign io_dram_0_wdata_bits_wdata_51 = Fringe_io_dram_0_wdata_bits_wdata_51; // @[SimTarget.scala 27:13:@159185.4]
  assign io_dram_0_wdata_bits_wdata_52 = Fringe_io_dram_0_wdata_bits_wdata_52; // @[SimTarget.scala 27:13:@159186.4]
  assign io_dram_0_wdata_bits_wdata_53 = Fringe_io_dram_0_wdata_bits_wdata_53; // @[SimTarget.scala 27:13:@159187.4]
  assign io_dram_0_wdata_bits_wdata_54 = Fringe_io_dram_0_wdata_bits_wdata_54; // @[SimTarget.scala 27:13:@159188.4]
  assign io_dram_0_wdata_bits_wdata_55 = Fringe_io_dram_0_wdata_bits_wdata_55; // @[SimTarget.scala 27:13:@159189.4]
  assign io_dram_0_wdata_bits_wdata_56 = Fringe_io_dram_0_wdata_bits_wdata_56; // @[SimTarget.scala 27:13:@159190.4]
  assign io_dram_0_wdata_bits_wdata_57 = Fringe_io_dram_0_wdata_bits_wdata_57; // @[SimTarget.scala 27:13:@159191.4]
  assign io_dram_0_wdata_bits_wdata_58 = Fringe_io_dram_0_wdata_bits_wdata_58; // @[SimTarget.scala 27:13:@159192.4]
  assign io_dram_0_wdata_bits_wdata_59 = Fringe_io_dram_0_wdata_bits_wdata_59; // @[SimTarget.scala 27:13:@159193.4]
  assign io_dram_0_wdata_bits_wdata_60 = Fringe_io_dram_0_wdata_bits_wdata_60; // @[SimTarget.scala 27:13:@159194.4]
  assign io_dram_0_wdata_bits_wdata_61 = Fringe_io_dram_0_wdata_bits_wdata_61; // @[SimTarget.scala 27:13:@159195.4]
  assign io_dram_0_wdata_bits_wdata_62 = Fringe_io_dram_0_wdata_bits_wdata_62; // @[SimTarget.scala 27:13:@159196.4]
  assign io_dram_0_wdata_bits_wdata_63 = Fringe_io_dram_0_wdata_bits_wdata_63; // @[SimTarget.scala 27:13:@159197.4]
  assign io_dram_0_wdata_bits_wstrb_0 = Fringe_io_dram_0_wdata_bits_wstrb_0; // @[SimTarget.scala 27:13:@159070.4]
  assign io_dram_0_wdata_bits_wstrb_1 = Fringe_io_dram_0_wdata_bits_wstrb_1; // @[SimTarget.scala 27:13:@159071.4]
  assign io_dram_0_wdata_bits_wstrb_2 = Fringe_io_dram_0_wdata_bits_wstrb_2; // @[SimTarget.scala 27:13:@159072.4]
  assign io_dram_0_wdata_bits_wstrb_3 = Fringe_io_dram_0_wdata_bits_wstrb_3; // @[SimTarget.scala 27:13:@159073.4]
  assign io_dram_0_wdata_bits_wstrb_4 = Fringe_io_dram_0_wdata_bits_wstrb_4; // @[SimTarget.scala 27:13:@159074.4]
  assign io_dram_0_wdata_bits_wstrb_5 = Fringe_io_dram_0_wdata_bits_wstrb_5; // @[SimTarget.scala 27:13:@159075.4]
  assign io_dram_0_wdata_bits_wstrb_6 = Fringe_io_dram_0_wdata_bits_wstrb_6; // @[SimTarget.scala 27:13:@159076.4]
  assign io_dram_0_wdata_bits_wstrb_7 = Fringe_io_dram_0_wdata_bits_wstrb_7; // @[SimTarget.scala 27:13:@159077.4]
  assign io_dram_0_wdata_bits_wstrb_8 = Fringe_io_dram_0_wdata_bits_wstrb_8; // @[SimTarget.scala 27:13:@159078.4]
  assign io_dram_0_wdata_bits_wstrb_9 = Fringe_io_dram_0_wdata_bits_wstrb_9; // @[SimTarget.scala 27:13:@159079.4]
  assign io_dram_0_wdata_bits_wstrb_10 = Fringe_io_dram_0_wdata_bits_wstrb_10; // @[SimTarget.scala 27:13:@159080.4]
  assign io_dram_0_wdata_bits_wstrb_11 = Fringe_io_dram_0_wdata_bits_wstrb_11; // @[SimTarget.scala 27:13:@159081.4]
  assign io_dram_0_wdata_bits_wstrb_12 = Fringe_io_dram_0_wdata_bits_wstrb_12; // @[SimTarget.scala 27:13:@159082.4]
  assign io_dram_0_wdata_bits_wstrb_13 = Fringe_io_dram_0_wdata_bits_wstrb_13; // @[SimTarget.scala 27:13:@159083.4]
  assign io_dram_0_wdata_bits_wstrb_14 = Fringe_io_dram_0_wdata_bits_wstrb_14; // @[SimTarget.scala 27:13:@159084.4]
  assign io_dram_0_wdata_bits_wstrb_15 = Fringe_io_dram_0_wdata_bits_wstrb_15; // @[SimTarget.scala 27:13:@159085.4]
  assign io_dram_0_wdata_bits_wstrb_16 = Fringe_io_dram_0_wdata_bits_wstrb_16; // @[SimTarget.scala 27:13:@159086.4]
  assign io_dram_0_wdata_bits_wstrb_17 = Fringe_io_dram_0_wdata_bits_wstrb_17; // @[SimTarget.scala 27:13:@159087.4]
  assign io_dram_0_wdata_bits_wstrb_18 = Fringe_io_dram_0_wdata_bits_wstrb_18; // @[SimTarget.scala 27:13:@159088.4]
  assign io_dram_0_wdata_bits_wstrb_19 = Fringe_io_dram_0_wdata_bits_wstrb_19; // @[SimTarget.scala 27:13:@159089.4]
  assign io_dram_0_wdata_bits_wstrb_20 = Fringe_io_dram_0_wdata_bits_wstrb_20; // @[SimTarget.scala 27:13:@159090.4]
  assign io_dram_0_wdata_bits_wstrb_21 = Fringe_io_dram_0_wdata_bits_wstrb_21; // @[SimTarget.scala 27:13:@159091.4]
  assign io_dram_0_wdata_bits_wstrb_22 = Fringe_io_dram_0_wdata_bits_wstrb_22; // @[SimTarget.scala 27:13:@159092.4]
  assign io_dram_0_wdata_bits_wstrb_23 = Fringe_io_dram_0_wdata_bits_wstrb_23; // @[SimTarget.scala 27:13:@159093.4]
  assign io_dram_0_wdata_bits_wstrb_24 = Fringe_io_dram_0_wdata_bits_wstrb_24; // @[SimTarget.scala 27:13:@159094.4]
  assign io_dram_0_wdata_bits_wstrb_25 = Fringe_io_dram_0_wdata_bits_wstrb_25; // @[SimTarget.scala 27:13:@159095.4]
  assign io_dram_0_wdata_bits_wstrb_26 = Fringe_io_dram_0_wdata_bits_wstrb_26; // @[SimTarget.scala 27:13:@159096.4]
  assign io_dram_0_wdata_bits_wstrb_27 = Fringe_io_dram_0_wdata_bits_wstrb_27; // @[SimTarget.scala 27:13:@159097.4]
  assign io_dram_0_wdata_bits_wstrb_28 = Fringe_io_dram_0_wdata_bits_wstrb_28; // @[SimTarget.scala 27:13:@159098.4]
  assign io_dram_0_wdata_bits_wstrb_29 = Fringe_io_dram_0_wdata_bits_wstrb_29; // @[SimTarget.scala 27:13:@159099.4]
  assign io_dram_0_wdata_bits_wstrb_30 = Fringe_io_dram_0_wdata_bits_wstrb_30; // @[SimTarget.scala 27:13:@159100.4]
  assign io_dram_0_wdata_bits_wstrb_31 = Fringe_io_dram_0_wdata_bits_wstrb_31; // @[SimTarget.scala 27:13:@159101.4]
  assign io_dram_0_wdata_bits_wstrb_32 = Fringe_io_dram_0_wdata_bits_wstrb_32; // @[SimTarget.scala 27:13:@159102.4]
  assign io_dram_0_wdata_bits_wstrb_33 = Fringe_io_dram_0_wdata_bits_wstrb_33; // @[SimTarget.scala 27:13:@159103.4]
  assign io_dram_0_wdata_bits_wstrb_34 = Fringe_io_dram_0_wdata_bits_wstrb_34; // @[SimTarget.scala 27:13:@159104.4]
  assign io_dram_0_wdata_bits_wstrb_35 = Fringe_io_dram_0_wdata_bits_wstrb_35; // @[SimTarget.scala 27:13:@159105.4]
  assign io_dram_0_wdata_bits_wstrb_36 = Fringe_io_dram_0_wdata_bits_wstrb_36; // @[SimTarget.scala 27:13:@159106.4]
  assign io_dram_0_wdata_bits_wstrb_37 = Fringe_io_dram_0_wdata_bits_wstrb_37; // @[SimTarget.scala 27:13:@159107.4]
  assign io_dram_0_wdata_bits_wstrb_38 = Fringe_io_dram_0_wdata_bits_wstrb_38; // @[SimTarget.scala 27:13:@159108.4]
  assign io_dram_0_wdata_bits_wstrb_39 = Fringe_io_dram_0_wdata_bits_wstrb_39; // @[SimTarget.scala 27:13:@159109.4]
  assign io_dram_0_wdata_bits_wstrb_40 = Fringe_io_dram_0_wdata_bits_wstrb_40; // @[SimTarget.scala 27:13:@159110.4]
  assign io_dram_0_wdata_bits_wstrb_41 = Fringe_io_dram_0_wdata_bits_wstrb_41; // @[SimTarget.scala 27:13:@159111.4]
  assign io_dram_0_wdata_bits_wstrb_42 = Fringe_io_dram_0_wdata_bits_wstrb_42; // @[SimTarget.scala 27:13:@159112.4]
  assign io_dram_0_wdata_bits_wstrb_43 = Fringe_io_dram_0_wdata_bits_wstrb_43; // @[SimTarget.scala 27:13:@159113.4]
  assign io_dram_0_wdata_bits_wstrb_44 = Fringe_io_dram_0_wdata_bits_wstrb_44; // @[SimTarget.scala 27:13:@159114.4]
  assign io_dram_0_wdata_bits_wstrb_45 = Fringe_io_dram_0_wdata_bits_wstrb_45; // @[SimTarget.scala 27:13:@159115.4]
  assign io_dram_0_wdata_bits_wstrb_46 = Fringe_io_dram_0_wdata_bits_wstrb_46; // @[SimTarget.scala 27:13:@159116.4]
  assign io_dram_0_wdata_bits_wstrb_47 = Fringe_io_dram_0_wdata_bits_wstrb_47; // @[SimTarget.scala 27:13:@159117.4]
  assign io_dram_0_wdata_bits_wstrb_48 = Fringe_io_dram_0_wdata_bits_wstrb_48; // @[SimTarget.scala 27:13:@159118.4]
  assign io_dram_0_wdata_bits_wstrb_49 = Fringe_io_dram_0_wdata_bits_wstrb_49; // @[SimTarget.scala 27:13:@159119.4]
  assign io_dram_0_wdata_bits_wstrb_50 = Fringe_io_dram_0_wdata_bits_wstrb_50; // @[SimTarget.scala 27:13:@159120.4]
  assign io_dram_0_wdata_bits_wstrb_51 = Fringe_io_dram_0_wdata_bits_wstrb_51; // @[SimTarget.scala 27:13:@159121.4]
  assign io_dram_0_wdata_bits_wstrb_52 = Fringe_io_dram_0_wdata_bits_wstrb_52; // @[SimTarget.scala 27:13:@159122.4]
  assign io_dram_0_wdata_bits_wstrb_53 = Fringe_io_dram_0_wdata_bits_wstrb_53; // @[SimTarget.scala 27:13:@159123.4]
  assign io_dram_0_wdata_bits_wstrb_54 = Fringe_io_dram_0_wdata_bits_wstrb_54; // @[SimTarget.scala 27:13:@159124.4]
  assign io_dram_0_wdata_bits_wstrb_55 = Fringe_io_dram_0_wdata_bits_wstrb_55; // @[SimTarget.scala 27:13:@159125.4]
  assign io_dram_0_wdata_bits_wstrb_56 = Fringe_io_dram_0_wdata_bits_wstrb_56; // @[SimTarget.scala 27:13:@159126.4]
  assign io_dram_0_wdata_bits_wstrb_57 = Fringe_io_dram_0_wdata_bits_wstrb_57; // @[SimTarget.scala 27:13:@159127.4]
  assign io_dram_0_wdata_bits_wstrb_58 = Fringe_io_dram_0_wdata_bits_wstrb_58; // @[SimTarget.scala 27:13:@159128.4]
  assign io_dram_0_wdata_bits_wstrb_59 = Fringe_io_dram_0_wdata_bits_wstrb_59; // @[SimTarget.scala 27:13:@159129.4]
  assign io_dram_0_wdata_bits_wstrb_60 = Fringe_io_dram_0_wdata_bits_wstrb_60; // @[SimTarget.scala 27:13:@159130.4]
  assign io_dram_0_wdata_bits_wstrb_61 = Fringe_io_dram_0_wdata_bits_wstrb_61; // @[SimTarget.scala 27:13:@159131.4]
  assign io_dram_0_wdata_bits_wstrb_62 = Fringe_io_dram_0_wdata_bits_wstrb_62; // @[SimTarget.scala 27:13:@159132.4]
  assign io_dram_0_wdata_bits_wstrb_63 = Fringe_io_dram_0_wdata_bits_wstrb_63; // @[SimTarget.scala 27:13:@159133.4]
  assign io_dram_0_wdata_bits_wlast = Fringe_io_dram_0_wdata_bits_wlast; // @[SimTarget.scala 27:13:@159069.4]
  assign io_dram_0_rresp_ready = Fringe_io_dram_0_rresp_ready; // @[SimTarget.scala 27:13:@159068.4]
  assign io_dram_0_wresp_ready = Fringe_io_dram_0_wresp_ready; // @[SimTarget.scala 27:13:@159001.4]
  assign accel_clock = clock; // @[:@157689.4]
  assign accel_reset = reset; // @[:@157690.4]
  assign accel_io_enable = Fringe_io_enable; // @[SimTarget.scala 45:21:@159738.4]
  assign accel_io_reset = Fringe_io_reset; // @[SimTarget.scala 47:20:@159740.4]
  assign accel_io_memStreams_loads_0_cmd_ready = Fringe_io_memStreams_loads_0_cmd_ready; // @[SimTarget.scala 43:26:@159731.4]
  assign accel_io_memStreams_loads_0_data_valid = Fringe_io_memStreams_loads_0_data_valid; // @[SimTarget.scala 43:26:@159726.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = Fringe_io_memStreams_loads_0_data_bits_rdata_0; // @[SimTarget.scala 43:26:@159725.4]
  assign accel_io_memStreams_stores_0_cmd_ready = Fringe_io_memStreams_stores_0_cmd_ready; // @[SimTarget.scala 43:26:@159724.4]
  assign accel_io_memStreams_stores_0_data_ready = Fringe_io_memStreams_stores_0_data_ready; // @[SimTarget.scala 43:26:@159720.4]
  assign accel_io_memStreams_stores_0_wresp_valid = Fringe_io_memStreams_stores_0_wresp_valid; // @[SimTarget.scala 43:26:@159715.4]
  assign accel_io_memStreams_stores_0_wresp_bits = Fringe_io_memStreams_stores_0_wresp_bits; // @[SimTarget.scala 43:26:@159714.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[SimTarget.scala 43:26:@159713.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[SimTarget.scala 43:26:@159646.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 8'h0; // @[SimTarget.scala 43:26:@159582.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 8'h0; // @[SimTarget.scala 43:26:@159583.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 8'h0; // @[SimTarget.scala 43:26:@159584.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 8'h0; // @[SimTarget.scala 43:26:@159585.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 8'h0; // @[SimTarget.scala 43:26:@159586.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 8'h0; // @[SimTarget.scala 43:26:@159587.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 8'h0; // @[SimTarget.scala 43:26:@159588.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 8'h0; // @[SimTarget.scala 43:26:@159589.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 8'h0; // @[SimTarget.scala 43:26:@159590.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 8'h0; // @[SimTarget.scala 43:26:@159591.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 8'h0; // @[SimTarget.scala 43:26:@159592.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 8'h0; // @[SimTarget.scala 43:26:@159593.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 8'h0; // @[SimTarget.scala 43:26:@159594.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 8'h0; // @[SimTarget.scala 43:26:@159595.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 8'h0; // @[SimTarget.scala 43:26:@159596.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 8'h0; // @[SimTarget.scala 43:26:@159597.4]
  assign accel_io_memStreams_gathers_0_data_bits_16 = 8'h0; // @[SimTarget.scala 43:26:@159598.4]
  assign accel_io_memStreams_gathers_0_data_bits_17 = 8'h0; // @[SimTarget.scala 43:26:@159599.4]
  assign accel_io_memStreams_gathers_0_data_bits_18 = 8'h0; // @[SimTarget.scala 43:26:@159600.4]
  assign accel_io_memStreams_gathers_0_data_bits_19 = 8'h0; // @[SimTarget.scala 43:26:@159601.4]
  assign accel_io_memStreams_gathers_0_data_bits_20 = 8'h0; // @[SimTarget.scala 43:26:@159602.4]
  assign accel_io_memStreams_gathers_0_data_bits_21 = 8'h0; // @[SimTarget.scala 43:26:@159603.4]
  assign accel_io_memStreams_gathers_0_data_bits_22 = 8'h0; // @[SimTarget.scala 43:26:@159604.4]
  assign accel_io_memStreams_gathers_0_data_bits_23 = 8'h0; // @[SimTarget.scala 43:26:@159605.4]
  assign accel_io_memStreams_gathers_0_data_bits_24 = 8'h0; // @[SimTarget.scala 43:26:@159606.4]
  assign accel_io_memStreams_gathers_0_data_bits_25 = 8'h0; // @[SimTarget.scala 43:26:@159607.4]
  assign accel_io_memStreams_gathers_0_data_bits_26 = 8'h0; // @[SimTarget.scala 43:26:@159608.4]
  assign accel_io_memStreams_gathers_0_data_bits_27 = 8'h0; // @[SimTarget.scala 43:26:@159609.4]
  assign accel_io_memStreams_gathers_0_data_bits_28 = 8'h0; // @[SimTarget.scala 43:26:@159610.4]
  assign accel_io_memStreams_gathers_0_data_bits_29 = 8'h0; // @[SimTarget.scala 43:26:@159611.4]
  assign accel_io_memStreams_gathers_0_data_bits_30 = 8'h0; // @[SimTarget.scala 43:26:@159612.4]
  assign accel_io_memStreams_gathers_0_data_bits_31 = 8'h0; // @[SimTarget.scala 43:26:@159613.4]
  assign accel_io_memStreams_gathers_0_data_bits_32 = 8'h0; // @[SimTarget.scala 43:26:@159614.4]
  assign accel_io_memStreams_gathers_0_data_bits_33 = 8'h0; // @[SimTarget.scala 43:26:@159615.4]
  assign accel_io_memStreams_gathers_0_data_bits_34 = 8'h0; // @[SimTarget.scala 43:26:@159616.4]
  assign accel_io_memStreams_gathers_0_data_bits_35 = 8'h0; // @[SimTarget.scala 43:26:@159617.4]
  assign accel_io_memStreams_gathers_0_data_bits_36 = 8'h0; // @[SimTarget.scala 43:26:@159618.4]
  assign accel_io_memStreams_gathers_0_data_bits_37 = 8'h0; // @[SimTarget.scala 43:26:@159619.4]
  assign accel_io_memStreams_gathers_0_data_bits_38 = 8'h0; // @[SimTarget.scala 43:26:@159620.4]
  assign accel_io_memStreams_gathers_0_data_bits_39 = 8'h0; // @[SimTarget.scala 43:26:@159621.4]
  assign accel_io_memStreams_gathers_0_data_bits_40 = 8'h0; // @[SimTarget.scala 43:26:@159622.4]
  assign accel_io_memStreams_gathers_0_data_bits_41 = 8'h0; // @[SimTarget.scala 43:26:@159623.4]
  assign accel_io_memStreams_gathers_0_data_bits_42 = 8'h0; // @[SimTarget.scala 43:26:@159624.4]
  assign accel_io_memStreams_gathers_0_data_bits_43 = 8'h0; // @[SimTarget.scala 43:26:@159625.4]
  assign accel_io_memStreams_gathers_0_data_bits_44 = 8'h0; // @[SimTarget.scala 43:26:@159626.4]
  assign accel_io_memStreams_gathers_0_data_bits_45 = 8'h0; // @[SimTarget.scala 43:26:@159627.4]
  assign accel_io_memStreams_gathers_0_data_bits_46 = 8'h0; // @[SimTarget.scala 43:26:@159628.4]
  assign accel_io_memStreams_gathers_0_data_bits_47 = 8'h0; // @[SimTarget.scala 43:26:@159629.4]
  assign accel_io_memStreams_gathers_0_data_bits_48 = 8'h0; // @[SimTarget.scala 43:26:@159630.4]
  assign accel_io_memStreams_gathers_0_data_bits_49 = 8'h0; // @[SimTarget.scala 43:26:@159631.4]
  assign accel_io_memStreams_gathers_0_data_bits_50 = 8'h0; // @[SimTarget.scala 43:26:@159632.4]
  assign accel_io_memStreams_gathers_0_data_bits_51 = 8'h0; // @[SimTarget.scala 43:26:@159633.4]
  assign accel_io_memStreams_gathers_0_data_bits_52 = 8'h0; // @[SimTarget.scala 43:26:@159634.4]
  assign accel_io_memStreams_gathers_0_data_bits_53 = 8'h0; // @[SimTarget.scala 43:26:@159635.4]
  assign accel_io_memStreams_gathers_0_data_bits_54 = 8'h0; // @[SimTarget.scala 43:26:@159636.4]
  assign accel_io_memStreams_gathers_0_data_bits_55 = 8'h0; // @[SimTarget.scala 43:26:@159637.4]
  assign accel_io_memStreams_gathers_0_data_bits_56 = 8'h0; // @[SimTarget.scala 43:26:@159638.4]
  assign accel_io_memStreams_gathers_0_data_bits_57 = 8'h0; // @[SimTarget.scala 43:26:@159639.4]
  assign accel_io_memStreams_gathers_0_data_bits_58 = 8'h0; // @[SimTarget.scala 43:26:@159640.4]
  assign accel_io_memStreams_gathers_0_data_bits_59 = 8'h0; // @[SimTarget.scala 43:26:@159641.4]
  assign accel_io_memStreams_gathers_0_data_bits_60 = 8'h0; // @[SimTarget.scala 43:26:@159642.4]
  assign accel_io_memStreams_gathers_0_data_bits_61 = 8'h0; // @[SimTarget.scala 43:26:@159643.4]
  assign accel_io_memStreams_gathers_0_data_bits_62 = 8'h0; // @[SimTarget.scala 43:26:@159644.4]
  assign accel_io_memStreams_gathers_0_data_bits_63 = 8'h0; // @[SimTarget.scala 43:26:@159645.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[SimTarget.scala 43:26:@159581.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[SimTarget.scala 43:26:@159450.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[SimTarget.scala 43:26:@159449.4]
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = Fringe_io_heap_0_resp_valid; // @[SimTarget.scala 44:20:@159734.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = Fringe_io_heap_0_resp_bits_allocDealloc; // @[SimTarget.scala 44:20:@159733.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = Fringe_io_heap_0_resp_bits_sizeAddr; // @[SimTarget.scala 44:20:@159732.4]
  assign accel_io_argIns_0 = Fringe_io_argIns_0; // @[SimTarget.scala 30:23:@159207.4]
  assign accel_io_argIns_1 = Fringe_io_argIns_1; // @[SimTarget.scala 30:23:@159208.4]
  assign accel_io_argOuts_0_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159211.4]
  assign accel_io_argOuts_0_echo = Fringe_io_argEchos_0; // @[SimTarget.scala 40:26:@159389.4]
  assign accel_io_argOuts_1_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159214.4]
  assign accel_io_argOuts_1_echo = Fringe_io_argEchos_1; // @[SimTarget.scala 40:26:@159390.4]
  assign accel_io_argOuts_2_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159217.4]
  assign accel_io_argOuts_2_echo = Fringe_io_argEchos_2; // @[SimTarget.scala 40:26:@159391.4]
  assign accel_io_argOuts_3_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159220.4]
  assign accel_io_argOuts_3_echo = Fringe_io_argEchos_3; // @[SimTarget.scala 40:26:@159392.4]
  assign accel_io_argOuts_4_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159223.4]
  assign accel_io_argOuts_4_echo = Fringe_io_argEchos_4; // @[SimTarget.scala 40:26:@159393.4]
  assign accel_io_argOuts_5_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159226.4]
  assign accel_io_argOuts_5_echo = Fringe_io_argEchos_5; // @[SimTarget.scala 40:26:@159394.4]
  assign accel_io_argOuts_6_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159229.4]
  assign accel_io_argOuts_6_echo = Fringe_io_argEchos_6; // @[SimTarget.scala 40:26:@159395.4]
  assign accel_io_argOuts_7_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159232.4]
  assign accel_io_argOuts_7_echo = Fringe_io_argEchos_7; // @[SimTarget.scala 40:26:@159396.4]
  assign accel_io_argOuts_8_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159235.4]
  assign accel_io_argOuts_8_echo = Fringe_io_argEchos_8; // @[SimTarget.scala 40:26:@159397.4]
  assign accel_io_argOuts_9_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159238.4]
  assign accel_io_argOuts_9_echo = Fringe_io_argEchos_9; // @[SimTarget.scala 40:26:@159398.4]
  assign accel_io_argOuts_10_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159241.4]
  assign accel_io_argOuts_10_echo = Fringe_io_argEchos_10; // @[SimTarget.scala 40:26:@159399.4]
  assign accel_io_argOuts_11_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159244.4]
  assign accel_io_argOuts_11_echo = Fringe_io_argEchos_11; // @[SimTarget.scala 40:26:@159400.4]
  assign accel_io_argOuts_12_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159247.4]
  assign accel_io_argOuts_12_echo = Fringe_io_argEchos_12; // @[SimTarget.scala 40:26:@159401.4]
  assign accel_io_argOuts_13_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159250.4]
  assign accel_io_argOuts_13_echo = Fringe_io_argEchos_13; // @[SimTarget.scala 40:26:@159402.4]
  assign accel_io_argOuts_14_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159253.4]
  assign accel_io_argOuts_14_echo = Fringe_io_argEchos_14; // @[SimTarget.scala 40:26:@159403.4]
  assign accel_io_argOuts_15_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159256.4]
  assign accel_io_argOuts_15_echo = Fringe_io_argEchos_15; // @[SimTarget.scala 40:26:@159404.4]
  assign accel_io_argOuts_16_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159259.4]
  assign accel_io_argOuts_16_echo = Fringe_io_argEchos_16; // @[SimTarget.scala 40:26:@159405.4]
  assign accel_io_argOuts_17_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159262.4]
  assign accel_io_argOuts_17_echo = Fringe_io_argEchos_17; // @[SimTarget.scala 40:26:@159406.4]
  assign accel_io_argOuts_18_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159265.4]
  assign accel_io_argOuts_18_echo = Fringe_io_argEchos_18; // @[SimTarget.scala 40:26:@159407.4]
  assign accel_io_argOuts_19_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159268.4]
  assign accel_io_argOuts_19_echo = Fringe_io_argEchos_19; // @[SimTarget.scala 40:26:@159408.4]
  assign accel_io_argOuts_20_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159271.4]
  assign accel_io_argOuts_20_echo = Fringe_io_argEchos_20; // @[SimTarget.scala 40:26:@159409.4]
  assign accel_io_argOuts_21_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159274.4]
  assign accel_io_argOuts_21_echo = Fringe_io_argEchos_21; // @[SimTarget.scala 40:26:@159410.4]
  assign accel_io_argOuts_22_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159277.4]
  assign accel_io_argOuts_22_echo = Fringe_io_argEchos_22; // @[SimTarget.scala 40:26:@159411.4]
  assign accel_io_argOuts_23_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159280.4]
  assign accel_io_argOuts_23_echo = Fringe_io_argEchos_23; // @[SimTarget.scala 40:26:@159412.4]
  assign accel_io_argOuts_24_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159283.4]
  assign accel_io_argOuts_24_echo = Fringe_io_argEchos_24; // @[SimTarget.scala 40:26:@159413.4]
  assign accel_io_argOuts_25_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159286.4]
  assign accel_io_argOuts_25_echo = Fringe_io_argEchos_25; // @[SimTarget.scala 40:26:@159414.4]
  assign accel_io_argOuts_26_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159289.4]
  assign accel_io_argOuts_26_echo = Fringe_io_argEchos_26; // @[SimTarget.scala 40:26:@159415.4]
  assign accel_io_argOuts_27_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159292.4]
  assign accel_io_argOuts_27_echo = Fringe_io_argEchos_27; // @[SimTarget.scala 40:26:@159416.4]
  assign accel_io_argOuts_28_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159295.4]
  assign accel_io_argOuts_28_echo = Fringe_io_argEchos_28; // @[SimTarget.scala 40:26:@159417.4]
  assign accel_io_argOuts_29_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159298.4]
  assign accel_io_argOuts_29_echo = Fringe_io_argEchos_29; // @[SimTarget.scala 40:26:@159418.4]
  assign accel_io_argOuts_30_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159301.4]
  assign accel_io_argOuts_30_echo = Fringe_io_argEchos_30; // @[SimTarget.scala 40:26:@159419.4]
  assign accel_io_argOuts_31_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159304.4]
  assign accel_io_argOuts_31_echo = Fringe_io_argEchos_31; // @[SimTarget.scala 40:26:@159420.4]
  assign accel_io_argOuts_32_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159307.4]
  assign accel_io_argOuts_32_echo = Fringe_io_argEchos_32; // @[SimTarget.scala 40:26:@159421.4]
  assign accel_io_argOuts_33_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159310.4]
  assign accel_io_argOuts_33_echo = Fringe_io_argEchos_33; // @[SimTarget.scala 40:26:@159422.4]
  assign accel_io_argOuts_34_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159313.4]
  assign accel_io_argOuts_34_echo = Fringe_io_argEchos_34; // @[SimTarget.scala 40:26:@159423.4]
  assign accel_io_argOuts_35_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159316.4]
  assign accel_io_argOuts_35_echo = Fringe_io_argEchos_35; // @[SimTarget.scala 40:26:@159424.4]
  assign accel_io_argOuts_36_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159319.4]
  assign accel_io_argOuts_36_echo = Fringe_io_argEchos_36; // @[SimTarget.scala 40:26:@159425.4]
  assign accel_io_argOuts_37_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159322.4]
  assign accel_io_argOuts_37_echo = Fringe_io_argEchos_37; // @[SimTarget.scala 40:26:@159426.4]
  assign accel_io_argOuts_38_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159325.4]
  assign accel_io_argOuts_38_echo = Fringe_io_argEchos_38; // @[SimTarget.scala 40:26:@159427.4]
  assign accel_io_argOuts_39_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159328.4]
  assign accel_io_argOuts_39_echo = Fringe_io_argEchos_39; // @[SimTarget.scala 40:26:@159428.4]
  assign accel_io_argOuts_40_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159331.4]
  assign accel_io_argOuts_40_echo = Fringe_io_argEchos_40; // @[SimTarget.scala 40:26:@159429.4]
  assign accel_io_argOuts_41_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159334.4]
  assign accel_io_argOuts_41_echo = Fringe_io_argEchos_41; // @[SimTarget.scala 40:26:@159430.4]
  assign accel_io_argOuts_42_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159337.4]
  assign accel_io_argOuts_42_echo = Fringe_io_argEchos_42; // @[SimTarget.scala 40:26:@159431.4]
  assign accel_io_argOuts_43_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159340.4]
  assign accel_io_argOuts_43_echo = Fringe_io_argEchos_43; // @[SimTarget.scala 40:26:@159432.4]
  assign accel_io_argOuts_44_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159343.4]
  assign accel_io_argOuts_44_echo = Fringe_io_argEchos_44; // @[SimTarget.scala 40:26:@159433.4]
  assign accel_io_argOuts_45_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159346.4]
  assign accel_io_argOuts_45_echo = Fringe_io_argEchos_45; // @[SimTarget.scala 40:26:@159434.4]
  assign accel_io_argOuts_46_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159349.4]
  assign accel_io_argOuts_46_echo = Fringe_io_argEchos_46; // @[SimTarget.scala 40:26:@159435.4]
  assign accel_io_argOuts_47_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159352.4]
  assign accel_io_argOuts_47_echo = Fringe_io_argEchos_47; // @[SimTarget.scala 40:26:@159436.4]
  assign accel_io_argOuts_48_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159355.4]
  assign accel_io_argOuts_48_echo = Fringe_io_argEchos_48; // @[SimTarget.scala 40:26:@159437.4]
  assign accel_io_argOuts_49_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159358.4]
  assign accel_io_argOuts_49_echo = Fringe_io_argEchos_49; // @[SimTarget.scala 40:26:@159438.4]
  assign accel_io_argOuts_50_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159361.4]
  assign accel_io_argOuts_50_echo = Fringe_io_argEchos_50; // @[SimTarget.scala 40:26:@159439.4]
  assign accel_io_argOuts_51_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159364.4]
  assign accel_io_argOuts_51_echo = Fringe_io_argEchos_51; // @[SimTarget.scala 40:26:@159440.4]
  assign accel_io_argOuts_52_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159367.4]
  assign accel_io_argOuts_52_echo = Fringe_io_argEchos_52; // @[SimTarget.scala 40:26:@159441.4]
  assign accel_io_argOuts_53_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159370.4]
  assign accel_io_argOuts_53_echo = Fringe_io_argEchos_53; // @[SimTarget.scala 40:26:@159442.4]
  assign accel_io_argOuts_54_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159373.4]
  assign accel_io_argOuts_54_echo = Fringe_io_argEchos_54; // @[SimTarget.scala 40:26:@159443.4]
  assign accel_io_argOuts_55_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159376.4]
  assign accel_io_argOuts_55_echo = Fringe_io_argEchos_55; // @[SimTarget.scala 40:26:@159444.4]
  assign accel_io_argOuts_56_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159379.4]
  assign accel_io_argOuts_56_echo = Fringe_io_argEchos_56; // @[SimTarget.scala 40:26:@159445.4]
  assign accel_io_argOuts_57_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159382.4]
  assign accel_io_argOuts_57_echo = Fringe_io_argEchos_57; // @[SimTarget.scala 40:26:@159446.4]
  assign accel_io_argOuts_58_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159385.4]
  assign accel_io_argOuts_58_echo = Fringe_io_argEchos_58; // @[SimTarget.scala 40:26:@159447.4]
  assign accel_io_argOuts_59_port_ready = 1'h1; // @[SimTarget.scala 37:32:@159388.4]
  assign accel_io_argOuts_59_echo = Fringe_io_argEchos_59; // @[SimTarget.scala 40:26:@159448.4]
  assign Fringe_clock = clock; // @[:@158244.4]
  assign Fringe_reset = reset; // @[:@158245.4]
  assign Fringe_io_raddr = io_raddr; // @[SimTarget.scala 20:21:@158994.4]
  assign Fringe_io_wen = io_wen; // @[SimTarget.scala 21:21:@158995.4]
  assign Fringe_io_waddr = io_waddr; // @[SimTarget.scala 22:21:@158996.4]
  assign Fringe_io_wdata = io_wdata; // @[SimTarget.scala 23:21:@158997.4]
  assign Fringe_io_done = accel_io_done; // @[SimTarget.scala 46:20:@159739.4]
  assign Fringe_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[SimTarget.scala 36:28:@159210.4]
  assign Fringe_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[SimTarget.scala 35:27:@159209.4]
  assign Fringe_io_argOuts_1_valid = accel_io_argOuts_1_port_valid; // @[SimTarget.scala 36:28:@159213.4]
  assign Fringe_io_argOuts_1_bits = accel_io_argOuts_1_port_bits; // @[SimTarget.scala 35:27:@159212.4]
  assign Fringe_io_argOuts_2_valid = accel_io_argOuts_2_port_valid; // @[SimTarget.scala 36:28:@159216.4]
  assign Fringe_io_argOuts_2_bits = accel_io_argOuts_2_port_bits; // @[SimTarget.scala 35:27:@159215.4]
  assign Fringe_io_argOuts_3_valid = accel_io_argOuts_3_port_valid; // @[SimTarget.scala 36:28:@159219.4]
  assign Fringe_io_argOuts_3_bits = accel_io_argOuts_3_port_bits; // @[SimTarget.scala 35:27:@159218.4]
  assign Fringe_io_argOuts_4_valid = accel_io_argOuts_4_port_valid; // @[SimTarget.scala 36:28:@159222.4]
  assign Fringe_io_argOuts_4_bits = accel_io_argOuts_4_port_bits; // @[SimTarget.scala 35:27:@159221.4]
  assign Fringe_io_argOuts_5_valid = accel_io_argOuts_5_port_valid; // @[SimTarget.scala 36:28:@159225.4]
  assign Fringe_io_argOuts_5_bits = accel_io_argOuts_5_port_bits; // @[SimTarget.scala 35:27:@159224.4]
  assign Fringe_io_argOuts_6_valid = accel_io_argOuts_6_port_valid; // @[SimTarget.scala 36:28:@159228.4]
  assign Fringe_io_argOuts_6_bits = accel_io_argOuts_6_port_bits; // @[SimTarget.scala 35:27:@159227.4]
  assign Fringe_io_argOuts_7_valid = accel_io_argOuts_7_port_valid; // @[SimTarget.scala 36:28:@159231.4]
  assign Fringe_io_argOuts_7_bits = accel_io_argOuts_7_port_bits; // @[SimTarget.scala 35:27:@159230.4]
  assign Fringe_io_argOuts_8_valid = accel_io_argOuts_8_port_valid; // @[SimTarget.scala 36:28:@159234.4]
  assign Fringe_io_argOuts_8_bits = accel_io_argOuts_8_port_bits; // @[SimTarget.scala 35:27:@159233.4]
  assign Fringe_io_argOuts_9_valid = accel_io_argOuts_9_port_valid; // @[SimTarget.scala 36:28:@159237.4]
  assign Fringe_io_argOuts_9_bits = accel_io_argOuts_9_port_bits; // @[SimTarget.scala 35:27:@159236.4]
  assign Fringe_io_argOuts_10_valid = accel_io_argOuts_10_port_valid; // @[SimTarget.scala 36:28:@159240.4]
  assign Fringe_io_argOuts_10_bits = accel_io_argOuts_10_port_bits; // @[SimTarget.scala 35:27:@159239.4]
  assign Fringe_io_argOuts_11_valid = accel_io_argOuts_11_port_valid; // @[SimTarget.scala 36:28:@159243.4]
  assign Fringe_io_argOuts_11_bits = accel_io_argOuts_11_port_bits; // @[SimTarget.scala 35:27:@159242.4]
  assign Fringe_io_argOuts_12_valid = accel_io_argOuts_12_port_valid; // @[SimTarget.scala 36:28:@159246.4]
  assign Fringe_io_argOuts_12_bits = accel_io_argOuts_12_port_bits; // @[SimTarget.scala 35:27:@159245.4]
  assign Fringe_io_argOuts_13_valid = accel_io_argOuts_13_port_valid; // @[SimTarget.scala 36:28:@159249.4]
  assign Fringe_io_argOuts_13_bits = accel_io_argOuts_13_port_bits; // @[SimTarget.scala 35:27:@159248.4]
  assign Fringe_io_argOuts_14_valid = accel_io_argOuts_14_port_valid; // @[SimTarget.scala 36:28:@159252.4]
  assign Fringe_io_argOuts_14_bits = accel_io_argOuts_14_port_bits; // @[SimTarget.scala 35:27:@159251.4]
  assign Fringe_io_argOuts_15_valid = accel_io_argOuts_15_port_valid; // @[SimTarget.scala 36:28:@159255.4]
  assign Fringe_io_argOuts_15_bits = accel_io_argOuts_15_port_bits; // @[SimTarget.scala 35:27:@159254.4]
  assign Fringe_io_argOuts_16_valid = accel_io_argOuts_16_port_valid; // @[SimTarget.scala 36:28:@159258.4]
  assign Fringe_io_argOuts_16_bits = accel_io_argOuts_16_port_bits; // @[SimTarget.scala 35:27:@159257.4]
  assign Fringe_io_argOuts_17_valid = accel_io_argOuts_17_port_valid; // @[SimTarget.scala 36:28:@159261.4]
  assign Fringe_io_argOuts_17_bits = accel_io_argOuts_17_port_bits; // @[SimTarget.scala 35:27:@159260.4]
  assign Fringe_io_argOuts_18_valid = accel_io_argOuts_18_port_valid; // @[SimTarget.scala 36:28:@159264.4]
  assign Fringe_io_argOuts_18_bits = accel_io_argOuts_18_port_bits; // @[SimTarget.scala 35:27:@159263.4]
  assign Fringe_io_argOuts_19_valid = accel_io_argOuts_19_port_valid; // @[SimTarget.scala 36:28:@159267.4]
  assign Fringe_io_argOuts_19_bits = accel_io_argOuts_19_port_bits; // @[SimTarget.scala 35:27:@159266.4]
  assign Fringe_io_argOuts_20_valid = accel_io_argOuts_20_port_valid; // @[SimTarget.scala 36:28:@159270.4]
  assign Fringe_io_argOuts_20_bits = accel_io_argOuts_20_port_bits; // @[SimTarget.scala 35:27:@159269.4]
  assign Fringe_io_argOuts_21_valid = accel_io_argOuts_21_port_valid; // @[SimTarget.scala 36:28:@159273.4]
  assign Fringe_io_argOuts_21_bits = accel_io_argOuts_21_port_bits; // @[SimTarget.scala 35:27:@159272.4]
  assign Fringe_io_argOuts_22_valid = accel_io_argOuts_22_port_valid; // @[SimTarget.scala 36:28:@159276.4]
  assign Fringe_io_argOuts_22_bits = accel_io_argOuts_22_port_bits; // @[SimTarget.scala 35:27:@159275.4]
  assign Fringe_io_argOuts_23_valid = accel_io_argOuts_23_port_valid; // @[SimTarget.scala 36:28:@159279.4]
  assign Fringe_io_argOuts_23_bits = accel_io_argOuts_23_port_bits; // @[SimTarget.scala 35:27:@159278.4]
  assign Fringe_io_argOuts_24_valid = accel_io_argOuts_24_port_valid; // @[SimTarget.scala 36:28:@159282.4]
  assign Fringe_io_argOuts_24_bits = accel_io_argOuts_24_port_bits; // @[SimTarget.scala 35:27:@159281.4]
  assign Fringe_io_argOuts_25_valid = accel_io_argOuts_25_port_valid; // @[SimTarget.scala 36:28:@159285.4]
  assign Fringe_io_argOuts_25_bits = accel_io_argOuts_25_port_bits; // @[SimTarget.scala 35:27:@159284.4]
  assign Fringe_io_argOuts_26_valid = accel_io_argOuts_26_port_valid; // @[SimTarget.scala 36:28:@159288.4]
  assign Fringe_io_argOuts_26_bits = accel_io_argOuts_26_port_bits; // @[SimTarget.scala 35:27:@159287.4]
  assign Fringe_io_argOuts_27_valid = accel_io_argOuts_27_port_valid; // @[SimTarget.scala 36:28:@159291.4]
  assign Fringe_io_argOuts_27_bits = accel_io_argOuts_27_port_bits; // @[SimTarget.scala 35:27:@159290.4]
  assign Fringe_io_argOuts_28_valid = accel_io_argOuts_28_port_valid; // @[SimTarget.scala 36:28:@159294.4]
  assign Fringe_io_argOuts_28_bits = accel_io_argOuts_28_port_bits; // @[SimTarget.scala 35:27:@159293.4]
  assign Fringe_io_argOuts_29_valid = accel_io_argOuts_29_port_valid; // @[SimTarget.scala 36:28:@159297.4]
  assign Fringe_io_argOuts_29_bits = accel_io_argOuts_29_port_bits; // @[SimTarget.scala 35:27:@159296.4]
  assign Fringe_io_argOuts_30_valid = accel_io_argOuts_30_port_valid; // @[SimTarget.scala 36:28:@159300.4]
  assign Fringe_io_argOuts_30_bits = accel_io_argOuts_30_port_bits; // @[SimTarget.scala 35:27:@159299.4]
  assign Fringe_io_argOuts_31_valid = accel_io_argOuts_31_port_valid; // @[SimTarget.scala 36:28:@159303.4]
  assign Fringe_io_argOuts_31_bits = accel_io_argOuts_31_port_bits; // @[SimTarget.scala 35:27:@159302.4]
  assign Fringe_io_argOuts_32_valid = accel_io_argOuts_32_port_valid; // @[SimTarget.scala 36:28:@159306.4]
  assign Fringe_io_argOuts_32_bits = accel_io_argOuts_32_port_bits; // @[SimTarget.scala 35:27:@159305.4]
  assign Fringe_io_argOuts_33_valid = accel_io_argOuts_33_port_valid; // @[SimTarget.scala 36:28:@159309.4]
  assign Fringe_io_argOuts_33_bits = accel_io_argOuts_33_port_bits; // @[SimTarget.scala 35:27:@159308.4]
  assign Fringe_io_argOuts_34_valid = accel_io_argOuts_34_port_valid; // @[SimTarget.scala 36:28:@159312.4]
  assign Fringe_io_argOuts_34_bits = accel_io_argOuts_34_port_bits; // @[SimTarget.scala 35:27:@159311.4]
  assign Fringe_io_argOuts_35_valid = accel_io_argOuts_35_port_valid; // @[SimTarget.scala 36:28:@159315.4]
  assign Fringe_io_argOuts_35_bits = accel_io_argOuts_35_port_bits; // @[SimTarget.scala 35:27:@159314.4]
  assign Fringe_io_argOuts_36_valid = accel_io_argOuts_36_port_valid; // @[SimTarget.scala 36:28:@159318.4]
  assign Fringe_io_argOuts_36_bits = accel_io_argOuts_36_port_bits; // @[SimTarget.scala 35:27:@159317.4]
  assign Fringe_io_argOuts_37_valid = accel_io_argOuts_37_port_valid; // @[SimTarget.scala 36:28:@159321.4]
  assign Fringe_io_argOuts_37_bits = accel_io_argOuts_37_port_bits; // @[SimTarget.scala 35:27:@159320.4]
  assign Fringe_io_argOuts_38_valid = accel_io_argOuts_38_port_valid; // @[SimTarget.scala 36:28:@159324.4]
  assign Fringe_io_argOuts_38_bits = accel_io_argOuts_38_port_bits; // @[SimTarget.scala 35:27:@159323.4]
  assign Fringe_io_argOuts_39_valid = accel_io_argOuts_39_port_valid; // @[SimTarget.scala 36:28:@159327.4]
  assign Fringe_io_argOuts_39_bits = accel_io_argOuts_39_port_bits; // @[SimTarget.scala 35:27:@159326.4]
  assign Fringe_io_argOuts_40_valid = accel_io_argOuts_40_port_valid; // @[SimTarget.scala 36:28:@159330.4]
  assign Fringe_io_argOuts_40_bits = accel_io_argOuts_40_port_bits; // @[SimTarget.scala 35:27:@159329.4]
  assign Fringe_io_argOuts_41_valid = accel_io_argOuts_41_port_valid; // @[SimTarget.scala 36:28:@159333.4]
  assign Fringe_io_argOuts_41_bits = accel_io_argOuts_41_port_bits; // @[SimTarget.scala 35:27:@159332.4]
  assign Fringe_io_argOuts_42_valid = accel_io_argOuts_42_port_valid; // @[SimTarget.scala 36:28:@159336.4]
  assign Fringe_io_argOuts_42_bits = accel_io_argOuts_42_port_bits; // @[SimTarget.scala 35:27:@159335.4]
  assign Fringe_io_argOuts_43_valid = accel_io_argOuts_43_port_valid; // @[SimTarget.scala 36:28:@159339.4]
  assign Fringe_io_argOuts_43_bits = accel_io_argOuts_43_port_bits; // @[SimTarget.scala 35:27:@159338.4]
  assign Fringe_io_argOuts_44_valid = accel_io_argOuts_44_port_valid; // @[SimTarget.scala 36:28:@159342.4]
  assign Fringe_io_argOuts_44_bits = accel_io_argOuts_44_port_bits; // @[SimTarget.scala 35:27:@159341.4]
  assign Fringe_io_argOuts_45_valid = accel_io_argOuts_45_port_valid; // @[SimTarget.scala 36:28:@159345.4]
  assign Fringe_io_argOuts_45_bits = accel_io_argOuts_45_port_bits; // @[SimTarget.scala 35:27:@159344.4]
  assign Fringe_io_argOuts_46_valid = accel_io_argOuts_46_port_valid; // @[SimTarget.scala 36:28:@159348.4]
  assign Fringe_io_argOuts_46_bits = accel_io_argOuts_46_port_bits; // @[SimTarget.scala 35:27:@159347.4]
  assign Fringe_io_argOuts_47_valid = accel_io_argOuts_47_port_valid; // @[SimTarget.scala 36:28:@159351.4]
  assign Fringe_io_argOuts_47_bits = accel_io_argOuts_47_port_bits; // @[SimTarget.scala 35:27:@159350.4]
  assign Fringe_io_argOuts_48_valid = accel_io_argOuts_48_port_valid; // @[SimTarget.scala 36:28:@159354.4]
  assign Fringe_io_argOuts_48_bits = accel_io_argOuts_48_port_bits; // @[SimTarget.scala 35:27:@159353.4]
  assign Fringe_io_argOuts_49_valid = accel_io_argOuts_49_port_valid; // @[SimTarget.scala 36:28:@159357.4]
  assign Fringe_io_argOuts_49_bits = accel_io_argOuts_49_port_bits; // @[SimTarget.scala 35:27:@159356.4]
  assign Fringe_io_argOuts_50_valid = accel_io_argOuts_50_port_valid; // @[SimTarget.scala 36:28:@159360.4]
  assign Fringe_io_argOuts_50_bits = accel_io_argOuts_50_port_bits; // @[SimTarget.scala 35:27:@159359.4]
  assign Fringe_io_argOuts_51_valid = accel_io_argOuts_51_port_valid; // @[SimTarget.scala 36:28:@159363.4]
  assign Fringe_io_argOuts_51_bits = accel_io_argOuts_51_port_bits; // @[SimTarget.scala 35:27:@159362.4]
  assign Fringe_io_argOuts_52_valid = accel_io_argOuts_52_port_valid; // @[SimTarget.scala 36:28:@159366.4]
  assign Fringe_io_argOuts_52_bits = accel_io_argOuts_52_port_bits; // @[SimTarget.scala 35:27:@159365.4]
  assign Fringe_io_argOuts_53_valid = accel_io_argOuts_53_port_valid; // @[SimTarget.scala 36:28:@159369.4]
  assign Fringe_io_argOuts_53_bits = accel_io_argOuts_53_port_bits; // @[SimTarget.scala 35:27:@159368.4]
  assign Fringe_io_argOuts_54_valid = accel_io_argOuts_54_port_valid; // @[SimTarget.scala 36:28:@159372.4]
  assign Fringe_io_argOuts_54_bits = accel_io_argOuts_54_port_bits; // @[SimTarget.scala 35:27:@159371.4]
  assign Fringe_io_argOuts_55_valid = accel_io_argOuts_55_port_valid; // @[SimTarget.scala 36:28:@159375.4]
  assign Fringe_io_argOuts_55_bits = accel_io_argOuts_55_port_bits; // @[SimTarget.scala 35:27:@159374.4]
  assign Fringe_io_argOuts_56_valid = accel_io_argOuts_56_port_valid; // @[SimTarget.scala 36:28:@159378.4]
  assign Fringe_io_argOuts_56_bits = accel_io_argOuts_56_port_bits; // @[SimTarget.scala 35:27:@159377.4]
  assign Fringe_io_argOuts_57_valid = accel_io_argOuts_57_port_valid; // @[SimTarget.scala 36:28:@159381.4]
  assign Fringe_io_argOuts_57_bits = accel_io_argOuts_57_port_bits; // @[SimTarget.scala 35:27:@159380.4]
  assign Fringe_io_argOuts_58_valid = accel_io_argOuts_58_port_valid; // @[SimTarget.scala 36:28:@159384.4]
  assign Fringe_io_argOuts_58_bits = accel_io_argOuts_58_port_bits; // @[SimTarget.scala 35:27:@159383.4]
  assign Fringe_io_argOuts_59_valid = accel_io_argOuts_59_port_valid; // @[SimTarget.scala 36:28:@159387.4]
  assign Fringe_io_argOuts_59_bits = accel_io_argOuts_59_port_bits; // @[SimTarget.scala 35:27:@159386.4]
  assign Fringe_io_memStreams_loads_0_cmd_valid = accel_io_memStreams_loads_0_cmd_valid; // @[SimTarget.scala 43:26:@159730.4]
  assign Fringe_io_memStreams_loads_0_cmd_bits_addr = accel_io_memStreams_loads_0_cmd_bits_addr; // @[SimTarget.scala 43:26:@159729.4]
  assign Fringe_io_memStreams_loads_0_cmd_bits_size = accel_io_memStreams_loads_0_cmd_bits_size; // @[SimTarget.scala 43:26:@159728.4]
  assign Fringe_io_memStreams_loads_0_data_ready = accel_io_memStreams_loads_0_data_ready; // @[SimTarget.scala 43:26:@159727.4]
  assign Fringe_io_memStreams_stores_0_cmd_valid = accel_io_memStreams_stores_0_cmd_valid; // @[SimTarget.scala 43:26:@159723.4]
  assign Fringe_io_memStreams_stores_0_cmd_bits_addr = accel_io_memStreams_stores_0_cmd_bits_addr; // @[SimTarget.scala 43:26:@159722.4]
  assign Fringe_io_memStreams_stores_0_cmd_bits_size = accel_io_memStreams_stores_0_cmd_bits_size; // @[SimTarget.scala 43:26:@159721.4]
  assign Fringe_io_memStreams_stores_0_data_valid = accel_io_memStreams_stores_0_data_valid; // @[SimTarget.scala 43:26:@159719.4]
  assign Fringe_io_memStreams_stores_0_data_bits_wdata_0 = accel_io_memStreams_stores_0_data_bits_wdata_0; // @[SimTarget.scala 43:26:@159718.4]
  assign Fringe_io_memStreams_stores_0_data_bits_wstrb = accel_io_memStreams_stores_0_data_bits_wstrb; // @[SimTarget.scala 43:26:@159717.4]
  assign Fringe_io_memStreams_stores_0_wresp_ready = accel_io_memStreams_stores_0_wresp_ready; // @[SimTarget.scala 43:26:@159716.4]
  assign Fringe_io_dram_0_cmd_ready = io_dram_0_cmd_ready; // @[SimTarget.scala 27:13:@159206.4]
  assign Fringe_io_dram_0_wdata_ready = io_dram_0_wdata_ready; // @[SimTarget.scala 27:13:@159199.4]
  assign Fringe_io_dram_0_rresp_valid = io_dram_0_rresp_valid; // @[SimTarget.scala 27:13:@159067.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_0 = io_dram_0_rresp_bits_rdata_0; // @[SimTarget.scala 27:13:@159003.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_1 = io_dram_0_rresp_bits_rdata_1; // @[SimTarget.scala 27:13:@159004.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_2 = io_dram_0_rresp_bits_rdata_2; // @[SimTarget.scala 27:13:@159005.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_3 = io_dram_0_rresp_bits_rdata_3; // @[SimTarget.scala 27:13:@159006.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_4 = io_dram_0_rresp_bits_rdata_4; // @[SimTarget.scala 27:13:@159007.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_5 = io_dram_0_rresp_bits_rdata_5; // @[SimTarget.scala 27:13:@159008.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_6 = io_dram_0_rresp_bits_rdata_6; // @[SimTarget.scala 27:13:@159009.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_7 = io_dram_0_rresp_bits_rdata_7; // @[SimTarget.scala 27:13:@159010.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_8 = io_dram_0_rresp_bits_rdata_8; // @[SimTarget.scala 27:13:@159011.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_9 = io_dram_0_rresp_bits_rdata_9; // @[SimTarget.scala 27:13:@159012.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_10 = io_dram_0_rresp_bits_rdata_10; // @[SimTarget.scala 27:13:@159013.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_11 = io_dram_0_rresp_bits_rdata_11; // @[SimTarget.scala 27:13:@159014.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_12 = io_dram_0_rresp_bits_rdata_12; // @[SimTarget.scala 27:13:@159015.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_13 = io_dram_0_rresp_bits_rdata_13; // @[SimTarget.scala 27:13:@159016.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_14 = io_dram_0_rresp_bits_rdata_14; // @[SimTarget.scala 27:13:@159017.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_15 = io_dram_0_rresp_bits_rdata_15; // @[SimTarget.scala 27:13:@159018.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_16 = io_dram_0_rresp_bits_rdata_16; // @[SimTarget.scala 27:13:@159019.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_17 = io_dram_0_rresp_bits_rdata_17; // @[SimTarget.scala 27:13:@159020.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_18 = io_dram_0_rresp_bits_rdata_18; // @[SimTarget.scala 27:13:@159021.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_19 = io_dram_0_rresp_bits_rdata_19; // @[SimTarget.scala 27:13:@159022.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_20 = io_dram_0_rresp_bits_rdata_20; // @[SimTarget.scala 27:13:@159023.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_21 = io_dram_0_rresp_bits_rdata_21; // @[SimTarget.scala 27:13:@159024.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_22 = io_dram_0_rresp_bits_rdata_22; // @[SimTarget.scala 27:13:@159025.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_23 = io_dram_0_rresp_bits_rdata_23; // @[SimTarget.scala 27:13:@159026.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_24 = io_dram_0_rresp_bits_rdata_24; // @[SimTarget.scala 27:13:@159027.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_25 = io_dram_0_rresp_bits_rdata_25; // @[SimTarget.scala 27:13:@159028.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_26 = io_dram_0_rresp_bits_rdata_26; // @[SimTarget.scala 27:13:@159029.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_27 = io_dram_0_rresp_bits_rdata_27; // @[SimTarget.scala 27:13:@159030.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_28 = io_dram_0_rresp_bits_rdata_28; // @[SimTarget.scala 27:13:@159031.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_29 = io_dram_0_rresp_bits_rdata_29; // @[SimTarget.scala 27:13:@159032.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_30 = io_dram_0_rresp_bits_rdata_30; // @[SimTarget.scala 27:13:@159033.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_31 = io_dram_0_rresp_bits_rdata_31; // @[SimTarget.scala 27:13:@159034.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_32 = io_dram_0_rresp_bits_rdata_32; // @[SimTarget.scala 27:13:@159035.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_33 = io_dram_0_rresp_bits_rdata_33; // @[SimTarget.scala 27:13:@159036.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_34 = io_dram_0_rresp_bits_rdata_34; // @[SimTarget.scala 27:13:@159037.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_35 = io_dram_0_rresp_bits_rdata_35; // @[SimTarget.scala 27:13:@159038.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_36 = io_dram_0_rresp_bits_rdata_36; // @[SimTarget.scala 27:13:@159039.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_37 = io_dram_0_rresp_bits_rdata_37; // @[SimTarget.scala 27:13:@159040.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_38 = io_dram_0_rresp_bits_rdata_38; // @[SimTarget.scala 27:13:@159041.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_39 = io_dram_0_rresp_bits_rdata_39; // @[SimTarget.scala 27:13:@159042.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_40 = io_dram_0_rresp_bits_rdata_40; // @[SimTarget.scala 27:13:@159043.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_41 = io_dram_0_rresp_bits_rdata_41; // @[SimTarget.scala 27:13:@159044.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_42 = io_dram_0_rresp_bits_rdata_42; // @[SimTarget.scala 27:13:@159045.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_43 = io_dram_0_rresp_bits_rdata_43; // @[SimTarget.scala 27:13:@159046.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_44 = io_dram_0_rresp_bits_rdata_44; // @[SimTarget.scala 27:13:@159047.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_45 = io_dram_0_rresp_bits_rdata_45; // @[SimTarget.scala 27:13:@159048.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_46 = io_dram_0_rresp_bits_rdata_46; // @[SimTarget.scala 27:13:@159049.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_47 = io_dram_0_rresp_bits_rdata_47; // @[SimTarget.scala 27:13:@159050.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_48 = io_dram_0_rresp_bits_rdata_48; // @[SimTarget.scala 27:13:@159051.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_49 = io_dram_0_rresp_bits_rdata_49; // @[SimTarget.scala 27:13:@159052.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_50 = io_dram_0_rresp_bits_rdata_50; // @[SimTarget.scala 27:13:@159053.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_51 = io_dram_0_rresp_bits_rdata_51; // @[SimTarget.scala 27:13:@159054.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_52 = io_dram_0_rresp_bits_rdata_52; // @[SimTarget.scala 27:13:@159055.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_53 = io_dram_0_rresp_bits_rdata_53; // @[SimTarget.scala 27:13:@159056.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_54 = io_dram_0_rresp_bits_rdata_54; // @[SimTarget.scala 27:13:@159057.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_55 = io_dram_0_rresp_bits_rdata_55; // @[SimTarget.scala 27:13:@159058.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_56 = io_dram_0_rresp_bits_rdata_56; // @[SimTarget.scala 27:13:@159059.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_57 = io_dram_0_rresp_bits_rdata_57; // @[SimTarget.scala 27:13:@159060.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_58 = io_dram_0_rresp_bits_rdata_58; // @[SimTarget.scala 27:13:@159061.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_59 = io_dram_0_rresp_bits_rdata_59; // @[SimTarget.scala 27:13:@159062.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_60 = io_dram_0_rresp_bits_rdata_60; // @[SimTarget.scala 27:13:@159063.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_61 = io_dram_0_rresp_bits_rdata_61; // @[SimTarget.scala 27:13:@159064.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_62 = io_dram_0_rresp_bits_rdata_62; // @[SimTarget.scala 27:13:@159065.4]
  assign Fringe_io_dram_0_rresp_bits_rdata_63 = io_dram_0_rresp_bits_rdata_63; // @[SimTarget.scala 27:13:@159066.4]
  assign Fringe_io_dram_0_rresp_bits_tag = io_dram_0_rresp_bits_tag; // @[SimTarget.scala 27:13:@159002.4]
  assign Fringe_io_dram_0_wresp_valid = io_dram_0_wresp_valid; // @[SimTarget.scala 27:13:@159000.4]
  assign Fringe_io_dram_0_wresp_bits_tag = io_dram_0_wresp_bits_tag; // @[SimTarget.scala 27:13:@158999.4]
  assign Fringe_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[SimTarget.scala 44:20:@159737.4]
  assign Fringe_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[SimTarget.scala 44:20:@159736.4]
  assign Fringe_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[SimTarget.scala 44:20:@159735.4]
endmodule
