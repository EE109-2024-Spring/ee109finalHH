module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 325:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 325:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 325:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 262:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 262:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 262:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 262:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 262:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 262:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 264:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 264:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 264:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 264:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 264:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 264:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 288:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 292:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 292:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 292:33:@104.4]
  wire  _T_57; // @[Counter.scala 294:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 300:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 300:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 300:74:@118.4]
  FF bases_0 ( // @[Counter.scala 262:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 264:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 288:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 292:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 292:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 292:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh50); // @[Counter.scala 294:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 300:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 300:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 300:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh50); // @[Counter.scala 334:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 300:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 282:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 285:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 265:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 266:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 267:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@390.2]
  input   clock, // @[:@391.4]
  input   reset, // @[:@392.4]
  input   io_enable, // @[:@393.4]
  output  io_done, // @[:@393.4]
  input   io_rst, // @[:@393.4]
  input   io_ctrDone, // @[:@393.4]
  output  io_ctrInc, // @[:@393.4]
  input   io_doneIn_0, // @[:@393.4]
  input   io_doneIn_1, // @[:@393.4]
  input   io_doneIn_2, // @[:@393.4]
  output  io_enableOut_0, // @[:@393.4]
  output  io_enableOut_1, // @[:@393.4]
  output  io_enableOut_2, // @[:@393.4]
  output  io_childAck_0, // @[:@393.4]
  output  io_childAck_1, // @[:@393.4]
  output  io_childAck_2 // @[:@393.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@396.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@396.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@396.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@396.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@396.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@396.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@399.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@399.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@399.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@399.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@399.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@399.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@402.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@402.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@402.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@402.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@402.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@402.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@405.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@405.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@405.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@405.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@405.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@405.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@408.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@408.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@408.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@408.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@408.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@408.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@411.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@411.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@411.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@411.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@411.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@411.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@452.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@452.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@452.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@452.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@452.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@452.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@455.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@455.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@455.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@455.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@455.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@455.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@458.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@458.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@458.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@458.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@458.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@458.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@497.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@497.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@497.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@497.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@497.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@630.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@630.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@630.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@630.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@630.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@647.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@647.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@647.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@647.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@647.4]
  wire  _T_77; // @[Controllers.scala 80:47:@414.4]
  wire  allDone; // @[Controllers.scala 80:47:@415.4]
  wire  _T_78; // @[Controllers.scala 81:26:@416.4]
  wire  finished; // @[Controllers.scala 81:37:@417.4]
  wire  synchronize; // @[package.scala 96:25:@502.4 package.scala 96:25:@503.4]
  wire  _T_168; // @[Controllers.scala 128:33:@511.4]
  wire  _T_170; // @[Controllers.scala 128:54:@512.4]
  wire  _T_171; // @[Controllers.scala 128:52:@513.4]
  wire  _T_172; // @[Controllers.scala 128:66:@514.4]
  wire  _T_174; // @[Controllers.scala 128:98:@516.4]
  wire  _T_175; // @[Controllers.scala 128:96:@517.4]
  wire  _T_177; // @[Controllers.scala 128:123:@518.4]
  wire  _T_179; // @[Controllers.scala 129:48:@521.4]
  wire  _T_184; // @[Controllers.scala 130:52:@526.4]
  wire  _T_185; // @[Controllers.scala 130:50:@527.4]
  wire  _T_193; // @[Controllers.scala 130:129:@533.4]
  wire  _T_196; // @[Controllers.scala 131:45:@536.4]
  wire  _T_199; // @[Controllers.scala 135:80:@540.4]
  wire  _T_200; // @[Controllers.scala 135:78:@541.4]
  wire  _T_202; // @[Controllers.scala 135:105:@542.4]
  wire  _T_203; // @[Controllers.scala 135:103:@543.4]
  wire  _T_204; // @[Controllers.scala 135:119:@544.4]
  wire  _T_206; // @[Controllers.scala 135:51:@546.4]
  wire  _T_227; // @[Controllers.scala 135:80:@567.4]
  wire  _T_228; // @[Controllers.scala 135:78:@568.4]
  wire  _T_230; // @[Controllers.scala 135:105:@569.4]
  wire  _T_231; // @[Controllers.scala 135:103:@570.4]
  wire  _T_232; // @[Controllers.scala 135:119:@571.4]
  wire  _T_234; // @[Controllers.scala 135:51:@573.4]
  wire  _T_258; // @[Controllers.scala 213:68:@600.4]
  wire  _T_260; // @[Controllers.scala 213:90:@602.4]
  wire  _T_262; // @[Controllers.scala 213:132:@604.4]
  wire  _T_263; // @[Controllers.scala 213:130:@605.4]
  wire  _T_264; // @[Controllers.scala 213:156:@606.4]
  wire  _T_266; // @[Controllers.scala 213:68:@609.4]
  wire  _T_268; // @[Controllers.scala 213:90:@611.4]
  wire  _T_274; // @[Controllers.scala 213:68:@617.4]
  wire  _T_276; // @[Controllers.scala 213:90:@619.4]
  wire  _T_283; // @[package.scala 100:49:@625.4]
  reg  _T_286; // @[package.scala 48:56:@626.4]
  reg [31:0] _RAND_0;
  reg  _T_300; // @[package.scala 48:56:@644.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@396.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@399.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@402.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@405.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@408.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@411.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@452.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@455.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@458.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@497.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@630.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@647.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@414.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@415.4]
  assign _T_78 = allDone | io_done; // @[Controllers.scala 81:26:@416.4]
  assign finished = _T_78 | done_2_io_input_set; // @[Controllers.scala 81:37:@417.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@502.4 package.scala 96:25:@503.4]
  assign _T_168 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@511.4]
  assign _T_170 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@512.4]
  assign _T_171 = _T_168 & _T_170; // @[Controllers.scala 128:52:@513.4]
  assign _T_172 = _T_171 & io_enable; // @[Controllers.scala 128:66:@514.4]
  assign _T_174 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@516.4]
  assign _T_175 = _T_172 & _T_174; // @[Controllers.scala 128:96:@517.4]
  assign _T_177 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@518.4]
  assign _T_179 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@521.4]
  assign _T_184 = synchronize == 1'h0; // @[Controllers.scala 130:52:@526.4]
  assign _T_185 = io_doneIn_0 & _T_184; // @[Controllers.scala 130:50:@527.4]
  assign _T_193 = finished == 1'h0; // @[Controllers.scala 130:129:@533.4]
  assign _T_196 = io_rst == 1'h0; // @[Controllers.scala 131:45:@536.4]
  assign _T_199 = ~ iterDone_1_io_output; // @[Controllers.scala 135:80:@540.4]
  assign _T_200 = iterDone_0_io_output & _T_199; // @[Controllers.scala 135:78:@541.4]
  assign _T_202 = io_doneIn_1 == 1'h0; // @[Controllers.scala 135:105:@542.4]
  assign _T_203 = _T_200 & _T_202; // @[Controllers.scala 135:103:@543.4]
  assign _T_204 = _T_203 & io_enable; // @[Controllers.scala 135:119:@544.4]
  assign _T_206 = io_doneIn_0 | _T_204; // @[Controllers.scala 135:51:@546.4]
  assign _T_227 = ~ iterDone_2_io_output; // @[Controllers.scala 135:80:@567.4]
  assign _T_228 = iterDone_1_io_output & _T_227; // @[Controllers.scala 135:78:@568.4]
  assign _T_230 = io_doneIn_2 == 1'h0; // @[Controllers.scala 135:105:@569.4]
  assign _T_231 = _T_228 & _T_230; // @[Controllers.scala 135:103:@570.4]
  assign _T_232 = _T_231 & io_enable; // @[Controllers.scala 135:119:@571.4]
  assign _T_234 = io_doneIn_1 | _T_232; // @[Controllers.scala 135:51:@573.4]
  assign _T_258 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@600.4]
  assign _T_260 = _T_258 & _T_174; // @[Controllers.scala 213:90:@602.4]
  assign _T_262 = ~ allDone; // @[Controllers.scala 213:132:@604.4]
  assign _T_263 = _T_260 & _T_262; // @[Controllers.scala 213:130:@605.4]
  assign _T_264 = ~ io_ctrDone; // @[Controllers.scala 213:156:@606.4]
  assign _T_266 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@609.4]
  assign _T_268 = _T_266 & _T_199; // @[Controllers.scala 213:90:@611.4]
  assign _T_274 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@617.4]
  assign _T_276 = _T_274 & _T_227; // @[Controllers.scala 213:90:@619.4]
  assign _T_283 = allDone == 1'h0; // @[package.scala 100:49:@625.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@654.4]
  assign io_ctrInc = io_doneIn_2; // @[Controllers.scala 122:17:@496.4]
  assign io_enableOut_0 = _T_263 & _T_264; // @[Controllers.scala 213:55:@608.4]
  assign io_enableOut_1 = _T_268 & _T_262; // @[Controllers.scala 213:55:@616.4]
  assign io_enableOut_2 = _T_276 & _T_262; // @[Controllers.scala 213:55:@624.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@595.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@597.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@599.4]
  assign active_0_clock = clock; // @[:@397.4]
  assign active_0_reset = reset; // @[:@398.4]
  assign active_0_io_input_set = _T_175 & _T_177; // @[Controllers.scala 128:30:@520.4]
  assign active_0_io_input_reset = _T_179 | allDone; // @[Controllers.scala 129:32:@525.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@418.4]
  assign active_1_clock = clock; // @[:@400.4]
  assign active_1_reset = reset; // @[:@401.4]
  assign active_1_io_input_set = _T_206 & _T_184; // @[Controllers.scala 135:32:@549.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_rst; // @[Controllers.scala 136:34:@553.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@419.4]
  assign active_2_clock = clock; // @[:@403.4]
  assign active_2_reset = reset; // @[:@404.4]
  assign active_2_io_input_set = _T_234 & _T_184; // @[Controllers.scala 135:32:@576.4]
  assign active_2_io_input_reset = io_doneIn_2 | io_rst; // @[Controllers.scala 136:34:@580.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@420.4]
  assign done_0_clock = clock; // @[:@406.4]
  assign done_0_reset = reset; // @[:@407.4]
  assign done_0_io_input_set = io_ctrDone & _T_196; // @[Controllers.scala 131:28:@539.4]
  assign done_0_io_input_reset = io_rst | allDone; // @[Controllers.scala 86:33:@432.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@421.4]
  assign done_1_clock = clock; // @[:@409.4]
  assign done_1_reset = reset; // @[:@410.4]
  assign done_1_io_input_set = io_ctrDone & _T_196; // @[Controllers.scala 138:30:@566.4]
  assign done_1_io_input_reset = io_rst | allDone; // @[Controllers.scala 86:33:@441.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@422.4]
  assign done_2_clock = clock; // @[:@412.4]
  assign done_2_reset = reset; // @[:@413.4]
  assign done_2_io_input_set = io_ctrDone & _T_196; // @[Controllers.scala 138:30:@593.4]
  assign done_2_io_input_reset = io_rst | allDone; // @[Controllers.scala 86:33:@450.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@423.4]
  assign iterDone_0_clock = clock; // @[:@453.4]
  assign iterDone_0_reset = reset; // @[:@454.4]
  assign iterDone_0_io_input_set = _T_185 & _T_193; // @[Controllers.scala 130:32:@535.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@472.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@461.4]
  assign iterDone_1_clock = clock; // @[:@456.4]
  assign iterDone_1_reset = reset; // @[:@457.4]
  assign iterDone_1_io_input_set = io_doneIn_1 & _T_184; // @[Controllers.scala 137:34:@562.4]
  assign iterDone_1_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@481.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@462.4]
  assign iterDone_2_clock = clock; // @[:@459.4]
  assign iterDone_2_reset = reset; // @[:@460.4]
  assign iterDone_2_io_input_set = io_doneIn_2 & _T_184; // @[Controllers.scala 137:34:@589.4]
  assign iterDone_2_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@490.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@463.4]
  assign RetimeWrapper_clock = clock; // @[:@498.4]
  assign RetimeWrapper_reset = reset; // @[:@499.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@501.4]
  assign RetimeWrapper_io_in = io_doneIn_2; // @[package.scala 94:16:@500.4]
  assign RetimeWrapper_1_clock = clock; // @[:@631.4]
  assign RetimeWrapper_1_reset = reset; // @[:@632.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@634.4]
  assign RetimeWrapper_1_io_in = allDone & _T_286; // @[package.scala 94:16:@633.4]
  assign RetimeWrapper_2_clock = clock; // @[:@648.4]
  assign RetimeWrapper_2_reset = reset; // @[:@649.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@651.4]
  assign RetimeWrapper_2_io_in = allDone & _T_300; // @[package.scala 94:16:@650.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_286 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_300 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_286 <= 1'h0;
    end else begin
      _T_286 <= _T_283;
    end
    if (reset) begin
      _T_300 <= 1'h0;
    end else begin
      _T_300 <= _T_283;
    end
  end
endmodule
module SRAM( // @[:@721.2]
  input         clock, // @[:@722.4]
  input         reset, // @[:@723.4]
  input  [8:0]  io_raddr, // @[:@724.4]
  input         io_wen, // @[:@724.4]
  input  [8:0]  io_waddr, // @[:@724.4]
  input  [31:0] io_wdata, // @[:@724.4]
  output [31:0] io_rdata, // @[:@724.4]
  input         io_backpressure // @[:@724.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@726.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@726.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@726.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@726.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@726.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@726.4]
  wire [8:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@726.4]
  wire [8:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@726.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@726.4]
  wire  _T_19; // @[SRAM.scala 182:49:@744.4]
  wire  _T_20; // @[SRAM.scala 182:37:@745.4]
  reg  _T_23; // @[SRAM.scala 182:29:@746.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@748.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(300), .AWIDTH(9)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@726.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@744.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@745.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@753.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@740.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@741.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@738.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@743.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@742.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@739.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@737.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@736.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_5( // @[:@767.2]
  input        clock, // @[:@768.4]
  input        reset, // @[:@769.4]
  input        io_flow, // @[:@770.4]
  input  [8:0] io_in, // @[:@770.4]
  output [8:0] io_out // @[:@770.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@772.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@772.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@772.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@772.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@772.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@772.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@772.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@785.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@784.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@783.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@782.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@781.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@779.4]
endmodule
module Mem1D( // @[:@787.2]
  input         clock, // @[:@788.4]
  input         reset, // @[:@789.4]
  input  [8:0]  io_r_ofs_0, // @[:@790.4]
  input         io_r_backpressure, // @[:@790.4]
  input  [8:0]  io_w_ofs_0, // @[:@790.4]
  input  [31:0] io_w_data_0, // @[:@790.4]
  input         io_w_en_0, // @[:@790.4]
  output [31:0] io_output // @[:@790.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 753:21:@794.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 753:21:@794.4]
  wire [8:0] SRAM_io_raddr; // @[MemPrimitives.scala 753:21:@794.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 753:21:@794.4]
  wire [8:0] SRAM_io_waddr; // @[MemPrimitives.scala 753:21:@794.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 753:21:@794.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 753:21:@794.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 753:21:@794.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@797.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@797.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@797.4]
  wire [8:0] RetimeWrapper_io_in; // @[package.scala 93:22:@797.4]
  wire [8:0] RetimeWrapper_io_out; // @[package.scala 93:22:@797.4]
  wire  wInBound; // @[MemPrimitives.scala 740:32:@792.4]
  SRAM SRAM ( // @[MemPrimitives.scala 753:21:@794.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@797.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 9'h12c; // @[MemPrimitives.scala 740:32:@792.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 760:17:@810.4]
  assign SRAM_clock = clock; // @[:@795.4]
  assign SRAM_reset = reset; // @[:@796.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 754:37:@804.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 757:22:@807.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 756:22:@805.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 758:22:@808.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 759:30:@809.4]
  assign RetimeWrapper_clock = clock; // @[:@798.4]
  assign RetimeWrapper_reset = reset; // @[:@799.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@801.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@800.4]
endmodule
module StickySelects( // @[:@812.2]
  input   io_ins_0, // @[:@815.4]
  output  io_outs_0 // @[:@815.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@817.4]
endmodule
module RetimeWrapper_6( // @[:@831.2]
  input   clock, // @[:@832.4]
  input   reset, // @[:@833.4]
  input   io_flow, // @[:@834.4]
  input   io_in, // @[:@834.4]
  output  io_out // @[:@834.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@836.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@836.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@836.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@836.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@836.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@836.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@836.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@849.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@848.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@847.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@846.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@845.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@843.4]
endmodule
module x471_A_sram_0( // @[:@851.2]
  input         clock, // @[:@852.4]
  input         reset, // @[:@853.4]
  input  [8:0]  io_rPort_0_ofs_0, // @[:@854.4]
  input         io_rPort_0_en_0, // @[:@854.4]
  input         io_rPort_0_backpressure, // @[:@854.4]
  output [31:0] io_rPort_0_output_0, // @[:@854.4]
  input  [8:0]  io_wPort_0_ofs_0, // @[:@854.4]
  input  [31:0] io_wPort_0_data_0, // @[:@854.4]
  input         io_wPort_0_en_0 // @[:@854.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@869.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@869.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@869.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@869.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@869.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@869.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@869.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@869.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@895.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@895.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@909.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@909.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@909.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@909.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@909.4]
  wire [41:0] _T_70; // @[Cat.scala 30:58:@887.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@899.4]
  wire [10:0] _T_78; // @[Cat.scala 30:58:@901.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@869.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@895.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@909.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_70 = {io_wPort_0_en_0,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@887.4]
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@899.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@901.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@916.4]
  assign Mem1D_clock = clock; // @[:@870.4]
  assign Mem1D_reset = reset; // @[:@871.4]
  assign Mem1D_io_r_ofs_0 = _T_78[8:0]; // @[MemPrimitives.scala 131:28:@905.4]
  assign Mem1D_io_r_backpressure = _T_78[9]; // @[MemPrimitives.scala 132:32:@906.4]
  assign Mem1D_io_w_ofs_0 = _T_70[8:0]; // @[MemPrimitives.scala 94:28:@891.4]
  assign Mem1D_io_w_data_0 = _T_70[40:9]; // @[MemPrimitives.scala 95:29:@892.4]
  assign Mem1D_io_w_en_0 = _T_70[41]; // @[MemPrimitives.scala 96:27:@893.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@898.4]
  assign RetimeWrapper_clock = clock; // @[:@910.4]
  assign RetimeWrapper_reset = reset; // @[:@911.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@913.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@912.4]
endmodule
module x538_outr_UnitPipe_DenseTransfer_sm( // @[:@1678.2]
  input   clock, // @[:@1679.4]
  input   reset, // @[:@1680.4]
  input   io_enable, // @[:@1681.4]
  output  io_done, // @[:@1681.4]
  input   io_parentAck, // @[:@1681.4]
  input   io_doneIn_0, // @[:@1681.4]
  input   io_doneIn_1, // @[:@1681.4]
  output  io_enableOut_0, // @[:@1681.4]
  output  io_enableOut_1, // @[:@1681.4]
  output  io_childAck_0, // @[:@1681.4]
  output  io_childAck_1, // @[:@1681.4]
  input   io_ctrCopyDone_0, // @[:@1681.4]
  input   io_ctrCopyDone_1 // @[:@1681.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1684.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1684.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1684.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1684.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1684.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1684.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1687.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1687.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1687.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1687.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1687.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1687.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1690.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1690.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1690.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1690.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1690.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1690.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1693.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1693.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1693.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1693.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1693.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1693.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1722.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1722.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1722.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1722.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1722.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1722.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1725.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1725.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1725.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1725.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1725.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1725.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1766.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1766.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1766.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1766.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1766.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1780.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1780.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1780.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1780.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1780.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1798.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1798.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1798.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1798.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1798.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1835.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1835.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1835.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1835.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1835.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1849.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1849.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1849.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1849.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1849.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1867.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1867.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1867.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1867.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1867.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1914.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1914.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1914.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1914.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1914.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1931.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1931.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1931.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1931.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1931.4]
  wire  allDone; // @[Controllers.scala 80:47:@1696.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1750.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1751.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1752.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1753.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1754.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1757.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1759.4]
  wire  _T_148; // @[package.scala 96:25:@1771.4 package.scala 96:25:@1772.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1774.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1775.4]
  wire  _T_160; // @[package.scala 96:25:@1785.4 package.scala 96:25:@1786.4]
  wire  _T_178; // @[package.scala 96:25:@1803.4 package.scala 96:25:@1804.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1806.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1807.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1819.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1820.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1821.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1822.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1823.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1826.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1828.4]
  wire  _T_216; // @[package.scala 96:25:@1840.4 package.scala 96:25:@1841.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1843.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1844.4]
  wire  _T_228; // @[package.scala 96:25:@1854.4 package.scala 96:25:@1855.4]
  wire  _T_246; // @[package.scala 96:25:@1872.4 package.scala 96:25:@1873.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1875.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1876.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1892.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1894.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1896.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1901.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1903.4]
  wire  _T_282; // @[package.scala 100:49:@1909.4]
  reg  _T_285; // @[package.scala 48:56:@1910.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1912.4]
  reg  _T_299; // @[package.scala 48:56:@1928.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1684.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1687.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1690.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1693.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1722.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1725.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1766.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1780.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1798.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1835.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1849.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1867.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1914.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1931.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1696.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1750.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1751.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1752.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1753.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1754.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1757.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1759.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1771.4 package.scala 96:25:@1772.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1774.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1775.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1785.4 package.scala 96:25:@1786.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1803.4 package.scala 96:25:@1804.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1806.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1807.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1819.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1820.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1821.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1822.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1823.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1826.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1828.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1840.4 package.scala 96:25:@1841.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1843.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1844.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1854.4 package.scala 96:25:@1855.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1872.4 package.scala 96:25:@1873.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1875.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1876.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1892.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1894.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1896.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1901.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1903.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1909.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1912.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1938.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1900.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1908.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1889.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1891.4]
  assign active_0_clock = clock; // @[:@1685.4]
  assign active_0_reset = reset; // @[:@1686.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1761.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1765.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1699.4]
  assign active_1_clock = clock; // @[:@1688.4]
  assign active_1_reset = reset; // @[:@1689.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1830.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1834.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1700.4]
  assign done_0_clock = clock; // @[:@1691.4]
  assign done_0_reset = reset; // @[:@1692.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1811.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1711.4 Controllers.scala 170:32:@1818.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1701.4]
  assign done_1_clock = clock; // @[:@1694.4]
  assign done_1_reset = reset; // @[:@1695.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1880.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1720.4 Controllers.scala 170:32:@1887.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1702.4]
  assign iterDone_0_clock = clock; // @[:@1723.4]
  assign iterDone_0_reset = reset; // @[:@1724.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1779.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1738.4 Controllers.scala 168:36:@1795.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1728.4]
  assign iterDone_1_clock = clock; // @[:@1726.4]
  assign iterDone_1_reset = reset; // @[:@1727.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1848.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1747.4 Controllers.scala 168:36:@1864.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1729.4]
  assign RetimeWrapper_clock = clock; // @[:@1767.4]
  assign RetimeWrapper_reset = reset; // @[:@1768.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1770.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1769.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1781.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1782.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1784.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1783.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1799.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1800.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1802.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1801.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1836.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1837.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1839.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1838.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1850.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1851.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1853.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1852.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1868.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1869.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1871.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1870.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1915.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1916.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1918.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1917.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1932.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1933.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1935.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1934.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module FF_1( // @[:@2021.2]
  input        clock, // @[:@2022.4]
  input        reset, // @[:@2023.4]
  output [6:0] io_rPort_0_output_0, // @[:@2024.4]
  input  [6:0] io_wPort_0_data_0, // @[:@2024.4]
  input        io_wPort_0_reset, // @[:@2024.4]
  input  [6:0] io_wPort_0_init, // @[:@2024.4]
  input        io_wPort_0_en_0, // @[:@2024.4]
  input        io_reset // @[:@2024.4]
);
  reg [6:0] ff; // @[MemPrimitives.scala 321:19:@2039.4]
  reg [31:0] _RAND_0;
  wire  anyReset; // @[MemPrimitives.scala 322:65:@2040.4]
  wire [6:0] _T_68; // @[MemPrimitives.scala 325:32:@2041.4]
  wire [6:0] _T_69; // @[MemPrimitives.scala 325:12:@2042.4]
  assign anyReset = io_wPort_0_reset | io_reset; // @[MemPrimitives.scala 322:65:@2040.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@2041.4]
  assign _T_69 = anyReset ? io_wPort_0_init : _T_68; // @[MemPrimitives.scala 325:12:@2042.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@2044.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= io_wPort_0_init;
    end else begin
      if (anyReset) begin
        ff <= io_wPort_0_init;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module CompactingCounter( // @[:@2046.2]
  input        clock, // @[:@2047.4]
  input        reset, // @[:@2048.4]
  input        io_input_reset, // @[:@2049.4]
  input        io_input_enables_0, // @[:@2049.4]
  output [6:0] io_output_count // @[:@2049.4]
);
  wire  base_clock; // @[Counter.scala 200:20:@2051.4]
  wire  base_reset; // @[Counter.scala 200:20:@2051.4]
  wire [6:0] base_io_rPort_0_output_0; // @[Counter.scala 200:20:@2051.4]
  wire [6:0] base_io_wPort_0_data_0; // @[Counter.scala 200:20:@2051.4]
  wire  base_io_wPort_0_reset; // @[Counter.scala 200:20:@2051.4]
  wire [6:0] base_io_wPort_0_init; // @[Counter.scala 200:20:@2051.4]
  wire  base_io_wPort_0_en_0; // @[Counter.scala 200:20:@2051.4]
  wire  base_io_reset; // @[Counter.scala 200:20:@2051.4]
  wire [6:0] count; // @[Counter.scala 206:42:@2070.4]
  wire [6:0] num_enabled; // @[Counter.scala 207:56:@2071.4]
  wire [7:0] _T_27; // @[Counter.scala 208:22:@2076.4]
  wire [6:0] _T_28; // @[Counter.scala 208:22:@2077.4]
  wire [6:0] newval; // @[Counter.scala 208:22:@2078.4]
  wire  isMax; // @[Counter.scala 209:40:@2079.4]
  wire [7:0] _T_34; // @[Counter.scala 210:32:@2082.4]
  wire [6:0] _T_35; // @[Counter.scala 210:32:@2083.4]
  wire [6:0] _T_36; // @[Counter.scala 210:32:@2084.4]
  wire [6:0] next; // @[Counter.scala 210:17:@2085.4]
  wire [6:0] _T_38; // @[Counter.scala 211:68:@2086.4]
  FF_1 base ( // @[Counter.scala 200:20:@2051.4]
    .clock(base_clock),
    .reset(base_reset),
    .io_rPort_0_output_0(base_io_rPort_0_output_0),
    .io_wPort_0_data_0(base_io_wPort_0_data_0),
    .io_wPort_0_reset(base_io_wPort_0_reset),
    .io_wPort_0_init(base_io_wPort_0_init),
    .io_wPort_0_en_0(base_io_wPort_0_en_0),
    .io_reset(base_io_reset)
  );
  assign count = $signed(base_io_rPort_0_output_0); // @[Counter.scala 206:42:@2070.4]
  assign num_enabled = io_input_enables_0 ? $signed(7'sh1) : $signed(7'sh0); // @[Counter.scala 207:56:@2071.4]
  assign _T_27 = $signed(count) + $signed(num_enabled); // @[Counter.scala 208:22:@2076.4]
  assign _T_28 = $signed(count) + $signed(num_enabled); // @[Counter.scala 208:22:@2077.4]
  assign newval = $signed(_T_28); // @[Counter.scala 208:22:@2078.4]
  assign isMax = $signed(newval) >= $signed(7'sh10); // @[Counter.scala 209:40:@2079.4]
  assign _T_34 = $signed(newval) - $signed(7'sh10); // @[Counter.scala 210:32:@2082.4]
  assign _T_35 = $signed(newval) - $signed(7'sh10); // @[Counter.scala 210:32:@2083.4]
  assign _T_36 = $signed(_T_35); // @[Counter.scala 210:32:@2084.4]
  assign next = isMax ? $signed(_T_36) : $signed(newval); // @[Counter.scala 210:17:@2085.4]
  assign _T_38 = $unsigned(next); // @[Counter.scala 211:68:@2086.4]
  assign io_output_count = $signed(base_io_rPort_0_output_0); // @[Counter.scala 213:19:@2090.4]
  assign base_clock = clock; // @[:@2052.4]
  assign base_reset = reset; // @[:@2053.4]
  assign base_io_wPort_0_data_0 = io_input_reset ? 7'h0 : _T_38; // @[Counter.scala 211:30:@2088.4]
  assign base_io_wPort_0_reset = io_input_reset; // @[Counter.scala 203:26:@2068.4]
  assign base_io_wPort_0_init = 7'h0; // @[Counter.scala 202:25:@2067.4]
  assign base_io_wPort_0_en_0 = io_input_enables_0; // @[Counter.scala 204:28:@2069.4]
  assign base_io_reset = 1'h0;
endmodule
module CompactingIncDincCtr( // @[:@2167.2]
  input   clock, // @[:@2168.4]
  input   reset, // @[:@2169.4]
  input   io_input_inc_en_0, // @[:@2170.4]
  input   io_input_dinc_en_0, // @[:@2170.4]
  output  io_output_empty, // @[:@2170.4]
  output  io_output_full // @[:@2170.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@2172.4]
  reg [31:0] _RAND_0;
  wire [6:0] numPushed; // @[Counter.scala 172:47:@2173.4]
  wire [6:0] numPopped; // @[Counter.scala 173:48:@2174.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@2175.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@2175.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@2176.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@2177.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@2178.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@2178.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@2179.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@2180.4]
  assign numPushed = io_input_inc_en_0 ? $signed(7'sh1) : $signed(7'sh0); // @[Counter.scala 172:47:@2173.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(7'sh1) : $signed(7'sh0); // @[Counter.scala 173:48:@2174.4]
  assign _GEN_0 = {{25{numPushed[6]}},numPushed}; // @[Counter.scala 174:14:@2175.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@2175.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@2176.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@2177.4]
  assign _GEN_1 = {{25{numPopped[6]}},numPopped}; // @[Counter.scala 174:26:@2178.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@2178.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@2179.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@2180.4]
  assign io_output_empty = $signed(cnt) < $signed(32'sh1); // @[Counter.scala 179:19:@2187.4]
  assign io_output_full = $signed(cnt) > $signed(32'shf); // @[Counter.scala 181:18:@2194.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module Mem1D_3( // @[:@2202.2]
  input         clock, // @[:@2203.4]
  input  [4:0]  io_r_ofs_0, // @[:@2205.4]
  input  [4:0]  io_w_ofs_0, // @[:@2205.4]
  input  [95:0] io_w_data_0, // @[:@2205.4]
  input         io_w_en_0, // @[:@2205.4]
  output [95:0] io_output // @[:@2205.4]
);
  reg [95:0] _T_127 [0:15]; // @[MemPrimitives.scala 771:18:@2209.4]
  reg [95:0] _RAND_0;
  wire [95:0] _T_127__T_132_data; // @[MemPrimitives.scala 771:18:@2209.4]
  wire [3:0] _T_127__T_132_addr; // @[MemPrimitives.scala 771:18:@2209.4]
  wire [95:0] _T_127__T_130_data; // @[MemPrimitives.scala 771:18:@2209.4]
  wire [3:0] _T_127__T_130_addr; // @[MemPrimitives.scala 771:18:@2209.4]
  wire  _T_127__T_130_mask; // @[MemPrimitives.scala 771:18:@2209.4]
  wire  _T_127__T_130_en; // @[MemPrimitives.scala 771:18:@2209.4]
  wire  wInBound; // @[MemPrimitives.scala 740:32:@2207.4]
  assign _T_127__T_132_addr = io_r_ofs_0[3:0];
  assign _T_127__T_132_data = _T_127[_T_127__T_132_addr]; // @[MemPrimitives.scala 771:18:@2209.4]
  assign _T_127__T_130_data = io_w_data_0;
  assign _T_127__T_130_addr = io_w_ofs_0[3:0];
  assign _T_127__T_130_mask = 1'h1;
  assign _T_127__T_130_en = io_w_en_0 & wInBound;
  assign wInBound = io_w_ofs_0 <= 5'h10; // @[MemPrimitives.scala 740:32:@2207.4]
  assign io_output = _T_127__T_132_data; // @[MemPrimitives.scala 773:17:@2218.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {3{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    _T_127[initvar] = _RAND_0[95:0];
  `endif // RANDOMIZE_MEM_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(_T_127__T_130_en & _T_127__T_130_mask) begin
      _T_127[_T_127__T_130_addr] <= _T_127__T_130_data; // @[MemPrimitives.scala 771:18:@2209.4]
    end
  end
endmodule
module Compactor( // @[:@2220.2]
  input  [95:0] io_in_0_data, // @[:@2223.4]
  output [95:0] io_out_0_data // @[:@2223.4]
);
  assign io_out_0_data = io_in_0_data; // @[MemPrimitives.scala 848:22:@2227.4]
endmodule
module CompactingEnqNetwork( // @[:@2231.2]
  input  [6:0]  io_headCnt, // @[:@2234.4]
  input  [95:0] io_in_0_data, // @[:@2234.4]
  input         io_in_0_en, // @[:@2234.4]
  output [95:0] io_out_0_data, // @[:@2234.4]
  output        io_out_0_en // @[:@2234.4]
);
  wire [95:0] compactor_io_in_0_data; // @[MemPrimitives.scala 870:25:@2237.4]
  wire [95:0] compactor_io_out_0_data; // @[MemPrimitives.scala 870:25:@2237.4]
  wire [6:0] numEnabled; // @[MemPrimitives.scala 866:38:@2236.4]
  wire [6:0] _GEN_0; // @[Math.scala 53:59:@2243.4]
  wire [6:0] current_base_bank; // @[Math.scala 53:59:@2243.4]
  wire [6:0] _T_22; // @[MemPrimitives.scala 876:46:@2244.4]
  wire [7:0] _T_23; // @[MemPrimitives.scala 876:33:@2245.4]
  wire [6:0] _T_24; // @[MemPrimitives.scala 876:33:@2246.4]
  wire [6:0] _T_25; // @[MemPrimitives.scala 876:33:@2247.4]
  wire [7:0] _T_27; // @[MemPrimitives.scala 876:53:@2248.4]
  wire [6:0] _T_28; // @[MemPrimitives.scala 876:53:@2249.4]
  wire [6:0] upper; // @[MemPrimitives.scala 876:53:@2250.4]
  wire  _T_30; // @[MemPrimitives.scala 877:34:@2251.4]
  wire [6:0] num_straddling; // @[MemPrimitives.scala 877:27:@2252.4]
  wire [7:0] _T_33; // @[MemPrimitives.scala 878:40:@2254.4]
  wire [6:0] _T_34; // @[MemPrimitives.scala 878:40:@2255.4]
  wire [6:0] num_straight; // @[MemPrimitives.scala 878:40:@2256.4]
  wire  _T_36; // @[MemPrimitives.scala 880:40:@2257.4]
  wire  _T_38; // @[MemPrimitives.scala 880:73:@2258.4]
  wire  _T_44; // @[MemPrimitives.scala 880:109:@2263.4]
  wire  _T_45; // @[MemPrimitives.scala 880:94:@2264.4]
  wire [7:0] _T_53; // @[MemPrimitives.scala 881:72:@2268.4]
  wire [6:0] _T_54; // @[MemPrimitives.scala 881:72:@2269.4]
  wire [6:0] _T_55; // @[MemPrimitives.scala 881:72:@2270.4]
  wire [7:0] _T_57; // @[MemPrimitives.scala 881:101:@2271.4]
  wire [6:0] _T_58; // @[MemPrimitives.scala 881:101:@2272.4]
  wire [6:0] _T_59; // @[MemPrimitives.scala 881:101:@2273.4]
  wire [6:0] _T_60; // @[MemPrimitives.scala 881:27:@2274.4]
  wire [6:0] _T_62; // @[MemPrimitives.scala 885:57:@2275.4]
  wire  _T_64; // @[Mux.scala 46:19:@2276.4]
  Compactor compactor ( // @[MemPrimitives.scala 870:25:@2237.4]
    .io_in_0_data(compactor_io_in_0_data),
    .io_out_0_data(compactor_io_out_0_data)
  );
  assign numEnabled = io_in_0_en ? 7'h1 : 7'h0; // @[MemPrimitives.scala 866:38:@2236.4]
  assign _GEN_0 = $signed(io_headCnt) % $signed(7'sh1); // @[Math.scala 53:59:@2243.4]
  assign current_base_bank = _GEN_0[6:0]; // @[Math.scala 53:59:@2243.4]
  assign _T_22 = $signed(numEnabled); // @[MemPrimitives.scala 876:46:@2244.4]
  assign _T_23 = $signed(current_base_bank) + $signed(_T_22); // @[MemPrimitives.scala 876:33:@2245.4]
  assign _T_24 = $signed(current_base_bank) + $signed(_T_22); // @[MemPrimitives.scala 876:33:@2246.4]
  assign _T_25 = $signed(_T_24); // @[MemPrimitives.scala 876:33:@2247.4]
  assign _T_27 = $signed(_T_25) - $signed(7'sh1); // @[MemPrimitives.scala 876:53:@2248.4]
  assign _T_28 = $signed(_T_25) - $signed(7'sh1); // @[MemPrimitives.scala 876:53:@2249.4]
  assign upper = $signed(_T_28); // @[MemPrimitives.scala 876:53:@2250.4]
  assign _T_30 = $signed(upper) < $signed(7'sh0); // @[MemPrimitives.scala 877:34:@2251.4]
  assign num_straddling = _T_30 ? $signed(7'sh0) : $signed(upper); // @[MemPrimitives.scala 877:27:@2252.4]
  assign _T_33 = $signed(_T_22) - $signed(num_straddling); // @[MemPrimitives.scala 878:40:@2254.4]
  assign _T_34 = $signed(_T_22) - $signed(num_straddling); // @[MemPrimitives.scala 878:40:@2255.4]
  assign num_straight = $signed(_T_34); // @[MemPrimitives.scala 878:40:@2256.4]
  assign _T_36 = $signed(7'sh0) < $signed(num_straddling); // @[MemPrimitives.scala 880:40:@2257.4]
  assign _T_38 = $signed(7'sh0) >= $signed(current_base_bank); // @[MemPrimitives.scala 880:73:@2258.4]
  assign _T_44 = $signed(7'sh0) < $signed(_T_25); // @[MemPrimitives.scala 880:109:@2263.4]
  assign _T_45 = _T_38 & _T_44; // @[MemPrimitives.scala 880:94:@2264.4]
  assign _T_53 = {{1{num_straight[6]}},num_straight}; // @[MemPrimitives.scala 881:72:@2268.4]
  assign _T_54 = _T_53[6:0]; // @[MemPrimitives.scala 881:72:@2269.4]
  assign _T_55 = $signed(_T_54); // @[MemPrimitives.scala 881:72:@2270.4]
  assign _T_57 = $signed(7'sh0) - $signed(current_base_bank); // @[MemPrimitives.scala 881:101:@2271.4]
  assign _T_58 = $signed(7'sh0) - $signed(current_base_bank); // @[MemPrimitives.scala 881:101:@2272.4]
  assign _T_59 = $signed(_T_58); // @[MemPrimitives.scala 881:101:@2273.4]
  assign _T_60 = _T_36 ? $signed(_T_55) : $signed(_T_59); // @[MemPrimitives.scala 881:27:@2274.4]
  assign _T_62 = $unsigned(_T_60); // @[MemPrimitives.scala 885:57:@2275.4]
  assign _T_64 = 7'h0 == _T_62; // @[Mux.scala 46:19:@2276.4]
  assign io_out_0_data = _T_64 ? compactor_io_out_0_data : 96'h0; // @[MemPrimitives.scala 890:63:@2278.4]
  assign io_out_0_en = _T_36 | _T_45; // @[MemPrimitives.scala 891:63:@2279.4]
  assign compactor_io_in_0_data = io_in_0_data; // @[MemPrimitives.scala 871:19:@2241.4]
endmodule
module CompactingDeqNetwork( // @[:@2281.2]
  input  [6:0]  io_tailCnt, // @[:@2284.4]
  input  [95:0] io_input_data_0, // @[:@2284.4]
  output [95:0] io_output_0 // @[:@2284.4]
);
  wire [6:0] _GEN_0; // @[Math.scala 53:59:@2288.4]
  wire [6:0] current_base_bank; // @[Math.scala 53:59:@2288.4]
  wire [6:0] _T_55; // @[MemPrimitives.scala 917:64:@2311.4]
  wire [7:0] _T_56; // @[MemPrimitives.scala 917:71:@2312.4]
  wire [6:0] _T_57; // @[MemPrimitives.scala 917:71:@2313.4]
  wire [6:0] _GEN_1; // @[Math.scala 55:59:@2314.4]
  wire [6:0] _T_59; // @[Math.scala 55:59:@2314.4]
  wire  _T_62; // @[Mux.scala 46:19:@2315.4]
  assign _GEN_0 = $signed(io_tailCnt) % $signed(7'sh1); // @[Math.scala 53:59:@2288.4]
  assign current_base_bank = _GEN_0[6:0]; // @[Math.scala 53:59:@2288.4]
  assign _T_55 = $unsigned(current_base_bank); // @[MemPrimitives.scala 917:64:@2311.4]
  assign _T_56 = {{1'd0}, _T_55}; // @[MemPrimitives.scala 917:71:@2312.4]
  assign _T_57 = _T_56[6:0]; // @[MemPrimitives.scala 917:71:@2313.4]
  assign _GEN_1 = _T_57 % 7'h1; // @[Math.scala 55:59:@2314.4]
  assign _T_59 = _GEN_1[6:0]; // @[Math.scala 55:59:@2314.4]
  assign _T_62 = 7'h0 == _T_59; // @[Mux.scala 46:19:@2315.4]
  assign io_output_0 = _T_62 ? io_input_data_0 : 96'h0; // @[MemPrimitives.scala 921:18:@2317.4]
endmodule
module x475_fifo( // @[:@2319.2]
  input         clock, // @[:@2320.4]
  input         reset, // @[:@2321.4]
  input         io_rPort_0_en_0, // @[:@2322.4]
  output [95:0] io_rPort_0_output_0, // @[:@2322.4]
  input  [95:0] io_wPort_0_data_0, // @[:@2322.4]
  input         io_wPort_0_en_0, // @[:@2322.4]
  output        io_full, // @[:@2322.4]
  output        io_empty, // @[:@2322.4]
  input         io_active_0_in, // @[:@2322.4]
  output        io_active_0_out // @[:@2322.4]
);
  wire  headCtr_clock; // @[MemPrimitives.scala 381:23:@2346.4]
  wire  headCtr_reset; // @[MemPrimitives.scala 381:23:@2346.4]
  wire  headCtr_io_input_reset; // @[MemPrimitives.scala 381:23:@2346.4]
  wire  headCtr_io_input_enables_0; // @[MemPrimitives.scala 381:23:@2346.4]
  wire [6:0] headCtr_io_output_count; // @[MemPrimitives.scala 381:23:@2346.4]
  wire  tailCtr_clock; // @[MemPrimitives.scala 382:23:@2354.4]
  wire  tailCtr_reset; // @[MemPrimitives.scala 382:23:@2354.4]
  wire  tailCtr_io_input_reset; // @[MemPrimitives.scala 382:23:@2354.4]
  wire  tailCtr_io_input_enables_0; // @[MemPrimitives.scala 382:23:@2354.4]
  wire [6:0] tailCtr_io_output_count; // @[MemPrimitives.scala 382:23:@2354.4]
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2368.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2368.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2368.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2368.4]
  wire  elements_io_output_empty; // @[MemPrimitives.scala 392:24:@2368.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2368.4]
  wire  m_0_clock; // @[MemPrimitives.scala 398:56:@2382.4]
  wire [4:0] m_0_io_r_ofs_0; // @[MemPrimitives.scala 398:56:@2382.4]
  wire [4:0] m_0_io_w_ofs_0; // @[MemPrimitives.scala 398:56:@2382.4]
  wire [95:0] m_0_io_w_data_0; // @[MemPrimitives.scala 398:56:@2382.4]
  wire  m_0_io_w_en_0; // @[MemPrimitives.scala 398:56:@2382.4]
  wire [95:0] m_0_io_output; // @[MemPrimitives.scala 398:56:@2382.4]
  wire [6:0] enqCompactor_io_headCnt; // @[MemPrimitives.scala 402:28:@2398.4]
  wire [95:0] enqCompactor_io_in_0_data; // @[MemPrimitives.scala 402:28:@2398.4]
  wire  enqCompactor_io_in_0_en; // @[MemPrimitives.scala 402:28:@2398.4]
  wire [95:0] enqCompactor_io_out_0_data; // @[MemPrimitives.scala 402:28:@2398.4]
  wire  enqCompactor_io_out_0_en; // @[MemPrimitives.scala 402:28:@2398.4]
  wire [6:0] deqCompactor_io_tailCnt; // @[MemPrimitives.scala 421:28:@2420.4]
  wire [95:0] deqCompactor_io_input_data_0; // @[MemPrimitives.scala 421:28:@2420.4]
  wire [95:0] deqCompactor_io_output_0; // @[MemPrimitives.scala 421:28:@2420.4]
  wire [6:0] _GEN_0; // @[Math.scala 53:59:@2409.4]
  wire [6:0] active_w_bank; // @[Math.scala 53:59:@2409.4]
  wire [7:0] active_w_addr; // @[Math.scala 52:59:@2410.4]
  wire  _T_102; // @[MemPrimitives.scala 414:38:@2411.4]
  wire [8:0] _T_104; // @[MemPrimitives.scala 414:69:@2412.4]
  wire [7:0] _T_105; // @[MemPrimitives.scala 414:69:@2413.4]
  wire [7:0] _T_106; // @[MemPrimitives.scala 414:69:@2414.4]
  wire [7:0] _T_107; // @[MemPrimitives.scala 414:19:@2415.4]
  wire [7:0] _T_108; // @[MemPrimitives.scala 415:32:@2416.4]
  wire [6:0] _GEN_1; // @[Math.scala 53:59:@2428.4]
  wire [6:0] active_r_bank; // @[Math.scala 53:59:@2428.4]
  wire [7:0] active_r_addr; // @[Math.scala 52:59:@2429.4]
  wire  _T_112; // @[MemPrimitives.scala 427:38:@2430.4]
  wire [8:0] _T_114; // @[MemPrimitives.scala 427:69:@2431.4]
  wire [7:0] _T_115; // @[MemPrimitives.scala 427:69:@2432.4]
  wire [7:0] _T_116; // @[MemPrimitives.scala 427:69:@2433.4]
  wire [7:0] _T_117; // @[MemPrimitives.scala 427:19:@2434.4]
  wire [7:0] _T_118; // @[MemPrimitives.scala 428:32:@2435.4]
  CompactingCounter headCtr ( // @[MemPrimitives.scala 381:23:@2346.4]
    .clock(headCtr_clock),
    .reset(headCtr_reset),
    .io_input_reset(headCtr_io_input_reset),
    .io_input_enables_0(headCtr_io_input_enables_0),
    .io_output_count(headCtr_io_output_count)
  );
  CompactingCounter tailCtr ( // @[MemPrimitives.scala 382:23:@2354.4]
    .clock(tailCtr_clock),
    .reset(tailCtr_reset),
    .io_input_reset(tailCtr_io_input_reset),
    .io_input_enables_0(tailCtr_io_input_enables_0),
    .io_output_count(tailCtr_io_output_count)
  );
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2368.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_empty(elements_io_output_empty),
    .io_output_full(elements_io_output_full)
  );
  Mem1D_3 m_0 ( // @[MemPrimitives.scala 398:56:@2382.4]
    .clock(m_0_clock),
    .io_r_ofs_0(m_0_io_r_ofs_0),
    .io_w_ofs_0(m_0_io_w_ofs_0),
    .io_w_data_0(m_0_io_w_data_0),
    .io_w_en_0(m_0_io_w_en_0),
    .io_output(m_0_io_output)
  );
  CompactingEnqNetwork enqCompactor ( // @[MemPrimitives.scala 402:28:@2398.4]
    .io_headCnt(enqCompactor_io_headCnt),
    .io_in_0_data(enqCompactor_io_in_0_data),
    .io_in_0_en(enqCompactor_io_in_0_en),
    .io_out_0_data(enqCompactor_io_out_0_data),
    .io_out_0_en(enqCompactor_io_out_0_en)
  );
  CompactingDeqNetwork deqCompactor ( // @[MemPrimitives.scala 421:28:@2420.4]
    .io_tailCnt(deqCompactor_io_tailCnt),
    .io_input_data_0(deqCompactor_io_input_data_0),
    .io_output_0(deqCompactor_io_output_0)
  );
  assign _GEN_0 = $signed(headCtr_io_output_count) % $signed(7'sh1); // @[Math.scala 53:59:@2409.4]
  assign active_w_bank = _GEN_0[6:0]; // @[Math.scala 53:59:@2409.4]
  assign active_w_addr = $signed(headCtr_io_output_count) / $signed(7'sh1); // @[Math.scala 52:59:@2410.4]
  assign _T_102 = $signed(7'sh0) < $signed(active_w_bank); // @[MemPrimitives.scala 414:38:@2411.4]
  assign _T_104 = $signed(active_w_addr) + $signed(8'sh1); // @[MemPrimitives.scala 414:69:@2412.4]
  assign _T_105 = $signed(active_w_addr) + $signed(8'sh1); // @[MemPrimitives.scala 414:69:@2413.4]
  assign _T_106 = $signed(_T_105); // @[MemPrimitives.scala 414:69:@2414.4]
  assign _T_107 = _T_102 ? $signed(_T_106) : $signed(active_w_addr); // @[MemPrimitives.scala 414:19:@2415.4]
  assign _T_108 = $unsigned(_T_107); // @[MemPrimitives.scala 415:32:@2416.4]
  assign _GEN_1 = $signed(tailCtr_io_output_count) % $signed(7'sh1); // @[Math.scala 53:59:@2428.4]
  assign active_r_bank = _GEN_1[6:0]; // @[Math.scala 53:59:@2428.4]
  assign active_r_addr = $signed(tailCtr_io_output_count) / $signed(7'sh1); // @[Math.scala 52:59:@2429.4]
  assign _T_112 = $signed(7'sh0) < $signed(active_r_bank); // @[MemPrimitives.scala 427:38:@2430.4]
  assign _T_114 = $signed(active_r_addr) + $signed(8'sh1); // @[MemPrimitives.scala 427:69:@2431.4]
  assign _T_115 = $signed(active_r_addr) + $signed(8'sh1); // @[MemPrimitives.scala 427:69:@2432.4]
  assign _T_116 = $signed(_T_115); // @[MemPrimitives.scala 427:69:@2433.4]
  assign _T_117 = _T_112 ? $signed(_T_116) : $signed(active_r_addr); // @[MemPrimitives.scala 427:19:@2434.4]
  assign _T_118 = $unsigned(_T_117); // @[MemPrimitives.scala 428:32:@2435.4]
  assign io_rPort_0_output_0 = deqCompactor_io_output_0; // @[MemPrimitives.scala 432:82:@2439.4]
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 439:39:@2443.4]
  assign io_empty = elements_io_output_empty; // @[MemPrimitives.scala 438:40:@2442.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 437:129:@2440.4]
  assign headCtr_clock = clock; // @[:@2347.4]
  assign headCtr_reset = reset; // @[:@2348.4]
  assign headCtr_io_input_reset = reset; // @[MemPrimitives.scala 385:26:@2364.4]
  assign headCtr_io_input_enables_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 383:129:@2362.4]
  assign tailCtr_clock = clock; // @[:@2355.4]
  assign tailCtr_reset = reset; // @[:@2356.4]
  assign tailCtr_io_input_reset = reset; // @[MemPrimitives.scala 386:26:@2365.4]
  assign tailCtr_io_input_enables_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 384:129:@2363.4]
  assign elements_clock = clock; // @[:@2369.4]
  assign elements_reset = reset; // @[:@2370.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 394:79:@2380.4]
  assign elements_io_input_dinc_en_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 395:80:@2381.4]
  assign m_0_clock = clock; // @[:@2383.4]
  assign m_0_io_r_ofs_0 = _T_118[4:0]; // @[MemPrimitives.scala 428:24:@2436.4]
  assign m_0_io_w_ofs_0 = _T_108[4:0]; // @[MemPrimitives.scala 415:24:@2417.4]
  assign m_0_io_w_data_0 = enqCompactor_io_out_0_data; // @[MemPrimitives.scala 416:25:@2418.4]
  assign m_0_io_w_en_0 = enqCompactor_io_out_0_en; // @[MemPrimitives.scala 417:25:@2419.4]
  assign enqCompactor_io_headCnt = headCtr_io_output_count; // @[MemPrimitives.scala 404:27:@2406.4]
  assign enqCompactor_io_in_0_data = io_wPort_0_data_0; // @[MemPrimitives.scala 406:90:@2407.4]
  assign enqCompactor_io_in_0_en = io_wPort_0_en_0; // @[MemPrimitives.scala 407:85:@2408.4]
  assign deqCompactor_io_tailCnt = tailCtr_io_output_count; // @[MemPrimitives.scala 423:27:@2427.4]
  assign deqCompactor_io_input_data_0 = m_0_io_output; // @[MemPrimitives.scala 429:35:@2437.4]
endmodule
module FF_3( // @[:@2449.2]
  input        clock, // @[:@2450.4]
  input        reset, // @[:@2451.4]
  output [8:0] io_rPort_0_output_0, // @[:@2452.4]
  input  [8:0] io_wPort_0_data_0, // @[:@2452.4]
  input        io_wPort_0_reset, // @[:@2452.4]
  input        io_wPort_0_en_0 // @[:@2452.4]
);
  reg [8:0] ff; // @[MemPrimitives.scala 321:19:@2467.4]
  reg [31:0] _RAND_0;
  wire [8:0] _T_68; // @[MemPrimitives.scala 325:32:@2469.4]
  wire [8:0] _T_69; // @[MemPrimitives.scala 325:12:@2470.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@2469.4]
  assign _T_69 = io_wPort_0_reset ? 9'h0 : _T_68; // @[MemPrimitives.scala 325:12:@2470.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@2472.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 9'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 9'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@2487.2]
  input        clock, // @[:@2488.4]
  input        reset, // @[:@2489.4]
  input        io_setup_saturate, // @[:@2490.4]
  input        io_input_reset, // @[:@2490.4]
  input        io_input_enable, // @[:@2490.4]
  output [8:0] io_output_count_0, // @[:@2490.4]
  output       io_output_oobs_0, // @[:@2490.4]
  output       io_output_done // @[:@2490.4]
);
  wire  bases_0_clock; // @[Counter.scala 262:53:@2503.4]
  wire  bases_0_reset; // @[Counter.scala 262:53:@2503.4]
  wire [8:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 262:53:@2503.4]
  wire [8:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 262:53:@2503.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 262:53:@2503.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 262:53:@2503.4]
  wire  SRFF_clock; // @[Counter.scala 264:22:@2519.4]
  wire  SRFF_reset; // @[Counter.scala 264:22:@2519.4]
  wire  SRFF_io_input_set; // @[Counter.scala 264:22:@2519.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 264:22:@2519.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 264:22:@2519.4]
  wire  SRFF_io_output; // @[Counter.scala 264:22:@2519.4]
  wire  _T_36; // @[Counter.scala 265:45:@2522.4]
  wire [8:0] _T_48; // @[Counter.scala 288:52:@2547.4]
  wire [9:0] _T_50; // @[Counter.scala 292:33:@2548.4]
  wire [8:0] _T_51; // @[Counter.scala 292:33:@2549.4]
  wire [8:0] _T_52; // @[Counter.scala 292:33:@2550.4]
  wire  _T_57; // @[Counter.scala 294:18:@2552.4]
  wire [8:0] _T_68; // @[Counter.scala 300:115:@2560.4]
  wire [8:0] _T_70; // @[Counter.scala 300:85:@2562.4]
  wire [8:0] _T_71; // @[Counter.scala 300:152:@2563.4]
  wire [8:0] _T_72; // @[Counter.scala 300:74:@2564.4]
  wire  _T_75; // @[Counter.scala 323:102:@2568.4]
  wire  _T_77; // @[Counter.scala 323:130:@2569.4]
  FF_3 bases_0 ( // @[Counter.scala 262:53:@2503.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 264:22:@2519.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 265:45:@2522.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 288:52:@2547.4]
  assign _T_50 = $signed(_T_48) + $signed(9'sh1); // @[Counter.scala 292:33:@2548.4]
  assign _T_51 = $signed(_T_48) + $signed(9'sh1); // @[Counter.scala 292:33:@2549.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 292:33:@2550.4]
  assign _T_57 = $signed(_T_52) >= $signed(9'sh64); // @[Counter.scala 294:18:@2552.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 300:115:@2560.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 9'h0; // @[Counter.scala 300:85:@2562.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 300:152:@2563.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 300:74:@2564.4]
  assign _T_75 = $signed(_T_48) < $signed(9'sh0); // @[Counter.scala 323:102:@2568.4]
  assign _T_77 = $signed(_T_48) >= $signed(9'sh64); // @[Counter.scala 323:130:@2569.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 305:28:@2567.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 323:60:@2571.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 334:20:@2573.4]
  assign bases_0_clock = clock; // @[:@2504.4]
  assign bases_0_reset = reset; // @[:@2505.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 9'h0 : _T_72; // @[Counter.scala 300:31:@2566.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 282:27:@2545.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 285:29:@2546.4]
  assign SRFF_clock = clock; // @[:@2520.4]
  assign SRFF_reset = reset; // @[:@2521.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 265:23:@2524.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 266:25:@2526.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 267:30:@2527.4]
endmodule
module x478_ctrchain( // @[:@2578.2]
  input        clock, // @[:@2579.4]
  input        reset, // @[:@2580.4]
  input        io_input_reset, // @[:@2581.4]
  input        io_input_enable, // @[:@2581.4]
  output [8:0] io_output_counts_0, // @[:@2581.4]
  output       io_output_oobs_0, // @[:@2581.4]
  output       io_output_done // @[:@2581.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 514:46:@2583.4]
  wire  ctrs_0_reset; // @[Counter.scala 514:46:@2583.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 514:46:@2583.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 514:46:@2583.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 514:46:@2583.4]
  wire [8:0] ctrs_0_io_output_count_0; // @[Counter.scala 514:46:@2583.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 514:46:@2583.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 514:46:@2583.4]
  reg  wasDone; // @[Counter.scala 543:24:@2592.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 547:69:@2598.4]
  wire  _T_47; // @[Counter.scala 547:80:@2599.4]
  reg  doneLatch; // @[Counter.scala 551:26:@2604.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 552:48:@2605.4]
  wire  _T_55; // @[Counter.scala 552:19:@2606.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 514:46:@2583.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 547:69:@2598.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 547:80:@2599.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 552:48:@2605.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 552:19:@2606.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 558:32:@2608.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 559:30:@2610.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 547:18:@2601.4]
  assign ctrs_0_clock = clock; // @[:@2584.4]
  assign ctrs_0_reset = reset; // @[:@2585.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 531:29:@2591.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 521:24:@2589.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 525:33:@2590.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@2650.2]
  input   clock, // @[:@2651.4]
  input   reset, // @[:@2652.4]
  input   io_flow, // @[:@2653.4]
  input   io_in, // @[:@2653.4]
  output  io_out // @[:@2653.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2655.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2655.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2655.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2655.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2655.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2655.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@2655.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2668.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2667.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2666.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2665.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2664.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2662.4]
endmodule
module RetimeWrapper_25( // @[:@2778.2]
  input   clock, // @[:@2779.4]
  input   reset, // @[:@2780.4]
  input   io_flow, // @[:@2781.4]
  input   io_in, // @[:@2781.4]
  output  io_out // @[:@2781.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2783.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2783.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2783.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2783.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2783.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2783.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@2783.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2796.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2795.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2794.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2793.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2792.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2790.4]
endmodule
module x499_inr_Foreach_sm( // @[:@2798.2]
  input   clock, // @[:@2799.4]
  input   reset, // @[:@2800.4]
  input   io_enable, // @[:@2801.4]
  output  io_done, // @[:@2801.4]
  output  io_doneLatch, // @[:@2801.4]
  input   io_rst, // @[:@2801.4]
  input   io_ctrDone, // @[:@2801.4]
  output  io_datapathEn, // @[:@2801.4]
  output  io_ctrInc, // @[:@2801.4]
  output  io_ctrRst, // @[:@2801.4]
  input   io_parentAck, // @[:@2801.4]
  input   io_backpressure, // @[:@2801.4]
  input   io_break // @[:@2801.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@2803.4]
  wire  active_reset; // @[Controllers.scala 261:22:@2803.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@2803.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@2803.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@2803.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@2803.4]
  wire  done_clock; // @[Controllers.scala 262:20:@2806.4]
  wire  done_reset; // @[Controllers.scala 262:20:@2806.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@2806.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@2806.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@2806.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@2806.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2840.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2840.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2840.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2840.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2840.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2862.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2862.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2862.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2862.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2862.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2874.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2874.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2874.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2874.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2874.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2882.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2882.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2882.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2882.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2882.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2898.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2898.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2898.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2898.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2898.4]
  wire  _T_80; // @[Controllers.scala 264:48:@2811.4]
  wire  _T_81; // @[Controllers.scala 264:46:@2812.4]
  wire  _T_82; // @[Controllers.scala 264:62:@2813.4]
  wire  _T_83; // @[Controllers.scala 264:60:@2814.4]
  wire  _T_100; // @[package.scala 100:49:@2831.4]
  reg  _T_103; // @[package.scala 48:56:@2832.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@2845.4 package.scala 96:25:@2846.4]
  wire  _T_110; // @[package.scala 100:49:@2847.4]
  reg  _T_113; // @[package.scala 48:56:@2848.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@2850.4]
  wire  _T_118; // @[Controllers.scala 283:41:@2855.4]
  wire  _T_119; // @[Controllers.scala 283:59:@2856.4]
  wire  _T_121; // @[Controllers.scala 284:37:@2859.4]
  wire  _T_124; // @[package.scala 96:25:@2867.4 package.scala 96:25:@2868.4]
  wire  _T_126; // @[package.scala 100:49:@2869.4]
  reg  _T_129; // @[package.scala 48:56:@2870.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@2892.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@2894.4]
  reg  _T_153; // @[package.scala 48:56:@2895.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@2903.4 package.scala 96:25:@2904.4]
  wire  _T_158; // @[Controllers.scala 292:61:@2905.4]
  wire  _T_159; // @[Controllers.scala 292:24:@2906.4]
  SRFF active ( // @[Controllers.scala 261:22:@2803.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@2806.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@2840.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@2862.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2874.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2882.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@2898.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@2811.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@2812.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@2813.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@2814.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@2831.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@2845.4 package.scala 96:25:@2846.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@2847.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@2850.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@2855.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@2856.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@2859.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2867.4 package.scala 96:25:@2868.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@2869.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@2894.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@2903.4 package.scala 96:25:@2904.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@2905.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@2906.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@2873.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@2908.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@2858.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@2861.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@2853.4]
  assign active_clock = clock; // @[:@2804.4]
  assign active_reset = reset; // @[:@2805.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@2816.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@2820.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@2821.4]
  assign done_clock = clock; // @[:@2807.4]
  assign done_reset = reset; // @[:@2808.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@2836.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@2829.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@2830.4]
  assign RetimeWrapper_clock = clock; // @[:@2841.4]
  assign RetimeWrapper_reset = reset; // @[:@2842.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@2844.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@2843.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2863.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2864.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@2866.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@2865.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2875.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2876.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2878.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@2877.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2883.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2884.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2886.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@2885.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2899.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2900.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@2902.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@2901.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x499_inr_Foreach_iiCtr( // @[:@2911.2]
  input   clock, // @[:@2912.4]
  input   reset, // @[:@2913.4]
  input   io_input_enable, // @[:@2914.4]
  input   io_input_reset, // @[:@2914.4]
  output  io_output_issue, // @[:@2914.4]
  output  io_output_done // @[:@2914.4]
);
  reg [4:0] _T_15; // @[Counter.scala 135:22:@2916.4]
  reg [31:0] _RAND_0;
  wire  _T_17; // @[Counter.scala 138:24:@2917.4]
  wire  _T_20; // @[Counter.scala 139:23:@2919.4]
  wire [5:0] _T_26; // @[Counter.scala 141:68:@2922.4]
  wire [4:0] _T_27; // @[Counter.scala 141:68:@2923.4]
  wire [4:0] _T_28; // @[Counter.scala 141:68:@2924.4]
  wire [4:0] _T_29; // @[Counter.scala 141:23:@2925.4]
  wire [4:0] _T_30; // @[Counter.scala 142:19:@2926.4]
  wire [4:0] _T_32; // @[Counter.scala 143:15:@2927.4]
  assign _T_17 = $signed(_T_15) == $signed(5'sh4); // @[Counter.scala 138:24:@2917.4]
  assign _T_20 = $signed(_T_15) == $signed(5'sh0); // @[Counter.scala 139:23:@2919.4]
  assign _T_26 = $signed(_T_15) - $signed(5'sh1); // @[Counter.scala 141:68:@2922.4]
  assign _T_27 = $signed(_T_15) - $signed(5'sh1); // @[Counter.scala 141:68:@2923.4]
  assign _T_28 = $signed(_T_27); // @[Counter.scala 141:68:@2924.4]
  assign _T_29 = _T_20 ? $signed(5'sh4) : $signed(_T_28); // @[Counter.scala 141:23:@2925.4]
  assign _T_30 = io_input_enable ? $signed(_T_29) : $signed(_T_15); // @[Counter.scala 142:19:@2926.4]
  assign _T_32 = io_input_reset ? $signed(5'sh4) : $signed(_T_30); // @[Counter.scala 143:15:@2927.4]
  assign io_output_issue = _T_17 & io_input_enable; // @[Counter.scala 146:21:@2930.4]
  assign io_output_done = _T_20 & io_input_enable; // @[Counter.scala 145:20:@2929.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 5'sh4;
    end else begin
      if (io_input_reset) begin
        _T_15 <= 5'sh4;
      end else begin
        if (io_input_enable) begin
          if (_T_20) begin
            _T_15 <= 5'sh4;
          end else begin
            _T_15 <= _T_28;
          end
        end
      end
    end
  end
endmodule
module fix2fixBox( // @[:@3060.2]
  input  [31:0] io_a, // @[:@3063.4]
  output [31:0] io_b // @[:@3063.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@3076.4]
endmodule
module _( // @[:@3078.2]
  input  [31:0] io_b, // @[:@3081.4]
  output [31:0] io_result // @[:@3081.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3086.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3086.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@3086.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3094.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3089.4]
endmodule
module fix2fixBox_1( // @[:@3128.2]
  input  [31:0] io_a, // @[:@3131.4]
  output [32:0] io_b // @[:@3131.4]
);
  wire  _T_20; // @[implicits.scala 70:16:@3141.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 70:16:@3141.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@3146.4]
endmodule
module __1( // @[:@3148.2]
  input  [31:0] io_b, // @[:@3151.4]
  output [32:0] io_result // @[:@3151.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3156.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3156.4]
  fix2fixBox_1 fix2fixBox ( // @[BigIPZynq.scala 219:30:@3156.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3164.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3159.4]
endmodule
module RetimeWrapper_31( // @[:@3216.2]
  input         clock, // @[:@3217.4]
  input         reset, // @[:@3218.4]
  input         io_flow, // @[:@3219.4]
  input  [31:0] io_in, // @[:@3219.4]
  output [31:0] io_out // @[:@3219.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3221.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3221.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3221.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3221.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3221.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3221.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3221.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3234.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3233.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3232.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3231.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3230.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3228.4]
endmodule
module fix2fixBox_3( // @[:@3236.2]
  input         clock, // @[:@3237.4]
  input         reset, // @[:@3238.4]
  input  [32:0] io_a, // @[:@3239.4]
  input         io_flow, // @[:@3239.4]
  output [31:0] io_b // @[:@3239.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3252.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3252.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3252.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3252.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3252.4]
  RetimeWrapper_31 RetimeWrapper ( // @[package.scala 93:22:@3252.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3259.4]
  assign RetimeWrapper_clock = clock; // @[:@3253.4]
  assign RetimeWrapper_reset = reset; // @[:@3254.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3256.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3255.4]
endmodule
module x739_sum( // @[:@3261.2]
  input         clock, // @[:@3262.4]
  input         reset, // @[:@3263.4]
  input  [31:0] io_a, // @[:@3264.4]
  input  [31:0] io_b, // @[:@3264.4]
  input         io_flow, // @[:@3264.4]
  output [31:0] io_result // @[:@3264.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@3272.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@3272.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@3279.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@3279.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@3297.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@3297.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@3297.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@3297.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@3297.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@3277.4 Math.scala 724:14:@3278.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@3284.4 Math.scala 724:14:@3285.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@3286.4]
  __1 _ ( // @[Math.scala 720:24:@3272.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __1 __1 ( // @[Math.scala 720:24:@3279.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_3 fix2fixBox ( // @[Math.scala 141:30:@3297.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@3277.4 Math.scala 724:14:@3278.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@3284.4 Math.scala 724:14:@3285.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@3286.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@3305.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@3275.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@3282.4]
  assign fix2fixBox_clock = clock; // @[:@3298.4]
  assign fix2fixBox_reset = reset; // @[:@3299.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@3300.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@3303.4]
endmodule
module x485_sub( // @[:@3440.2]
  input         clock, // @[:@3441.4]
  input         reset, // @[:@3442.4]
  input  [31:0] io_a, // @[:@3443.4]
  input  [31:0] io_b, // @[:@3443.4]
  input         io_flow, // @[:@3443.4]
  output [31:0] io_result // @[:@3443.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@3451.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@3451.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@3458.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@3458.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@3477.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@3477.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@3477.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@3477.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@3477.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@3456.4 Math.scala 724:14:@3457.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@3463.4 Math.scala 724:14:@3464.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@3465.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@3466.4]
  __1 _ ( // @[Math.scala 720:24:@3451.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __1 __1 ( // @[Math.scala 720:24:@3458.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_3 fix2fixBox ( // @[Math.scala 182:30:@3477.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@3456.4 Math.scala 724:14:@3457.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@3463.4 Math.scala 724:14:@3464.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@3465.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@3466.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@3485.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@3454.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@3461.4]
  assign fix2fixBox_clock = clock; // @[:@3478.4]
  assign fix2fixBox_reset = reset; // @[:@3479.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@3480.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@3483.4]
endmodule
module RetimeWrapper_35( // @[:@3857.2]
  input         clock, // @[:@3858.4]
  input         reset, // @[:@3859.4]
  input         io_flow, // @[:@3860.4]
  input  [35:0] io_in, // @[:@3860.4]
  output [35:0] io_out // @[:@3860.4]
);
  wire [35:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3862.4]
  wire [35:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3862.4]
  wire [35:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3862.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3862.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3862.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3862.4]
  RetimeShiftRegister #(.WIDTH(36), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3862.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3875.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3874.4]
  assign sr_init = 36'h0; // @[RetimeShiftRegister.scala 19:16:@3873.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3872.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3871.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3869.4]
endmodule
module RetimeWrapper_36( // @[:@3889.2]
  input         clock, // @[:@3890.4]
  input         reset, // @[:@3891.4]
  input         io_flow, // @[:@3892.4]
  input  [37:0] io_in, // @[:@3892.4]
  output [37:0] io_out // @[:@3892.4]
);
  wire [37:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3894.4]
  wire [37:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3894.4]
  wire [37:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3894.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3894.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3894.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3894.4]
  RetimeShiftRegister #(.WIDTH(38), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3894.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3907.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3906.4]
  assign sr_init = 38'h0; // @[RetimeShiftRegister.scala 19:16:@3905.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3904.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3903.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3901.4]
endmodule
module fix2fixBox_13( // @[:@3909.2]
  input  [31:0] io_a, // @[:@3912.4]
  output [63:0] io_b // @[:@3912.4]
);
  wire  _T_20; // @[implicits.scala 70:16:@3922.4]
  wire [31:0] _T_24; // @[Bitwise.scala 72:12:@3925.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 70:16:@3922.4]
  assign _T_24 = _T_20 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@3925.4]
  assign io_b = {_T_24,io_a}; // @[Converter.scala 95:38:@3929.4]
endmodule
module x491( // @[:@3931.2]
  input  [31:0] io_b, // @[:@3934.4]
  output [63:0] io_result // @[:@3934.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3939.4]
  wire [63:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3939.4]
  fix2fixBox_13 fix2fixBox ( // @[BigIPZynq.scala 219:30:@3939.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3947.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3942.4]
endmodule
module RetimeWrapper_37( // @[:@3961.2]
  input         clock, // @[:@3962.4]
  input         reset, // @[:@3963.4]
  input         io_flow, // @[:@3964.4]
  input  [63:0] io_in, // @[:@3964.4]
  output [63:0] io_out // @[:@3964.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3966.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3966.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3966.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3966.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3966.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3966.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3966.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3979.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3978.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@3977.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3976.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3975.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3973.4]
endmodule
module fix2fixBox_14( // @[:@3981.2]
  input  [63:0] io_a, // @[:@3984.4]
  output [64:0] io_b // @[:@3984.4]
);
  wire  _T_20; // @[implicits.scala 70:16:@3994.4]
  assign _T_20 = io_a[63]; // @[implicits.scala 70:16:@3994.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@3999.4]
endmodule
module __9( // @[:@4001.2]
  input  [63:0] io_b, // @[:@4004.4]
  output [64:0] io_result // @[:@4004.4]
);
  wire [63:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@4009.4]
  wire [64:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@4009.4]
  fix2fixBox_14 fix2fixBox ( // @[BigIPZynq.scala 219:30:@4009.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@4017.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@4012.4]
endmodule
module RetimeWrapper_38( // @[:@4069.2]
  input         clock, // @[:@4070.4]
  input         reset, // @[:@4071.4]
  input         io_flow, // @[:@4072.4]
  input  [63:0] io_in, // @[:@4072.4]
  output [63:0] io_out // @[:@4072.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@4074.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@4074.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@4074.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@4074.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@4074.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@4074.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@4074.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@4087.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@4086.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@4085.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@4084.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@4083.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@4081.4]
endmodule
module fix2fixBox_16( // @[:@4089.2]
  input         clock, // @[:@4090.4]
  input         reset, // @[:@4091.4]
  input  [64:0] io_a, // @[:@4092.4]
  input         io_flow, // @[:@4092.4]
  output [63:0] io_b // @[:@4092.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4105.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4105.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4105.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@4105.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@4105.4]
  RetimeWrapper_38 RetimeWrapper ( // @[package.scala 93:22:@4105.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@4112.4]
  assign RetimeWrapper_clock = clock; // @[:@4106.4]
  assign RetimeWrapper_reset = reset; // @[:@4107.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@4109.4]
  assign RetimeWrapper_io_in = io_a[63:0]; // @[package.scala 94:16:@4108.4]
endmodule
module x493_sum( // @[:@4114.2]
  input         clock, // @[:@4115.4]
  input         reset, // @[:@4116.4]
  input  [63:0] io_a, // @[:@4117.4]
  input  [63:0] io_b, // @[:@4117.4]
  input         io_flow, // @[:@4117.4]
  output [63:0] io_result // @[:@4117.4]
);
  wire [63:0] __io_b; // @[Math.scala 720:24:@4125.4]
  wire [64:0] __io_result; // @[Math.scala 720:24:@4125.4]
  wire [63:0] __1_io_b; // @[Math.scala 720:24:@4132.4]
  wire [64:0] __1_io_result; // @[Math.scala 720:24:@4132.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4150.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4150.4]
  wire [64:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4150.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4150.4]
  wire [63:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4150.4]
  wire [64:0] a_upcast_number; // @[Math.scala 723:22:@4130.4 Math.scala 724:14:@4131.4]
  wire [64:0] b_upcast_number; // @[Math.scala 723:22:@4137.4 Math.scala 724:14:@4138.4]
  wire [65:0] _T_21; // @[Math.scala 136:37:@4139.4]
  __9 _ ( // @[Math.scala 720:24:@4125.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __9 __1 ( // @[Math.scala 720:24:@4132.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_16 fix2fixBox ( // @[Math.scala 141:30:@4150.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@4130.4 Math.scala 724:14:@4131.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@4137.4 Math.scala 724:14:@4138.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4139.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4158.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@4128.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@4135.4]
  assign fix2fixBox_clock = clock; // @[:@4151.4]
  assign fix2fixBox_reset = reset; // @[:@4152.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4153.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4156.4]
endmodule
module RetimeWrapper_44( // @[:@4332.2]
  input         clock, // @[:@4333.4]
  input         reset, // @[:@4334.4]
  input         io_flow, // @[:@4335.4]
  input  [31:0] io_in, // @[:@4335.4]
  output [31:0] io_out // @[:@4335.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@4337.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@4337.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@4337.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@4337.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@4337.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@4337.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@4337.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@4350.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@4349.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@4348.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@4347.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@4346.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@4344.4]
endmodule
module x499_inr_Foreach_kernelx499_inr_Foreach_concrete1( // @[:@4384.2]
  input         clock, // @[:@4385.4]
  input         reset, // @[:@4386.4]
  input  [63:0] io_in_x468_A_dram_number, // @[:@4387.4]
  output [95:0] io_in_x475_fifo_wPort_0_data_0, // @[:@4387.4]
  output        io_in_x475_fifo_wPort_0_en_0, // @[:@4387.4]
  input         io_in_x475_fifo_full, // @[:@4387.4]
  output        io_in_x475_fifo_active_0_in, // @[:@4387.4]
  input         io_in_x475_fifo_active_0_out, // @[:@4387.4]
  input         io_in_x474_ready, // @[:@4387.4]
  output        io_in_x474_valid, // @[:@4387.4]
  output [63:0] io_in_x474_bits_addr, // @[:@4387.4]
  output [31:0] io_in_x474_bits_size, // @[:@4387.4]
  input         io_sigsIn_iiIssue, // @[:@4387.4]
  input         io_sigsIn_backpressure, // @[:@4387.4]
  input         io_sigsIn_datapathEn, // @[:@4387.4]
  input         io_sigsIn_break, // @[:@4387.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@4387.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@4387.4]
  input         io_rr // @[:@4387.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4423.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@4423.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4434.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4434.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4434.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@4434.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@4434.4]
  wire  x739_sum_1_clock; // @[Math.scala 150:24:@4452.4]
  wire  x739_sum_1_reset; // @[Math.scala 150:24:@4452.4]
  wire [31:0] x739_sum_1_io_a; // @[Math.scala 150:24:@4452.4]
  wire [31:0] x739_sum_1_io_b; // @[Math.scala 150:24:@4452.4]
  wire  x739_sum_1_io_flow; // @[Math.scala 150:24:@4452.4]
  wire [31:0] x739_sum_1_io_result; // @[Math.scala 150:24:@4452.4]
  wire  x485_sub_1_clock; // @[Math.scala 191:24:@4489.4]
  wire  x485_sub_1_reset; // @[Math.scala 191:24:@4489.4]
  wire [31:0] x485_sub_1_io_a; // @[Math.scala 191:24:@4489.4]
  wire [31:0] x485_sub_1_io_b; // @[Math.scala 191:24:@4489.4]
  wire  x485_sub_1_io_flow; // @[Math.scala 191:24:@4489.4]
  wire [31:0] x485_sub_1_io_result; // @[Math.scala 191:24:@4489.4]
  wire  x486_sum_1_clock; // @[Math.scala 150:24:@4501.4]
  wire  x486_sum_1_reset; // @[Math.scala 150:24:@4501.4]
  wire [31:0] x486_sum_1_io_a; // @[Math.scala 150:24:@4501.4]
  wire [31:0] x486_sum_1_io_b; // @[Math.scala 150:24:@4501.4]
  wire  x486_sum_1_io_flow; // @[Math.scala 150:24:@4501.4]
  wire [31:0] x486_sum_1_io_result; // @[Math.scala 150:24:@4501.4]
  wire  x487_sum_1_clock; // @[Math.scala 150:24:@4513.4]
  wire  x487_sum_1_reset; // @[Math.scala 150:24:@4513.4]
  wire [31:0] x487_sum_1_io_a; // @[Math.scala 150:24:@4513.4]
  wire [31:0] x487_sum_1_io_b; // @[Math.scala 150:24:@4513.4]
  wire  x487_sum_1_io_flow; // @[Math.scala 150:24:@4513.4]
  wire [31:0] x487_sum_1_io_result; // @[Math.scala 150:24:@4513.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4542.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4542.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@4542.4]
  wire [35:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@4542.4]
  wire [35:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@4542.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@4554.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@4554.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@4554.4]
  wire [37:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@4554.4]
  wire [37:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@4554.4]
  wire [31:0] x491_1_io_b; // @[Math.scala 720:24:@4564.4]
  wire [63:0] x491_1_io_result; // @[Math.scala 720:24:@4564.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@4574.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@4574.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@4574.4]
  wire [63:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@4574.4]
  wire [63:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@4574.4]
  wire  x493_sum_1_clock; // @[Math.scala 150:24:@4583.4]
  wire  x493_sum_1_reset; // @[Math.scala 150:24:@4583.4]
  wire [63:0] x493_sum_1_io_a; // @[Math.scala 150:24:@4583.4]
  wire [63:0] x493_sum_1_io_b; // @[Math.scala 150:24:@4583.4]
  wire  x493_sum_1_io_flow; // @[Math.scala 150:24:@4583.4]
  wire [63:0] x493_sum_1_io_result; // @[Math.scala 150:24:@4583.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@4594.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@4594.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@4594.4]
  wire [63:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@4594.4]
  wire [63:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@4594.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@4608.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@4608.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@4608.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@4608.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@4608.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@4618.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@4618.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@4618.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@4618.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@4618.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@4628.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@4628.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@4628.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@4628.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@4628.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@4646.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@4646.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@4646.4]
  wire [31:0] RetimeWrapper_8_io_in; // @[package.scala 93:22:@4646.4]
  wire [31:0] RetimeWrapper_8_io_out; // @[package.scala 93:22:@4646.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@4656.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@4656.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@4656.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@4656.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@4656.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@4672.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@4672.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@4672.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@4672.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@4672.4]
  wire  _T_323; // @[package.scala 96:25:@4439.4 package.scala 96:25:@4440.4]
  wire  _T_326; // @[sm_x499_inr_Foreach.scala 70:18:@4442.4]
  wire  _T_327; // @[sm_x499_inr_Foreach.scala 70:45:@4443.4]
  wire  _T_328; // @[sm_x499_inr_Foreach.scala 70:43:@4444.4]
  wire [31:0] b479_number; // @[Math.scala 723:22:@4428.4 Math.scala 724:14:@4429.4]
  wire [32:0] _GEN_0; // @[Math.scala 461:32:@4448.4]
  wire [32:0] _T_331; // @[Math.scala 461:32:@4448.4]
  wire [31:0] x739_sum_number; // @[Math.scala 154:22:@4458.4 Math.scala 155:14:@4459.4]
  wire  _T_337; // @[FixedPoint.scala 50:25:@4463.4]
  wire [3:0] _T_341; // @[Bitwise.scala 72:12:@4465.4]
  wire [27:0] _T_342; // @[FixedPoint.scala 18:52:@4466.4]
  wire  _T_348; // @[Math.scala 451:55:@4468.4]
  wire [3:0] _T_349; // @[FixedPoint.scala 18:52:@4469.4]
  wire  _T_355; // @[Math.scala 451:110:@4471.4]
  wire  _T_356; // @[Math.scala 451:94:@4472.4]
  wire [31:0] _T_358; // @[Cat.scala 30:58:@4474.4]
  wire [31:0] x482_1_number; // @[Math.scala 454:20:@4475.4]
  wire [35:0] _GEN_1; // @[Math.scala 461:32:@4480.4]
  wire [35:0] _T_363; // @[Math.scala 461:32:@4480.4]
  wire [37:0] _GEN_2; // @[Math.scala 461:32:@4485.4]
  wire [37:0] _T_366; // @[Math.scala 461:32:@4485.4]
  wire [31:0] x487_sum_number; // @[Math.scala 154:22:@4519.4 Math.scala 155:14:@4520.4]
  wire  _T_386; // @[FixedPoint.scala 50:25:@4524.4]
  wire [3:0] _T_390; // @[Bitwise.scala 72:12:@4526.4]
  wire [27:0] _T_391; // @[FixedPoint.scala 18:52:@4527.4]
  wire  _T_397; // @[Math.scala 451:55:@4529.4]
  wire [3:0] _T_398; // @[FixedPoint.scala 18:52:@4530.4]
  wire  _T_404; // @[Math.scala 451:110:@4532.4]
  wire  _T_405; // @[Math.scala 451:94:@4533.4]
  wire [31:0] _T_407; // @[Cat.scala 30:58:@4535.4]
  wire [31:0] x488_1_number; // @[Math.scala 454:20:@4536.4]
  wire [35:0] _GEN_3; // @[Math.scala 461:32:@4541.4]
  wire [37:0] _GEN_4; // @[Math.scala 461:32:@4553.4]
  wire [37:0] _T_419; // @[package.scala 96:25:@4559.4 package.scala 96:25:@4560.4]
  wire [31:0] x741_1_number; // @[Math.scala 459:22:@4552.4 Math.scala 461:14:@4561.4]
  wire [63:0] x759_x493_sum_D1_number; // @[package.scala 96:25:@4599.4 package.scala 96:25:@4600.4]
  wire [96:0] x494_tuple; // @[Cat.scala 30:58:@4604.4]
  wire  _T_454; // @[package.scala 96:25:@4633.4 package.scala 96:25:@4634.4]
  wire  _T_456; // @[implicits.scala 56:10:@4635.4]
  wire  x760_x495_D4; // @[package.scala 96:25:@4613.4 package.scala 96:25:@4614.4]
  wire  _T_457; // @[sm_x499_inr_Foreach.scala 108:121:@4636.4]
  wire  x761_b480_D4; // @[package.scala 96:25:@4623.4 package.scala 96:25:@4624.4]
  wire  _T_458; // @[sm_x499_inr_Foreach.scala 108:127:@4637.4]
  wire [31:0] x762_x486_sum_D1_number; // @[package.scala 96:25:@4651.4 package.scala 96:25:@4652.4]
  wire [31:0] x763_x485_sub_D2_number; // @[package.scala 96:25:@4661.4 package.scala 96:25:@4662.4]
  wire [63:0] _T_473; // @[Cat.scala 30:58:@4665.4]
  wire [35:0] _T_414; // @[package.scala 96:25:@4547.4 package.scala 96:25:@4548.4]
  wire [31:0] x489_1_number; // @[Math.scala 459:22:@4540.4 Math.scala 461:14:@4549.4]
  wire  _T_475; // @[sm_x499_inr_Foreach.scala 121:121:@4668.4]
  wire  _T_481; // @[package.scala 96:25:@4677.4 package.scala 96:25:@4678.4]
  wire  _T_483; // @[implicits.scala 56:10:@4679.4]
  wire  _T_484; // @[sm_x499_inr_Foreach.scala 121:138:@4680.4]
  wire  _T_486; // @[sm_x499_inr_Foreach.scala 121:235:@4682.4]
  wire  _T_487; // @[sm_x499_inr_Foreach.scala 121:254:@4683.4]
  _ _ ( // @[Math.scala 720:24:@4423.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_25 RetimeWrapper ( // @[package.scala 93:22:@4434.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x739_sum x739_sum_1 ( // @[Math.scala 150:24:@4452.4]
    .clock(x739_sum_1_clock),
    .reset(x739_sum_1_reset),
    .io_a(x739_sum_1_io_a),
    .io_b(x739_sum_1_io_b),
    .io_flow(x739_sum_1_io_flow),
    .io_result(x739_sum_1_io_result)
  );
  x485_sub x485_sub_1 ( // @[Math.scala 191:24:@4489.4]
    .clock(x485_sub_1_clock),
    .reset(x485_sub_1_reset),
    .io_a(x485_sub_1_io_a),
    .io_b(x485_sub_1_io_b),
    .io_flow(x485_sub_1_io_flow),
    .io_result(x485_sub_1_io_result)
  );
  x739_sum x486_sum_1 ( // @[Math.scala 150:24:@4501.4]
    .clock(x486_sum_1_clock),
    .reset(x486_sum_1_reset),
    .io_a(x486_sum_1_io_a),
    .io_b(x486_sum_1_io_b),
    .io_flow(x486_sum_1_io_flow),
    .io_result(x486_sum_1_io_result)
  );
  x739_sum x487_sum_1 ( // @[Math.scala 150:24:@4513.4]
    .clock(x487_sum_1_clock),
    .reset(x487_sum_1_reset),
    .io_a(x487_sum_1_io_a),
    .io_b(x487_sum_1_io_b),
    .io_flow(x487_sum_1_io_flow),
    .io_result(x487_sum_1_io_result)
  );
  RetimeWrapper_35 RetimeWrapper_1 ( // @[package.scala 93:22:@4542.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_2 ( // @[package.scala 93:22:@4554.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x491 x491_1 ( // @[Math.scala 720:24:@4564.4]
    .io_b(x491_1_io_b),
    .io_result(x491_1_io_result)
  );
  RetimeWrapper_37 RetimeWrapper_3 ( // @[package.scala 93:22:@4574.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x493_sum x493_sum_1 ( // @[Math.scala 150:24:@4583.4]
    .clock(x493_sum_1_clock),
    .reset(x493_sum_1_reset),
    .io_a(x493_sum_1_io_a),
    .io_b(x493_sum_1_io_b),
    .io_flow(x493_sum_1_io_flow),
    .io_result(x493_sum_1_io_result)
  );
  RetimeWrapper_37 RetimeWrapper_4 ( // @[package.scala 93:22:@4594.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_5 ( // @[package.scala 93:22:@4608.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_6 ( // @[package.scala 93:22:@4618.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_7 ( // @[package.scala 93:22:@4628.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_31 RetimeWrapper_8 ( // @[package.scala 93:22:@4646.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_9 ( // @[package.scala 93:22:@4656.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_10 ( // @[package.scala 93:22:@4672.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_323 = RetimeWrapper_io_out; // @[package.scala 96:25:@4439.4 package.scala 96:25:@4440.4]
  assign _T_326 = ~ _T_323; // @[sm_x499_inr_Foreach.scala 70:18:@4442.4]
  assign _T_327 = ~ io_in_x475_fifo_active_0_out; // @[sm_x499_inr_Foreach.scala 70:45:@4443.4]
  assign _T_328 = _T_326 | _T_327; // @[sm_x499_inr_Foreach.scala 70:43:@4444.4]
  assign b479_number = __io_result; // @[Math.scala 723:22:@4428.4 Math.scala 724:14:@4429.4]
  assign _GEN_0 = {{1'd0}, b479_number}; // @[Math.scala 461:32:@4448.4]
  assign _T_331 = _GEN_0 << 1; // @[Math.scala 461:32:@4448.4]
  assign x739_sum_number = x739_sum_1_io_result; // @[Math.scala 154:22:@4458.4 Math.scala 155:14:@4459.4]
  assign _T_337 = x739_sum_number[31]; // @[FixedPoint.scala 50:25:@4463.4]
  assign _T_341 = _T_337 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@4465.4]
  assign _T_342 = x739_sum_number[31:4]; // @[FixedPoint.scala 18:52:@4466.4]
  assign _T_348 = _T_342 == 28'hfffffff; // @[Math.scala 451:55:@4468.4]
  assign _T_349 = x739_sum_number[3:0]; // @[FixedPoint.scala 18:52:@4469.4]
  assign _T_355 = _T_349 != 4'h0; // @[Math.scala 451:110:@4471.4]
  assign _T_356 = _T_348 & _T_355; // @[Math.scala 451:94:@4472.4]
  assign _T_358 = {_T_341,_T_342}; // @[Cat.scala 30:58:@4474.4]
  assign x482_1_number = _T_356 ? 32'h0 : _T_358; // @[Math.scala 454:20:@4475.4]
  assign _GEN_1 = {{4'd0}, x482_1_number}; // @[Math.scala 461:32:@4480.4]
  assign _T_363 = _GEN_1 << 4; // @[Math.scala 461:32:@4480.4]
  assign _GEN_2 = {{6'd0}, x482_1_number}; // @[Math.scala 461:32:@4485.4]
  assign _T_366 = _GEN_2 << 6; // @[Math.scala 461:32:@4485.4]
  assign x487_sum_number = x487_sum_1_io_result; // @[Math.scala 154:22:@4519.4 Math.scala 155:14:@4520.4]
  assign _T_386 = x487_sum_number[31]; // @[FixedPoint.scala 50:25:@4524.4]
  assign _T_390 = _T_386 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@4526.4]
  assign _T_391 = x487_sum_number[31:4]; // @[FixedPoint.scala 18:52:@4527.4]
  assign _T_397 = _T_391 == 28'hfffffff; // @[Math.scala 451:55:@4529.4]
  assign _T_398 = x487_sum_number[3:0]; // @[FixedPoint.scala 18:52:@4530.4]
  assign _T_404 = _T_398 != 4'h0; // @[Math.scala 451:110:@4532.4]
  assign _T_405 = _T_397 & _T_404; // @[Math.scala 451:94:@4533.4]
  assign _T_407 = {_T_390,_T_391}; // @[Cat.scala 30:58:@4535.4]
  assign x488_1_number = _T_405 ? 32'h0 : _T_407; // @[Math.scala 454:20:@4536.4]
  assign _GEN_3 = {{4'd0}, x488_1_number}; // @[Math.scala 461:32:@4541.4]
  assign _GEN_4 = {{6'd0}, x488_1_number}; // @[Math.scala 461:32:@4553.4]
  assign _T_419 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@4559.4 package.scala 96:25:@4560.4]
  assign x741_1_number = _T_419[31:0]; // @[Math.scala 459:22:@4552.4 Math.scala 461:14:@4561.4]
  assign x759_x493_sum_D1_number = RetimeWrapper_4_io_out; // @[package.scala 96:25:@4599.4 package.scala 96:25:@4600.4]
  assign x494_tuple = {1'h1,x741_1_number,x759_x493_sum_D1_number}; // @[Cat.scala 30:58:@4604.4]
  assign _T_454 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@4633.4 package.scala 96:25:@4634.4]
  assign _T_456 = io_rr ? _T_454 : 1'h0; // @[implicits.scala 56:10:@4635.4]
  assign x760_x495_D4 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@4613.4 package.scala 96:25:@4614.4]
  assign _T_457 = _T_456 & x760_x495_D4; // @[sm_x499_inr_Foreach.scala 108:121:@4636.4]
  assign x761_b480_D4 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@4623.4 package.scala 96:25:@4624.4]
  assign _T_458 = _T_457 & x761_b480_D4; // @[sm_x499_inr_Foreach.scala 108:127:@4637.4]
  assign x762_x486_sum_D1_number = RetimeWrapper_8_io_out; // @[package.scala 96:25:@4651.4 package.scala 96:25:@4652.4]
  assign x763_x485_sub_D2_number = RetimeWrapper_9_io_out; // @[package.scala 96:25:@4661.4 package.scala 96:25:@4662.4]
  assign _T_473 = {x762_x486_sum_D1_number,x763_x485_sub_D2_number}; // @[Cat.scala 30:58:@4665.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@4547.4 package.scala 96:25:@4548.4]
  assign x489_1_number = _T_414[31:0]; // @[Math.scala 459:22:@4540.4 Math.scala 461:14:@4549.4]
  assign _T_475 = ~ io_sigsIn_break; // @[sm_x499_inr_Foreach.scala 121:121:@4668.4]
  assign _T_481 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@4677.4 package.scala 96:25:@4678.4]
  assign _T_483 = io_rr ? _T_481 : 1'h0; // @[implicits.scala 56:10:@4679.4]
  assign _T_484 = _T_475 & _T_483; // @[sm_x499_inr_Foreach.scala 121:138:@4680.4]
  assign _T_486 = _T_484 & _T_475; // @[sm_x499_inr_Foreach.scala 121:235:@4682.4]
  assign _T_487 = _T_486 & io_sigsIn_backpressure; // @[sm_x499_inr_Foreach.scala 121:254:@4683.4]
  assign io_in_x475_fifo_wPort_0_data_0 = {_T_473,x489_1_number}; // @[MemInterfaceType.scala 90:56:@4686.4]
  assign io_in_x475_fifo_wPort_0_en_0 = _T_487 & x761_b480_D4; // @[MemInterfaceType.scala 93:57:@4688.4]
  assign io_in_x475_fifo_active_0_in = RetimeWrapper_6_io_out; // @[MemInterfaceType.scala 147:18:@4690.4]
  assign io_in_x474_valid = _T_458 & io_sigsIn_backpressure; // @[sm_x499_inr_Foreach.scala 108:18:@4639.4]
  assign io_in_x474_bits_addr = x494_tuple[63:0]; // @[sm_x499_inr_Foreach.scala 109:22:@4641.4]
  assign io_in_x474_bits_size = x494_tuple[95:64]; // @[sm_x499_inr_Foreach.scala 110:22:@4643.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@4426.4]
  assign RetimeWrapper_clock = clock; // @[:@4435.4]
  assign RetimeWrapper_reset = reset; // @[:@4436.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@4438.4]
  assign RetimeWrapper_io_in = io_in_x475_fifo_full; // @[package.scala 94:16:@4437.4]
  assign x739_sum_1_clock = clock; // @[:@4453.4]
  assign x739_sum_1_reset = reset; // @[:@4454.4]
  assign x739_sum_1_io_a = _T_331[31:0]; // @[Math.scala 151:17:@4455.4]
  assign x739_sum_1_io_b = __io_result; // @[Math.scala 152:17:@4456.4]
  assign x739_sum_1_io_flow = _T_328 & io_in_x474_ready; // @[Math.scala 153:20:@4457.4]
  assign x485_sub_1_clock = clock; // @[:@4490.4]
  assign x485_sub_1_reset = reset; // @[:@4491.4]
  assign x485_sub_1_io_a = x739_sum_1_io_result; // @[Math.scala 192:17:@4492.4]
  assign x485_sub_1_io_b = _T_363[31:0]; // @[Math.scala 193:17:@4493.4]
  assign x485_sub_1_io_flow = _T_328 & io_in_x474_ready; // @[Math.scala 194:20:@4494.4]
  assign x486_sum_1_clock = clock; // @[:@4502.4]
  assign x486_sum_1_reset = reset; // @[:@4503.4]
  assign x486_sum_1_io_a = x485_sub_1_io_result; // @[Math.scala 151:17:@4504.4]
  assign x486_sum_1_io_b = 32'h3; // @[Math.scala 152:17:@4505.4]
  assign x486_sum_1_io_flow = _T_328 & io_in_x474_ready; // @[Math.scala 153:20:@4506.4]
  assign x487_sum_1_clock = clock; // @[:@4514.4]
  assign x487_sum_1_reset = reset; // @[:@4515.4]
  assign x487_sum_1_io_a = x485_sub_1_io_result; // @[Math.scala 151:17:@4516.4]
  assign x487_sum_1_io_b = 32'h12; // @[Math.scala 152:17:@4517.4]
  assign x487_sum_1_io_flow = _T_328 & io_in_x474_ready; // @[Math.scala 153:20:@4518.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4543.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4544.4]
  assign RetimeWrapper_1_io_flow = _T_328 & io_in_x474_ready; // @[package.scala 95:18:@4546.4]
  assign RetimeWrapper_1_io_in = _GEN_3 << 4; // @[package.scala 94:16:@4545.4]
  assign RetimeWrapper_2_clock = clock; // @[:@4555.4]
  assign RetimeWrapper_2_reset = reset; // @[:@4556.4]
  assign RetimeWrapper_2_io_flow = _T_328 & io_in_x474_ready; // @[package.scala 95:18:@4558.4]
  assign RetimeWrapper_2_io_in = _GEN_4 << 6; // @[package.scala 94:16:@4557.4]
  assign x491_1_io_b = _T_366[31:0]; // @[Math.scala 721:17:@4567.4]
  assign RetimeWrapper_3_clock = clock; // @[:@4575.4]
  assign RetimeWrapper_3_reset = reset; // @[:@4576.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4578.4]
  assign RetimeWrapper_3_io_in = io_in_x468_A_dram_number; // @[package.scala 94:16:@4577.4]
  assign x493_sum_1_clock = clock; // @[:@4584.4]
  assign x493_sum_1_reset = reset; // @[:@4585.4]
  assign x493_sum_1_io_a = x491_1_io_result; // @[Math.scala 151:17:@4586.4]
  assign x493_sum_1_io_b = RetimeWrapper_3_io_out; // @[Math.scala 152:17:@4587.4]
  assign x493_sum_1_io_flow = _T_328 & io_in_x474_ready; // @[Math.scala 153:20:@4588.4]
  assign RetimeWrapper_4_clock = clock; // @[:@4595.4]
  assign RetimeWrapper_4_reset = reset; // @[:@4596.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4598.4]
  assign RetimeWrapper_4_io_in = x493_sum_1_io_result; // @[package.scala 94:16:@4597.4]
  assign RetimeWrapper_5_clock = clock; // @[:@4609.4]
  assign RetimeWrapper_5_reset = reset; // @[:@4610.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4612.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@4611.4]
  assign RetimeWrapper_6_clock = clock; // @[:@4619.4]
  assign RetimeWrapper_6_reset = reset; // @[:@4620.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4622.4]
  assign RetimeWrapper_6_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@4621.4]
  assign RetimeWrapper_7_clock = clock; // @[:@4629.4]
  assign RetimeWrapper_7_reset = reset; // @[:@4630.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4632.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_datapathEn & io_sigsIn_iiIssue; // @[package.scala 94:16:@4631.4]
  assign RetimeWrapper_8_clock = clock; // @[:@4647.4]
  assign RetimeWrapper_8_reset = reset; // @[:@4648.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4650.4]
  assign RetimeWrapper_8_io_in = x486_sum_1_io_result; // @[package.scala 94:16:@4649.4]
  assign RetimeWrapper_9_clock = clock; // @[:@4657.4]
  assign RetimeWrapper_9_reset = reset; // @[:@4658.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4660.4]
  assign RetimeWrapper_9_io_in = x485_sub_1_io_result; // @[package.scala 94:16:@4659.4]
  assign RetimeWrapper_10_clock = clock; // @[:@4673.4]
  assign RetimeWrapper_10_reset = reset; // @[:@4674.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4676.4]
  assign RetimeWrapper_10_io_in = io_sigsIn_datapathEn & io_sigsIn_iiIssue; // @[package.scala 94:16:@4675.4]
endmodule
module x537_outr_Foreach_sm( // @[:@5029.2]
  input   clock, // @[:@5030.4]
  input   reset, // @[:@5031.4]
  input   io_enable, // @[:@5032.4]
  output  io_done, // @[:@5032.4]
  input   io_ctrDone, // @[:@5032.4]
  output  io_ctrInc, // @[:@5032.4]
  output  io_ctrRst, // @[:@5032.4]
  input   io_parentAck, // @[:@5032.4]
  input   io_doneIn_0, // @[:@5032.4]
  input   io_doneIn_1, // @[:@5032.4]
  input   io_maskIn_0, // @[:@5032.4]
  input   io_maskIn_1, // @[:@5032.4]
  output  io_enableOut_0, // @[:@5032.4]
  output  io_enableOut_1, // @[:@5032.4]
  output  io_childAck_0, // @[:@5032.4]
  output  io_childAck_1 // @[:@5032.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@5035.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@5035.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@5035.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@5035.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@5035.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@5035.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@5038.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@5038.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@5038.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@5038.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@5038.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@5038.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@5041.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@5041.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@5041.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@5041.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@5041.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@5041.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@5044.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@5044.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@5044.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@5044.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@5044.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@5044.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@5073.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@5073.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@5073.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@5073.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@5073.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@5073.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@5076.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@5076.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@5076.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@5076.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@5076.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@5076.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@5105.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@5105.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@5105.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@5105.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@5105.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@5201.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@5201.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@5201.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@5201.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@5201.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@5218.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@5218.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@5218.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@5218.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@5218.4]
  wire  allDone; // @[Controllers.scala 80:47:@5047.4]
  wire  _T_77; // @[Controllers.scala 81:26:@5048.4]
  wire  finished; // @[Controllers.scala 81:37:@5049.4]
  wire  _T_134; // @[package.scala 96:25:@5110.4 package.scala 96:25:@5111.4]
  wire  _T_138; // @[Controllers.scala 125:45:@5113.4]
  wire  _T_139; // @[Controllers.scala 125:61:@5114.4]
  wire  _T_140; // @[Controllers.scala 125:87:@5115.4]
  wire  synchronize; // @[Controllers.scala 125:42:@5117.4]
  wire  _T_144; // @[Controllers.scala 128:33:@5119.4]
  wire  _T_146; // @[Controllers.scala 128:54:@5120.4]
  wire  _T_147; // @[Controllers.scala 128:52:@5121.4]
  wire  _T_148; // @[Controllers.scala 128:66:@5122.4]
  wire  _T_150; // @[Controllers.scala 128:98:@5124.4]
  wire  _T_151; // @[Controllers.scala 128:96:@5125.4]
  wire  _T_153; // @[Controllers.scala 128:123:@5126.4]
  wire  _T_156; // @[Controllers.scala 129:57:@5130.4]
  wire  _T_160; // @[Controllers.scala 130:52:@5134.4]
  wire  _T_161; // @[Controllers.scala 130:50:@5135.4]
  wire  _T_163; // @[Controllers.scala 130:69:@5136.4]
  wire  _T_164; // @[Controllers.scala 130:83:@5137.4]
  wire  _T_166; // @[Controllers.scala 130:66:@5139.4]
  wire  _T_169; // @[Controllers.scala 130:129:@5141.4]
  wire  _T_175; // @[Controllers.scala 135:80:@5148.4]
  wire  _T_176; // @[Controllers.scala 135:78:@5149.4]
  wire  _T_178; // @[Controllers.scala 135:105:@5150.4]
  wire  _T_179; // @[Controllers.scala 135:103:@5151.4]
  wire  _T_180; // @[Controllers.scala 135:119:@5152.4]
  wire  _T_182; // @[Controllers.scala 135:51:@5154.4]
  wire  _T_191; // @[Controllers.scala 137:79:@5163.4]
  wire  _T_192; // @[Controllers.scala 137:95:@5164.4]
  wire  _T_194; // @[Controllers.scala 137:52:@5166.4]
  wire  _T_205; // @[Controllers.scala 213:68:@5179.4]
  wire  _T_207; // @[Controllers.scala 213:90:@5181.4]
  wire  _T_208; // @[Controllers.scala 213:115:@5182.4]
  wire  _T_209; // @[Controllers.scala 213:132:@5183.4]
  wire  _T_210; // @[Controllers.scala 213:130:@5184.4]
  wire  _T_211; // @[Controllers.scala 213:156:@5185.4]
  wire  _T_213; // @[Controllers.scala 213:68:@5188.4]
  wire  _T_215; // @[Controllers.scala 213:90:@5190.4]
  wire  _T_216; // @[Controllers.scala 213:115:@5191.4]
  wire  _T_222; // @[package.scala 100:49:@5196.4]
  reg  _T_225; // @[package.scala 48:56:@5197.4]
  reg [31:0] _RAND_0;
  wire  _T_226; // @[package.scala 100:41:@5199.4]
  reg  _T_239; // @[package.scala 48:56:@5215.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@5035.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@5038.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@5041.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@5044.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@5073.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@5076.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@5105.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@5201.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@5218.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@5047.4]
  assign _T_77 = allDone | io_done; // @[Controllers.scala 81:26:@5048.4]
  assign finished = _T_77 | done_1_io_input_set; // @[Controllers.scala 81:37:@5049.4]
  assign _T_134 = RetimeWrapper_io_out; // @[package.scala 96:25:@5110.4 package.scala 96:25:@5111.4]
  assign _T_138 = io_maskIn_1 == 1'h0; // @[Controllers.scala 125:45:@5113.4]
  assign _T_139 = _T_138 & iterDone_1_io_output; // @[Controllers.scala 125:61:@5114.4]
  assign _T_140 = _T_139 & io_enable; // @[Controllers.scala 125:87:@5115.4]
  assign synchronize = _T_134 | _T_140; // @[Controllers.scala 125:42:@5117.4]
  assign _T_144 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@5119.4]
  assign _T_146 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@5120.4]
  assign _T_147 = _T_144 & _T_146; // @[Controllers.scala 128:52:@5121.4]
  assign _T_148 = _T_147 & io_enable; // @[Controllers.scala 128:66:@5122.4]
  assign _T_150 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@5124.4]
  assign _T_151 = _T_148 & _T_150; // @[Controllers.scala 128:96:@5125.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@5126.4]
  assign _T_156 = io_doneIn_0 | io_parentAck; // @[Controllers.scala 129:57:@5130.4]
  assign _T_160 = synchronize == 1'h0; // @[Controllers.scala 130:52:@5134.4]
  assign _T_161 = io_doneIn_0 & _T_160; // @[Controllers.scala 130:50:@5135.4]
  assign _T_163 = io_maskIn_0 == 1'h0; // @[Controllers.scala 130:69:@5136.4]
  assign _T_164 = _T_163 & io_enable; // @[Controllers.scala 130:83:@5137.4]
  assign _T_166 = _T_161 | _T_164; // @[Controllers.scala 130:66:@5139.4]
  assign _T_169 = finished == 1'h0; // @[Controllers.scala 130:129:@5141.4]
  assign _T_175 = ~ iterDone_1_io_output; // @[Controllers.scala 135:80:@5148.4]
  assign _T_176 = iterDone_0_io_output & _T_175; // @[Controllers.scala 135:78:@5149.4]
  assign _T_178 = io_doneIn_1 == 1'h0; // @[Controllers.scala 135:105:@5150.4]
  assign _T_179 = _T_176 & _T_178; // @[Controllers.scala 135:103:@5151.4]
  assign _T_180 = _T_179 & io_enable; // @[Controllers.scala 135:119:@5152.4]
  assign _T_182 = io_doneIn_0 | _T_180; // @[Controllers.scala 135:51:@5154.4]
  assign _T_191 = iterDone_0_io_output & _T_138; // @[Controllers.scala 137:79:@5163.4]
  assign _T_192 = _T_191 & io_enable; // @[Controllers.scala 137:95:@5164.4]
  assign _T_194 = io_doneIn_1 | _T_192; // @[Controllers.scala 137:52:@5166.4]
  assign _T_205 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@5179.4]
  assign _T_207 = _T_205 & _T_150; // @[Controllers.scala 213:90:@5181.4]
  assign _T_208 = _T_207 & io_maskIn_0; // @[Controllers.scala 213:115:@5182.4]
  assign _T_209 = ~ allDone; // @[Controllers.scala 213:132:@5183.4]
  assign _T_210 = _T_208 & _T_209; // @[Controllers.scala 213:130:@5184.4]
  assign _T_211 = ~ io_ctrDone; // @[Controllers.scala 213:156:@5185.4]
  assign _T_213 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@5188.4]
  assign _T_215 = _T_213 & _T_175; // @[Controllers.scala 213:90:@5190.4]
  assign _T_216 = _T_215 & io_maskIn_1; // @[Controllers.scala 213:115:@5191.4]
  assign _T_222 = allDone == 1'h0; // @[package.scala 100:49:@5196.4]
  assign _T_226 = allDone & _T_225; // @[package.scala 100:41:@5199.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@5225.4]
  assign io_ctrInc = io_doneIn_1 | _T_140; // @[Controllers.scala 122:17:@5104.4]
  assign io_ctrRst = RetimeWrapper_1_io_out; // @[Controllers.scala 215:13:@5208.4]
  assign io_enableOut_0 = _T_210 & _T_211; // @[Controllers.scala 213:55:@5187.4]
  assign io_enableOut_1 = _T_216 & _T_209; // @[Controllers.scala 213:55:@5195.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@5176.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@5178.4]
  assign active_0_clock = clock; // @[:@5036.4]
  assign active_0_reset = reset; // @[:@5037.4]
  assign active_0_io_input_set = _T_151 & _T_153; // @[Controllers.scala 128:30:@5128.4]
  assign active_0_io_input_reset = _T_156 | allDone; // @[Controllers.scala 129:32:@5133.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@5050.4]
  assign active_1_clock = clock; // @[:@5039.4]
  assign active_1_reset = reset; // @[:@5040.4]
  assign active_1_io_input_set = _T_182 & _T_160; // @[Controllers.scala 135:32:@5157.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 136:34:@5161.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@5051.4]
  assign done_0_clock = clock; // @[:@5042.4]
  assign done_0_reset = reset; // @[:@5043.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 131:28:@5147.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@5062.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@5052.4]
  assign done_1_clock = clock; // @[:@5045.4]
  assign done_1_reset = reset; // @[:@5046.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 138:30:@5174.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@5071.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@5053.4]
  assign iterDone_0_clock = clock; // @[:@5074.4]
  assign iterDone_0_reset = reset; // @[:@5075.4]
  assign iterDone_0_io_input_set = _T_166 & _T_169; // @[Controllers.scala 130:32:@5143.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@5089.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@5079.4]
  assign iterDone_1_clock = clock; // @[:@5077.4]
  assign iterDone_1_reset = reset; // @[:@5078.4]
  assign iterDone_1_io_input_set = _T_194 & _T_160; // @[Controllers.scala 137:34:@5170.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@5098.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@5080.4]
  assign RetimeWrapper_clock = clock; // @[:@5106.4]
  assign RetimeWrapper_reset = reset; // @[:@5107.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@5109.4]
  assign RetimeWrapper_io_in = io_doneIn_1; // @[package.scala 94:16:@5108.4]
  assign RetimeWrapper_1_clock = clock; // @[:@5202.4]
  assign RetimeWrapper_1_reset = reset; // @[:@5203.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@5205.4]
  assign RetimeWrapper_1_io_in = _T_226 | io_parentAck; // @[package.scala 94:16:@5204.4]
  assign RetimeWrapper_2_clock = clock; // @[:@5219.4]
  assign RetimeWrapper_2_reset = reset; // @[:@5220.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@5222.4]
  assign RetimeWrapper_2_io_in = allDone & _T_239; // @[package.scala 94:16:@5221.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_225 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_239 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_225 <= 1'h0;
    end else begin
      _T_225 <= _T_222;
    end
    if (reset) begin
      _T_239 <= 1'h0;
    end else begin
      _T_239 <= _T_222;
    end
  end
endmodule
module x505_reg( // @[:@5376.2]
  input         clock, // @[:@5377.4]
  input         reset, // @[:@5378.4]
  output [31:0] io_rPort_0_output_0, // @[:@5379.4]
  input  [31:0] io_wPort_0_data_0, // @[:@5379.4]
  input         io_wPort_0_reset, // @[:@5379.4]
  input         io_wPort_0_en_0 // @[:@5379.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@5395.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 325:32:@5397.4]
  wire [31:0] _T_70; // @[MemPrimitives.scala 325:12:@5398.4]
  assign _T_69 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@5397.4]
  assign _T_70 = io_wPort_0_reset ? 32'h0 : _T_69; // @[MemPrimitives.scala 325:12:@5398.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@5400.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module x516_inr_UnitPipe_sm( // @[:@5608.2]
  input   clock, // @[:@5609.4]
  input   reset, // @[:@5610.4]
  input   io_enable, // @[:@5611.4]
  output  io_done, // @[:@5611.4]
  output  io_doneLatch, // @[:@5611.4]
  input   io_ctrDone, // @[:@5611.4]
  output  io_datapathEn, // @[:@5611.4]
  output  io_ctrInc, // @[:@5611.4]
  input   io_parentAck, // @[:@5611.4]
  input   io_backpressure, // @[:@5611.4]
  input   io_break // @[:@5611.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@5613.4]
  wire  active_reset; // @[Controllers.scala 261:22:@5613.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@5613.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@5613.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@5613.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@5613.4]
  wire  done_clock; // @[Controllers.scala 262:20:@5616.4]
  wire  done_reset; // @[Controllers.scala 262:20:@5616.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@5616.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@5616.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@5616.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@5616.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@5650.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@5650.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@5650.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@5650.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@5650.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@5672.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@5672.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@5672.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@5672.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@5672.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@5684.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@5684.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@5684.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@5684.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@5684.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@5692.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@5692.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@5692.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@5692.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@5692.4]
  wire  _T_80; // @[Controllers.scala 264:48:@5621.4]
  wire  _T_81; // @[Controllers.scala 264:46:@5622.4]
  wire  _T_82; // @[Controllers.scala 264:62:@5623.4]
  wire  _T_100; // @[package.scala 100:49:@5641.4]
  reg  _T_103; // @[package.scala 48:56:@5642.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@5665.4]
  wire  _T_124; // @[package.scala 96:25:@5677.4 package.scala 96:25:@5678.4]
  wire  _T_126; // @[package.scala 100:49:@5679.4]
  reg  _T_129; // @[package.scala 48:56:@5680.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@5702.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@5704.4]
  reg  _T_153; // @[package.scala 48:56:@5705.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@5707.4]
  wire  _T_156; // @[Controllers.scala 292:61:@5708.4]
  wire  _T_157; // @[Controllers.scala 292:24:@5709.4]
  SRFF active ( // @[Controllers.scala 261:22:@5613.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@5616.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@5650.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@5672.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@5684.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@5692.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@5621.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@5622.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@5623.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@5641.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@5665.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@5677.4 package.scala 96:25:@5678.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@5679.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@5704.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@5707.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@5708.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@5709.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@5683.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@5711.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@5668.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@5671.4]
  assign active_clock = clock; // @[:@5614.4]
  assign active_reset = reset; // @[:@5615.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@5626.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@5630.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@5631.4]
  assign done_clock = clock; // @[:@5617.4]
  assign done_reset = reset; // @[:@5618.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@5646.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@5639.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@5640.4]
  assign RetimeWrapper_clock = clock; // @[:@5651.4]
  assign RetimeWrapper_reset = reset; // @[:@5652.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@5654.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@5653.4]
  assign RetimeWrapper_1_clock = clock; // @[:@5673.4]
  assign RetimeWrapper_1_reset = reset; // @[:@5674.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@5676.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@5675.4]
  assign RetimeWrapper_2_clock = clock; // @[:@5685.4]
  assign RetimeWrapper_2_reset = reset; // @[:@5686.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@5688.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@5687.4]
  assign RetimeWrapper_3_clock = clock; // @[:@5693.4]
  assign RetimeWrapper_3_reset = reset; // @[:@5694.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@5696.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@5695.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1( // @[:@5786.2]
  output        io_in_x475_fifo_rPort_0_en_0, // @[:@5789.4]
  input  [95:0] io_in_x475_fifo_rPort_0_output_0, // @[:@5789.4]
  output [31:0] io_in_x507_reg_wPort_0_data_0, // @[:@5789.4]
  output        io_in_x507_reg_wPort_0_reset, // @[:@5789.4]
  output        io_in_x507_reg_wPort_0_en_0, // @[:@5789.4]
  output        io_in_x507_reg_reset, // @[:@5789.4]
  output [31:0] io_in_x505_reg_wPort_0_data_0, // @[:@5789.4]
  output        io_in_x505_reg_wPort_0_reset, // @[:@5789.4]
  output        io_in_x505_reg_wPort_0_en_0, // @[:@5789.4]
  output        io_in_x505_reg_reset, // @[:@5789.4]
  output [31:0] io_in_x506_reg_wPort_0_data_0, // @[:@5789.4]
  output        io_in_x506_reg_wPort_0_reset, // @[:@5789.4]
  output        io_in_x506_reg_wPort_0_en_0, // @[:@5789.4]
  output        io_in_x506_reg_reset, // @[:@5789.4]
  input         io_sigsIn_forwardpressure, // @[:@5789.4]
  input         io_sigsIn_datapathEn, // @[:@5789.4]
  input         io_sigsIn_break, // @[:@5789.4]
  input         io_rr // @[:@5789.4]
);
  wire  _T_692; // @[implicits.scala 56:10:@5862.4]
  wire  _T_693; // @[sm_x516_inr_UnitPipe.scala 78:120:@5863.4]
  wire  _T_694; // @[sm_x516_inr_UnitPipe.scala 78:117:@5864.4]
  wire  _T_699; // @[implicits.scala 56:10:@5867.4]
  wire  _T_714; // @[sm_x516_inr_UnitPipe.scala 90:133:@5885.4]
  assign _T_692 = io_rr ? io_sigsIn_forwardpressure : 1'h0; // @[implicits.scala 56:10:@5862.4]
  assign _T_693 = ~ io_sigsIn_break; // @[sm_x516_inr_UnitPipe.scala 78:120:@5863.4]
  assign _T_694 = _T_692 & _T_693; // @[sm_x516_inr_UnitPipe.scala 78:117:@5864.4]
  assign _T_699 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 56:10:@5867.4]
  assign _T_714 = _T_693 & _T_699; // @[sm_x516_inr_UnitPipe.scala 90:133:@5885.4]
  assign io_in_x475_fifo_rPort_0_en_0 = _T_694 & _T_699; // @[MemInterfaceType.scala 110:79:@5872.4]
  assign io_in_x507_reg_wPort_0_data_0 = io_in_x475_fifo_rPort_0_output_0[31:0]; // @[MemInterfaceType.scala 90:56:@5922.4]
  assign io_in_x507_reg_wPort_0_reset = io_in_x507_reg_reset; // @[MemInterfaceType.scala 91:23:@5923.4]
  assign io_in_x507_reg_wPort_0_en_0 = _T_714 & _T_693; // @[MemInterfaceType.scala 93:57:@5924.4]
  assign io_in_x507_reg_reset = 1'h0;
  assign io_in_x505_reg_wPort_0_data_0 = io_in_x475_fifo_rPort_0_output_0[63:32]; // @[MemInterfaceType.scala 90:56:@5890.4]
  assign io_in_x505_reg_wPort_0_reset = io_in_x505_reg_reset; // @[MemInterfaceType.scala 91:23:@5891.4]
  assign io_in_x505_reg_wPort_0_en_0 = _T_714 & _T_693; // @[MemInterfaceType.scala 93:57:@5892.4]
  assign io_in_x505_reg_reset = 1'h0;
  assign io_in_x506_reg_wPort_0_data_0 = io_in_x475_fifo_rPort_0_output_0[95:64]; // @[MemInterfaceType.scala 90:56:@5906.4]
  assign io_in_x506_reg_wPort_0_reset = io_in_x506_reg_reset; // @[MemInterfaceType.scala 91:23:@5907.4]
  assign io_in_x506_reg_wPort_0_en_0 = _T_714 & _T_693; // @[MemInterfaceType.scala 93:57:@5908.4]
  assign io_in_x506_reg_reset = 1'h0;
endmodule
module SingleCounter_3( // @[:@5964.2]
  input         clock, // @[:@5965.4]
  input         reset, // @[:@5966.4]
  input  [31:0] io_setup_stop, // @[:@5967.4]
  input         io_setup_saturate, // @[:@5967.4]
  input         io_input_reset, // @[:@5967.4]
  input         io_input_enable, // @[:@5967.4]
  output [31:0] io_output_count_0, // @[:@5967.4]
  output        io_output_oobs_0, // @[:@5967.4]
  output        io_output_noop, // @[:@5967.4]
  output        io_output_done // @[:@5967.4]
);
  wire  bases_0_clock; // @[Counter.scala 262:53:@5980.4]
  wire  bases_0_reset; // @[Counter.scala 262:53:@5980.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 262:53:@5980.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 262:53:@5980.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 262:53:@5980.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 262:53:@5980.4]
  wire  SRFF_clock; // @[Counter.scala 264:22:@5996.4]
  wire  SRFF_reset; // @[Counter.scala 264:22:@5996.4]
  wire  SRFF_io_input_set; // @[Counter.scala 264:22:@5996.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 264:22:@5996.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 264:22:@5996.4]
  wire  SRFF_io_output; // @[Counter.scala 264:22:@5996.4]
  wire  _T_36; // @[Counter.scala 265:45:@5999.4]
  wire [31:0] _T_48; // @[Counter.scala 288:52:@6024.4]
  wire [32:0] _T_50; // @[Counter.scala 292:33:@6025.4]
  wire [31:0] _T_51; // @[Counter.scala 292:33:@6026.4]
  wire [31:0] _T_52; // @[Counter.scala 292:33:@6027.4]
  wire  _T_56; // @[Counter.scala 294:18:@6029.4]
  wire [31:0] _T_66; // @[Counter.scala 300:115:@6037.4]
  wire [31:0] _T_68; // @[Counter.scala 300:85:@6039.4]
  wire [31:0] _T_69; // @[Counter.scala 300:152:@6040.4]
  wire [31:0] _T_70; // @[Counter.scala 300:74:@6041.4]
  wire  _T_73; // @[Counter.scala 325:102:@6045.4]
  wire  _T_74; // @[Counter.scala 325:130:@6046.4]
  FF bases_0 ( // @[Counter.scala 262:53:@5980.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 264:22:@5996.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 265:45:@5999.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 288:52:@6024.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 292:33:@6025.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 292:33:@6026.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 292:33:@6027.4]
  assign _T_56 = $signed(_T_52) >= $signed(io_setup_stop); // @[Counter.scala 294:18:@6029.4]
  assign _T_66 = $unsigned(_T_48); // @[Counter.scala 300:115:@6037.4]
  assign _T_68 = io_setup_saturate ? _T_66 : 32'h0; // @[Counter.scala 300:85:@6039.4]
  assign _T_69 = $unsigned(_T_52); // @[Counter.scala 300:152:@6040.4]
  assign _T_70 = _T_56 ? _T_68 : _T_69; // @[Counter.scala 300:74:@6041.4]
  assign _T_73 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 325:102:@6045.4]
  assign _T_74 = $signed(_T_48) >= $signed(io_setup_stop); // @[Counter.scala 325:130:@6046.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 305:28:@6044.4]
  assign io_output_oobs_0 = _T_73 | _T_74; // @[Counter.scala 325:60:@6048.4]
  assign io_output_noop = $signed(32'sh0) == $signed(io_setup_stop); // @[Counter.scala 337:40:@6052.4]
  assign io_output_done = io_input_enable & _T_56; // @[Counter.scala 334:20:@6050.4]
  assign bases_0_clock = clock; // @[:@5981.4]
  assign bases_0_reset = reset; // @[:@5982.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_70; // @[Counter.scala 300:31:@6043.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 282:27:@6022.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 285:29:@6023.4]
  assign SRFF_clock = clock; // @[:@5997.4]
  assign SRFF_reset = reset; // @[:@5998.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 265:23:@6001.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 266:25:@6003.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 267:30:@6004.4]
endmodule
module x519_ctrchain( // @[:@6056.2]
  input         clock, // @[:@6057.4]
  input         reset, // @[:@6058.4]
  input  [31:0] io_setup_stops_0, // @[:@6059.4]
  input         io_input_reset, // @[:@6059.4]
  input         io_input_enable, // @[:@6059.4]
  output [31:0] io_output_counts_0, // @[:@6059.4]
  output        io_output_oobs_0, // @[:@6059.4]
  output        io_output_noop, // @[:@6059.4]
  output        io_output_done // @[:@6059.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 514:46:@6061.4]
  wire  ctrs_0_reset; // @[Counter.scala 514:46:@6061.4]
  wire [31:0] ctrs_0_io_setup_stop; // @[Counter.scala 514:46:@6061.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 514:46:@6061.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 514:46:@6061.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 514:46:@6061.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 514:46:@6061.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 514:46:@6061.4]
  wire  ctrs_0_io_output_noop; // @[Counter.scala 514:46:@6061.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 514:46:@6061.4]
  reg  wasDone; // @[Counter.scala 543:24:@6070.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 547:69:@6076.4]
  wire  _T_47; // @[Counter.scala 547:80:@6077.4]
  reg  doneLatch; // @[Counter.scala 551:26:@6082.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 552:48:@6083.4]
  wire  _T_55; // @[Counter.scala 552:19:@6084.4]
  SingleCounter_3 ctrs_0 ( // @[Counter.scala 514:46:@6061.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_stop(ctrs_0_io_setup_stop),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_noop(ctrs_0_io_output_noop),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 547:69:@6076.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 547:80:@6077.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 552:48:@6083.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 552:19:@6084.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 558:32:@6086.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 559:30:@6088.4]
  assign io_output_noop = ctrs_0_io_output_noop; // @[Counter.scala 546:18:@6074.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 547:18:@6079.4]
  assign ctrs_0_clock = clock; // @[:@6062.4]
  assign ctrs_0_reset = reset; // @[:@6063.4]
  assign ctrs_0_io_setup_stop = io_setup_stops_0; // @[Counter.scala 519:23:@6065.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 531:29:@6069.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 521:24:@6067.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 525:33:@6068.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_58( // @[:@6128.2]
  input   clock, // @[:@6129.4]
  input   reset, // @[:@6130.4]
  input   io_flow, // @[:@6131.4]
  input   io_in, // @[:@6131.4]
  output  io_out // @[:@6131.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6133.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6133.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6133.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6133.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6133.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6133.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@6133.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6146.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6145.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6144.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6143.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6142.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6140.4]
endmodule
module x536_inr_Foreach_sm( // @[:@6276.2]
  input   clock, // @[:@6277.4]
  input   reset, // @[:@6278.4]
  input   io_enable, // @[:@6279.4]
  output  io_done, // @[:@6279.4]
  output  io_doneLatch, // @[:@6279.4]
  input   io_ctrDone, // @[:@6279.4]
  output  io_datapathEn, // @[:@6279.4]
  output  io_ctrInc, // @[:@6279.4]
  output  io_ctrRst, // @[:@6279.4]
  input   io_parentAck, // @[:@6279.4]
  input   io_backpressure, // @[:@6279.4]
  input   io_break // @[:@6279.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@6281.4]
  wire  active_reset; // @[Controllers.scala 261:22:@6281.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@6281.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@6281.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@6281.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@6281.4]
  wire  done_clock; // @[Controllers.scala 262:20:@6284.4]
  wire  done_reset; // @[Controllers.scala 262:20:@6284.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@6284.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@6284.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@6284.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@6284.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6318.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6318.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6318.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6318.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6318.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6340.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6340.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6340.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6340.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6340.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6352.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6352.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6352.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6352.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6352.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6360.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6360.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6360.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6360.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6360.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@6376.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@6376.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@6376.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@6376.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@6376.4]
  wire  _T_80; // @[Controllers.scala 264:48:@6289.4]
  wire  _T_81; // @[Controllers.scala 264:46:@6290.4]
  wire  _T_82; // @[Controllers.scala 264:62:@6291.4]
  wire  _T_100; // @[package.scala 100:49:@6309.4]
  reg  _T_103; // @[package.scala 48:56:@6310.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@6323.4 package.scala 96:25:@6324.4]
  wire  _T_110; // @[package.scala 100:49:@6325.4]
  reg  _T_113; // @[package.scala 48:56:@6326.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@6328.4]
  wire  _T_118; // @[Controllers.scala 283:41:@6333.4]
  wire  _T_124; // @[package.scala 96:25:@6345.4 package.scala 96:25:@6346.4]
  wire  _T_126; // @[package.scala 100:49:@6347.4]
  reg  _T_129; // @[package.scala 48:56:@6348.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@6370.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@6372.4]
  reg  _T_153; // @[package.scala 48:56:@6373.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@6381.4 package.scala 96:25:@6382.4]
  wire  _T_158; // @[Controllers.scala 292:61:@6383.4]
  wire  _T_159; // @[Controllers.scala 292:24:@6384.4]
  SRFF active ( // @[Controllers.scala 261:22:@6281.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@6284.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_58 RetimeWrapper ( // @[package.scala 93:22:@6318.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_58 RetimeWrapper_1 ( // @[package.scala 93:22:@6340.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6352.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6360.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@6376.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@6289.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@6290.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@6291.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@6309.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@6323.4 package.scala 96:25:@6324.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@6325.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@6328.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@6333.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6345.4 package.scala 96:25:@6346.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@6347.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@6372.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@6381.4 package.scala 96:25:@6382.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@6383.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@6384.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@6351.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@6386.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@6336.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@6339.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@6331.4]
  assign active_clock = clock; // @[:@6282.4]
  assign active_reset = reset; // @[:@6283.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@6294.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@6298.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@6299.4]
  assign done_clock = clock; // @[:@6285.4]
  assign done_reset = reset; // @[:@6286.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@6314.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@6307.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@6308.4]
  assign RetimeWrapper_clock = clock; // @[:@6319.4]
  assign RetimeWrapper_reset = reset; // @[:@6320.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@6322.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@6321.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6341.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6342.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@6344.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@6343.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6353.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6354.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6356.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@6355.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6361.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6362.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6364.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@6363.4]
  assign RetimeWrapper_4_clock = clock; // @[:@6377.4]
  assign RetimeWrapper_4_reset = reset; // @[:@6378.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@6380.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@6379.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x536_inr_Foreach_kernelx536_inr_Foreach_concrete1( // @[:@7323.2]
  input         clock, // @[:@7324.4]
  input         reset, // @[:@7325.4]
  output [8:0]  io_in_x472_A_sram_1_wPort_0_ofs_0, // @[:@7326.4]
  output [31:0] io_in_x472_A_sram_1_wPort_0_data_0, // @[:@7326.4]
  output        io_in_x472_A_sram_1_wPort_0_en_0, // @[:@7326.4]
  input         io_in_b504, // @[:@7326.4]
  output [8:0]  io_in_x471_A_sram_0_wPort_0_ofs_0, // @[:@7326.4]
  output [31:0] io_in_x471_A_sram_0_wPort_0_data_0, // @[:@7326.4]
  output        io_in_x471_A_sram_0_wPort_0_en_0, // @[:@7326.4]
  output        io_in_x476_ready, // @[:@7326.4]
  input  [31:0] io_in_x476_bits_rdata_0, // @[:@7326.4]
  input  [31:0] io_in_b503_number, // @[:@7326.4]
  input  [31:0] io_in_x505_reg_rPort_0_output_0, // @[:@7326.4]
  output [8:0]  io_in_x473_A_sram_2_wPort_0_ofs_0, // @[:@7326.4]
  output [31:0] io_in_x473_A_sram_2_wPort_0_data_0, // @[:@7326.4]
  output        io_in_x473_A_sram_2_wPort_0_en_0, // @[:@7326.4]
  input  [31:0] io_in_x506_reg_rPort_0_output_0, // @[:@7326.4]
  input         io_sigsIn_datapathEn, // @[:@7326.4]
  input         io_sigsIn_break, // @[:@7326.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@7326.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@7326.4]
  input         io_rr // @[:@7326.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@7405.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@7405.4]
  wire  x527_sub_1_clock; // @[Math.scala 191:24:@7456.4]
  wire  x527_sub_1_reset; // @[Math.scala 191:24:@7456.4]
  wire [31:0] x527_sub_1_io_a; // @[Math.scala 191:24:@7456.4]
  wire [31:0] x527_sub_1_io_b; // @[Math.scala 191:24:@7456.4]
  wire  x527_sub_1_io_flow; // @[Math.scala 191:24:@7456.4]
  wire [31:0] x527_sub_1_io_result; // @[Math.scala 191:24:@7456.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@7472.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@7472.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@7472.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@7472.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@7472.4]
  wire  x743_sum_1_clock; // @[Math.scala 150:24:@7488.4]
  wire  x743_sum_1_reset; // @[Math.scala 150:24:@7488.4]
  wire [31:0] x743_sum_1_io_a; // @[Math.scala 150:24:@7488.4]
  wire [31:0] x743_sum_1_io_b; // @[Math.scala 150:24:@7488.4]
  wire  x743_sum_1_io_flow; // @[Math.scala 150:24:@7488.4]
  wire [31:0] x743_sum_1_io_result; // @[Math.scala 150:24:@7488.4]
  wire  x532_sum_1_clock; // @[Math.scala 150:24:@7498.4]
  wire  x532_sum_1_reset; // @[Math.scala 150:24:@7498.4]
  wire [31:0] x532_sum_1_io_a; // @[Math.scala 150:24:@7498.4]
  wire [31:0] x532_sum_1_io_b; // @[Math.scala 150:24:@7498.4]
  wire  x532_sum_1_io_flow; // @[Math.scala 150:24:@7498.4]
  wire [31:0] x532_sum_1_io_result; // @[Math.scala 150:24:@7498.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@7509.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@7509.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@7509.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@7509.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@7509.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@7519.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@7519.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@7519.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@7519.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@7519.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@7529.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@7529.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@7529.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@7529.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@7529.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@7539.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@7539.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@7539.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@7539.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@7539.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@7553.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@7553.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@7553.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@7553.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@7553.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@7579.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@7579.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@7579.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@7579.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@7579.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@7605.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@7605.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@7605.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@7605.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@7605.4]
  wire  b521; // @[sm_x536_inr_Foreach.scala 88:18:@7413.4]
  wire  _T_787; // @[sm_x536_inr_Foreach.scala 93:119:@7417.4]
  wire [31:0] _T_799; // @[Math.scala 493:37:@7429.4]
  wire [31:0] b520_number; // @[Math.scala 723:22:@7410.4 Math.scala 724:14:@7411.4]
  wire [31:0] _T_800; // @[Math.scala 493:51:@7430.4]
  wire  x523; // @[Math.scala 493:44:@7431.4]
  wire [31:0] _T_820; // @[Math.scala 476:50:@7449.4]
  wire  x525; // @[Math.scala 476:44:@7450.4]
  wire  _T_834; // @[sm_x536_inr_Foreach.scala 110:26:@7466.4]
  wire [32:0] _GEN_0; // @[Math.scala 461:32:@7484.4]
  wire [32:0] _T_850; // @[Math.scala 461:32:@7484.4]
  wire  _T_889; // @[package.scala 96:25:@7558.4 package.scala 96:25:@7559.4]
  wire  _T_891; // @[implicits.scala 56:10:@7560.4]
  wire  _T_892; // @[sm_x536_inr_Foreach.scala 135:118:@7561.4]
  wire  _T_894; // @[sm_x536_inr_Foreach.scala 135:215:@7563.4]
  wire  x767_x526_D2; // @[package.scala 96:25:@7534.4 package.scala 96:25:@7535.4]
  wire  _T_896; // @[sm_x536_inr_Foreach.scala 135:260:@7565.4]
  wire  x768_b521_D2; // @[package.scala 96:25:@7544.4 package.scala 96:25:@7545.4]
  wire  _T_897; // @[sm_x536_inr_Foreach.scala 135:268:@7566.4]
  wire  x765_b504_D2; // @[package.scala 96:25:@7514.4 package.scala 96:25:@7515.4]
  wire  _T_909; // @[package.scala 96:25:@7584.4 package.scala 96:25:@7585.4]
  wire  _T_911; // @[implicits.scala 56:10:@7586.4]
  wire  _T_912; // @[sm_x536_inr_Foreach.scala 140:118:@7587.4]
  wire  _T_914; // @[sm_x536_inr_Foreach.scala 140:215:@7589.4]
  wire  _T_916; // @[sm_x536_inr_Foreach.scala 140:260:@7591.4]
  wire  _T_917; // @[sm_x536_inr_Foreach.scala 140:268:@7592.4]
  wire  _T_929; // @[package.scala 96:25:@7610.4 package.scala 96:25:@7611.4]
  wire  _T_931; // @[implicits.scala 56:10:@7612.4]
  wire  _T_932; // @[sm_x536_inr_Foreach.scala 145:118:@7613.4]
  wire  _T_934; // @[sm_x536_inr_Foreach.scala 145:215:@7615.4]
  wire  _T_936; // @[sm_x536_inr_Foreach.scala 145:260:@7617.4]
  wire  _T_937; // @[sm_x536_inr_Foreach.scala 145:268:@7618.4]
  wire [31:0] x532_sum_number; // @[Math.scala 154:22:@7504.4 Math.scala 155:14:@7505.4]
  _ _ ( // @[Math.scala 720:24:@7405.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x485_sub x527_sub_1 ( // @[Math.scala 191:24:@7456.4]
    .clock(x527_sub_1_clock),
    .reset(x527_sub_1_reset),
    .io_a(x527_sub_1_io_a),
    .io_b(x527_sub_1_io_b),
    .io_flow(x527_sub_1_io_flow),
    .io_result(x527_sub_1_io_result)
  );
  RetimeWrapper_31 RetimeWrapper ( // @[package.scala 93:22:@7472.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x739_sum x743_sum_1 ( // @[Math.scala 150:24:@7488.4]
    .clock(x743_sum_1_clock),
    .reset(x743_sum_1_reset),
    .io_a(x743_sum_1_io_a),
    .io_b(x743_sum_1_io_b),
    .io_flow(x743_sum_1_io_flow),
    .io_result(x743_sum_1_io_result)
  );
  x739_sum x532_sum_1 ( // @[Math.scala 150:24:@7498.4]
    .clock(x532_sum_1_clock),
    .reset(x532_sum_1_reset),
    .io_a(x532_sum_1_io_a),
    .io_b(x532_sum_1_io_b),
    .io_flow(x532_sum_1_io_flow),
    .io_result(x532_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@7509.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_31 RetimeWrapper_2 ( // @[package.scala 93:22:@7519.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@7529.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@7539.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@7553.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@7579.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@7605.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign b521 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x536_inr_Foreach.scala 88:18:@7413.4]
  assign _T_787 = ~ io_sigsIn_break; // @[sm_x536_inr_Foreach.scala 93:119:@7417.4]
  assign _T_799 = $signed(io_in_x505_reg_rPort_0_output_0); // @[Math.scala 493:37:@7429.4]
  assign b520_number = __io_result; // @[Math.scala 723:22:@7410.4 Math.scala 724:14:@7411.4]
  assign _T_800 = $signed(b520_number); // @[Math.scala 493:51:@7430.4]
  assign x523 = $signed(_T_799) <= $signed(_T_800); // @[Math.scala 493:44:@7431.4]
  assign _T_820 = $signed(io_in_x506_reg_rPort_0_output_0); // @[Math.scala 476:50:@7449.4]
  assign x525 = $signed(_T_800) < $signed(_T_820); // @[Math.scala 476:44:@7450.4]
  assign _T_834 = b521 & io_in_b504; // @[sm_x536_inr_Foreach.scala 110:26:@7466.4]
  assign _GEN_0 = {{1'd0}, io_in_b503_number}; // @[Math.scala 461:32:@7484.4]
  assign _T_850 = _GEN_0 << 1; // @[Math.scala 461:32:@7484.4]
  assign _T_889 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@7558.4 package.scala 96:25:@7559.4]
  assign _T_891 = io_rr ? _T_889 : 1'h0; // @[implicits.scala 56:10:@7560.4]
  assign _T_892 = _T_787 & _T_891; // @[sm_x536_inr_Foreach.scala 135:118:@7561.4]
  assign _T_894 = _T_892 & _T_787; // @[sm_x536_inr_Foreach.scala 135:215:@7563.4]
  assign x767_x526_D2 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@7534.4 package.scala 96:25:@7535.4]
  assign _T_896 = _T_894 & x767_x526_D2; // @[sm_x536_inr_Foreach.scala 135:260:@7565.4]
  assign x768_b521_D2 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@7544.4 package.scala 96:25:@7545.4]
  assign _T_897 = _T_896 & x768_b521_D2; // @[sm_x536_inr_Foreach.scala 135:268:@7566.4]
  assign x765_b504_D2 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@7514.4 package.scala 96:25:@7515.4]
  assign _T_909 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@7584.4 package.scala 96:25:@7585.4]
  assign _T_911 = io_rr ? _T_909 : 1'h0; // @[implicits.scala 56:10:@7586.4]
  assign _T_912 = _T_787 & _T_911; // @[sm_x536_inr_Foreach.scala 140:118:@7587.4]
  assign _T_914 = _T_912 & _T_787; // @[sm_x536_inr_Foreach.scala 140:215:@7589.4]
  assign _T_916 = _T_914 & x767_x526_D2; // @[sm_x536_inr_Foreach.scala 140:260:@7591.4]
  assign _T_917 = _T_916 & x768_b521_D2; // @[sm_x536_inr_Foreach.scala 140:268:@7592.4]
  assign _T_929 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@7610.4 package.scala 96:25:@7611.4]
  assign _T_931 = io_rr ? _T_929 : 1'h0; // @[implicits.scala 56:10:@7612.4]
  assign _T_932 = _T_787 & _T_931; // @[sm_x536_inr_Foreach.scala 145:118:@7613.4]
  assign _T_934 = _T_932 & _T_787; // @[sm_x536_inr_Foreach.scala 145:215:@7615.4]
  assign _T_936 = _T_934 & x767_x526_D2; // @[sm_x536_inr_Foreach.scala 145:260:@7617.4]
  assign _T_937 = _T_936 & x768_b521_D2; // @[sm_x536_inr_Foreach.scala 145:268:@7618.4]
  assign x532_sum_number = x532_sum_1_io_result; // @[Math.scala 154:22:@7504.4 Math.scala 155:14:@7505.4]
  assign io_in_x472_A_sram_1_wPort_0_ofs_0 = x532_sum_number[8:0]; // @[MemInterfaceType.scala 89:54:@7569.4]
  assign io_in_x472_A_sram_1_wPort_0_data_0 = RetimeWrapper_2_io_out; // @[MemInterfaceType.scala 90:56:@7570.4]
  assign io_in_x472_A_sram_1_wPort_0_en_0 = _T_897 & x765_b504_D2; // @[MemInterfaceType.scala 93:57:@7572.4]
  assign io_in_x471_A_sram_0_wPort_0_ofs_0 = x532_sum_number[8:0]; // @[MemInterfaceType.scala 89:54:@7595.4]
  assign io_in_x471_A_sram_0_wPort_0_data_0 = RetimeWrapper_2_io_out; // @[MemInterfaceType.scala 90:56:@7596.4]
  assign io_in_x471_A_sram_0_wPort_0_en_0 = _T_917 & x765_b504_D2; // @[MemInterfaceType.scala 93:57:@7598.4]
  assign io_in_x476_ready = _T_834 & io_sigsIn_datapathEn; // @[sm_x536_inr_Foreach.scala 110:18:@7468.4]
  assign io_in_x473_A_sram_2_wPort_0_ofs_0 = x532_sum_number[8:0]; // @[MemInterfaceType.scala 89:54:@7621.4]
  assign io_in_x473_A_sram_2_wPort_0_data_0 = RetimeWrapper_2_io_out; // @[MemInterfaceType.scala 90:56:@7622.4]
  assign io_in_x473_A_sram_2_wPort_0_en_0 = _T_937 & x765_b504_D2; // @[MemInterfaceType.scala 93:57:@7624.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@7408.4]
  assign x527_sub_1_clock = clock; // @[:@7457.4]
  assign x527_sub_1_reset = reset; // @[:@7458.4]
  assign x527_sub_1_io_a = __io_result; // @[Math.scala 192:17:@7459.4]
  assign x527_sub_1_io_b = io_in_x505_reg_rPort_0_output_0; // @[Math.scala 193:17:@7460.4]
  assign x527_sub_1_io_flow = 1'h1; // @[Math.scala 194:20:@7461.4]
  assign RetimeWrapper_clock = clock; // @[:@7473.4]
  assign RetimeWrapper_reset = reset; // @[:@7474.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@7476.4]
  assign RetimeWrapper_io_in = io_in_x476_bits_rdata_0; // @[package.scala 94:16:@7475.4]
  assign x743_sum_1_clock = clock; // @[:@7489.4]
  assign x743_sum_1_reset = reset; // @[:@7490.4]
  assign x743_sum_1_io_a = _T_850[31:0]; // @[Math.scala 151:17:@7491.4]
  assign x743_sum_1_io_b = io_in_b503_number; // @[Math.scala 152:17:@7492.4]
  assign x743_sum_1_io_flow = 1'h1; // @[Math.scala 153:20:@7493.4]
  assign x532_sum_1_clock = clock; // @[:@7499.4]
  assign x532_sum_1_reset = reset; // @[:@7500.4]
  assign x532_sum_1_io_a = x743_sum_1_io_result; // @[Math.scala 151:17:@7501.4]
  assign x532_sum_1_io_b = x527_sub_1_io_result; // @[Math.scala 152:17:@7502.4]
  assign x532_sum_1_io_flow = 1'h1; // @[Math.scala 153:20:@7503.4]
  assign RetimeWrapper_1_clock = clock; // @[:@7510.4]
  assign RetimeWrapper_1_reset = reset; // @[:@7511.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@7513.4]
  assign RetimeWrapper_1_io_in = io_in_b504; // @[package.scala 94:16:@7512.4]
  assign RetimeWrapper_2_clock = clock; // @[:@7520.4]
  assign RetimeWrapper_2_reset = reset; // @[:@7521.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@7523.4]
  assign RetimeWrapper_2_io_in = RetimeWrapper_io_out; // @[package.scala 94:16:@7522.4]
  assign RetimeWrapper_3_clock = clock; // @[:@7530.4]
  assign RetimeWrapper_3_reset = reset; // @[:@7531.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@7533.4]
  assign RetimeWrapper_3_io_in = x523 & x525; // @[package.scala 94:16:@7532.4]
  assign RetimeWrapper_4_clock = clock; // @[:@7540.4]
  assign RetimeWrapper_4_reset = reset; // @[:@7541.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@7543.4]
  assign RetimeWrapper_4_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@7542.4]
  assign RetimeWrapper_5_clock = clock; // @[:@7554.4]
  assign RetimeWrapper_5_reset = reset; // @[:@7555.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@7557.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7556.4]
  assign RetimeWrapper_6_clock = clock; // @[:@7580.4]
  assign RetimeWrapper_6_reset = reset; // @[:@7581.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@7583.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7582.4]
  assign RetimeWrapper_7_clock = clock; // @[:@7606.4]
  assign RetimeWrapper_7_reset = reset; // @[:@7607.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@7609.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@7608.4]
endmodule
module x537_outr_Foreach_kernelx537_outr_Foreach_concrete1( // @[:@7626.2]
  input         clock, // @[:@7627.4]
  input         reset, // @[:@7628.4]
  output [8:0]  io_in_x472_A_sram_1_wPort_0_ofs_0, // @[:@7629.4]
  output [31:0] io_in_x472_A_sram_1_wPort_0_data_0, // @[:@7629.4]
  output        io_in_x472_A_sram_1_wPort_0_en_0, // @[:@7629.4]
  output        io_in_x475_fifo_rPort_0_en_0, // @[:@7629.4]
  input  [95:0] io_in_x475_fifo_rPort_0_output_0, // @[:@7629.4]
  input         io_in_x475_fifo_empty, // @[:@7629.4]
  output [8:0]  io_in_x471_A_sram_0_wPort_0_ofs_0, // @[:@7629.4]
  output [31:0] io_in_x471_A_sram_0_wPort_0_data_0, // @[:@7629.4]
  output        io_in_x471_A_sram_0_wPort_0_en_0, // @[:@7629.4]
  output        io_in_x476_ready, // @[:@7629.4]
  input         io_in_x476_valid, // @[:@7629.4]
  input  [31:0] io_in_x476_bits_rdata_0, // @[:@7629.4]
  output [8:0]  io_in_x473_A_sram_2_wPort_0_ofs_0, // @[:@7629.4]
  output [31:0] io_in_x473_A_sram_2_wPort_0_data_0, // @[:@7629.4]
  output        io_in_x473_A_sram_2_wPort_0_en_0, // @[:@7629.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@7629.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@7629.4]
  input         io_sigsIn_smChildAcks_0, // @[:@7629.4]
  input         io_sigsIn_smChildAcks_1, // @[:@7629.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@7629.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@7629.4]
  output        io_sigsOut_smDoneIn_0, // @[:@7629.4]
  output        io_sigsOut_smDoneIn_1, // @[:@7629.4]
  output        io_sigsOut_smMaskIn_0, // @[:@7629.4]
  output        io_sigsOut_smMaskIn_1, // @[:@7629.4]
  input         io_rr // @[:@7629.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@7706.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@7706.4]
  wire  x505_reg_clock; // @[m_x505_reg.scala 27:22:@7715.4]
  wire  x505_reg_reset; // @[m_x505_reg.scala 27:22:@7715.4]
  wire [31:0] x505_reg_io_rPort_0_output_0; // @[m_x505_reg.scala 27:22:@7715.4]
  wire [31:0] x505_reg_io_wPort_0_data_0; // @[m_x505_reg.scala 27:22:@7715.4]
  wire  x505_reg_io_wPort_0_reset; // @[m_x505_reg.scala 27:22:@7715.4]
  wire  x505_reg_io_wPort_0_en_0; // @[m_x505_reg.scala 27:22:@7715.4]
  wire  x506_reg_clock; // @[m_x506_reg.scala 27:22:@7732.4]
  wire  x506_reg_reset; // @[m_x506_reg.scala 27:22:@7732.4]
  wire [31:0] x506_reg_io_rPort_0_output_0; // @[m_x506_reg.scala 27:22:@7732.4]
  wire [31:0] x506_reg_io_wPort_0_data_0; // @[m_x506_reg.scala 27:22:@7732.4]
  wire  x506_reg_io_wPort_0_reset; // @[m_x506_reg.scala 27:22:@7732.4]
  wire  x506_reg_io_wPort_0_en_0; // @[m_x506_reg.scala 27:22:@7732.4]
  wire  x507_reg_clock; // @[m_x507_reg.scala 27:22:@7749.4]
  wire  x507_reg_reset; // @[m_x507_reg.scala 27:22:@7749.4]
  wire [31:0] x507_reg_io_rPort_0_output_0; // @[m_x507_reg.scala 27:22:@7749.4]
  wire [31:0] x507_reg_io_wPort_0_data_0; // @[m_x507_reg.scala 27:22:@7749.4]
  wire  x507_reg_io_wPort_0_reset; // @[m_x507_reg.scala 27:22:@7749.4]
  wire  x507_reg_io_wPort_0_en_0; // @[m_x507_reg.scala 27:22:@7749.4]
  wire  x516_inr_UnitPipe_sm_clock; // @[sm_x516_inr_UnitPipe.scala 34:18:@7802.4]
  wire  x516_inr_UnitPipe_sm_reset; // @[sm_x516_inr_UnitPipe.scala 34:18:@7802.4]
  wire  x516_inr_UnitPipe_sm_io_enable; // @[sm_x516_inr_UnitPipe.scala 34:18:@7802.4]
  wire  x516_inr_UnitPipe_sm_io_done; // @[sm_x516_inr_UnitPipe.scala 34:18:@7802.4]
  wire  x516_inr_UnitPipe_sm_io_doneLatch; // @[sm_x516_inr_UnitPipe.scala 34:18:@7802.4]
  wire  x516_inr_UnitPipe_sm_io_ctrDone; // @[sm_x516_inr_UnitPipe.scala 34:18:@7802.4]
  wire  x516_inr_UnitPipe_sm_io_datapathEn; // @[sm_x516_inr_UnitPipe.scala 34:18:@7802.4]
  wire  x516_inr_UnitPipe_sm_io_ctrInc; // @[sm_x516_inr_UnitPipe.scala 34:18:@7802.4]
  wire  x516_inr_UnitPipe_sm_io_parentAck; // @[sm_x516_inr_UnitPipe.scala 34:18:@7802.4]
  wire  x516_inr_UnitPipe_sm_io_backpressure; // @[sm_x516_inr_UnitPipe.scala 34:18:@7802.4]
  wire  x516_inr_UnitPipe_sm_io_break; // @[sm_x516_inr_UnitPipe.scala 34:18:@7802.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@7864.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@7864.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@7864.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@7864.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@7864.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@7872.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@7872.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@7872.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@7872.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@7872.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x475_fifo_rPort_0_en_0; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire [95:0] x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x475_fifo_rPort_0_output_0; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire [31:0] x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_data_0; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_reset; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_en_0; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_reset; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire [31:0] x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_data_0; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_reset; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_en_0; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_reset; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire [31:0] x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_data_0; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_reset; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_en_0; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_reset; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_forwardpressure; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_break; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_rr; // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
  wire  x519_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@8070.4]
  wire  x519_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@8070.4]
  wire [31:0] x519_ctrchain_io_setup_stops_0; // @[SpatialBlocks.scala 37:22:@8070.4]
  wire  x519_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@8070.4]
  wire  x519_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@8070.4]
  wire [31:0] x519_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@8070.4]
  wire  x519_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@8070.4]
  wire  x519_ctrchain_io_output_noop; // @[SpatialBlocks.scala 37:22:@8070.4]
  wire  x519_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@8070.4]
  wire  x536_inr_Foreach_sm_clock; // @[sm_x536_inr_Foreach.scala 35:18:@8125.4]
  wire  x536_inr_Foreach_sm_reset; // @[sm_x536_inr_Foreach.scala 35:18:@8125.4]
  wire  x536_inr_Foreach_sm_io_enable; // @[sm_x536_inr_Foreach.scala 35:18:@8125.4]
  wire  x536_inr_Foreach_sm_io_done; // @[sm_x536_inr_Foreach.scala 35:18:@8125.4]
  wire  x536_inr_Foreach_sm_io_doneLatch; // @[sm_x536_inr_Foreach.scala 35:18:@8125.4]
  wire  x536_inr_Foreach_sm_io_ctrDone; // @[sm_x536_inr_Foreach.scala 35:18:@8125.4]
  wire  x536_inr_Foreach_sm_io_datapathEn; // @[sm_x536_inr_Foreach.scala 35:18:@8125.4]
  wire  x536_inr_Foreach_sm_io_ctrInc; // @[sm_x536_inr_Foreach.scala 35:18:@8125.4]
  wire  x536_inr_Foreach_sm_io_ctrRst; // @[sm_x536_inr_Foreach.scala 35:18:@8125.4]
  wire  x536_inr_Foreach_sm_io_parentAck; // @[sm_x536_inr_Foreach.scala 35:18:@8125.4]
  wire  x536_inr_Foreach_sm_io_backpressure; // @[sm_x536_inr_Foreach.scala 35:18:@8125.4]
  wire  x536_inr_Foreach_sm_io_break; // @[sm_x536_inr_Foreach.scala 35:18:@8125.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@8154.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@8154.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@8154.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@8154.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@8154.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@8194.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@8194.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@8194.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@8194.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@8194.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@8202.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@8202.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@8202.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@8202.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@8202.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_clock; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_reset; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire [8:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire [31:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_data_0; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_en_0; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_b504; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire [8:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire [31:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_data_0; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_en_0; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x476_ready; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire [31:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x476_bits_rdata_0; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire [31:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_b503_number; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire [31:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x505_reg_rPort_0_output_0; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire [8:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire [31:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_data_0; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_en_0; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire [31:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x506_reg_rPort_0_output_0; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire [31:0] x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_rr; // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
  wire  b504; // @[sm_x537_outr_Foreach.scala 75:18:@7714.4]
  wire  _T_773; // @[package.scala 100:49:@7830.4]
  reg  _T_776; // @[package.scala 48:56:@7831.4]
  reg [31:0] _RAND_0;
  wire  _T_784; // @[sm_x537_outr_Foreach.scala 82:46:@7838.4]
  wire  x516_inr_UnitPipe_mySignalsIn_forwardpressure; // @[sm_x537_outr_Foreach.scala 82:115:@7842.4]
  wire  _T_797; // @[package.scala 96:25:@7869.4 package.scala 96:25:@7870.4]
  wire  _T_803; // @[package.scala 96:25:@7877.4 package.scala 96:25:@7878.4]
  wire  _T_806; // @[SpatialBlocks.scala 137:99:@7880.4]
  wire  x516_inr_UnitPipe_mySignalsIn_baseEn; // @[SpatialBlocks.scala 137:96:@7881.4]
  wire [31:0] x734_rd_x507_number; // @[sm_x537_outr_Foreach.scala 88:30:@8056.4 sm_x537_outr_Foreach.scala 93:202:@8069.4]
  wire  _T_894; // @[package.scala 96:25:@8159.4 package.scala 96:25:@8160.4]
  wire  x536_inr_Foreach_mySignalsIn_forwardpressure; // @[sm_x537_outr_Foreach.scala 101:68:@8166.4]
  wire  _T_903; // @[sm_x537_outr_Foreach.scala 104:32:@8170.4]
  wire  x536_inr_Foreach_mySignalsIn_mask; // @[sm_x537_outr_Foreach.scala 104:74:@8171.4]
  wire  _T_909; // @[package.scala 96:25:@8199.4 package.scala 96:25:@8200.4]
  wire  _T_915; // @[package.scala 96:25:@8207.4 package.scala 96:25:@8208.4]
  wire  _T_918; // @[SpatialBlocks.scala 137:99:@8210.4]
  wire  x536_inr_Foreach_mySignalsIn_baseEn; // @[SpatialBlocks.scala 137:96:@8211.4]
  wire  _T_920; // @[SpatialBlocks.scala 156:36:@8219.4]
  wire  _T_921; // @[SpatialBlocks.scala 156:78:@8220.4]
  wire  _T_928; // @[SpatialBlocks.scala 158:58:@8232.4]
  _ _ ( // @[Math.scala 720:24:@7706.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x505_reg x505_reg ( // @[m_x505_reg.scala 27:22:@7715.4]
    .clock(x505_reg_clock),
    .reset(x505_reg_reset),
    .io_rPort_0_output_0(x505_reg_io_rPort_0_output_0),
    .io_wPort_0_data_0(x505_reg_io_wPort_0_data_0),
    .io_wPort_0_reset(x505_reg_io_wPort_0_reset),
    .io_wPort_0_en_0(x505_reg_io_wPort_0_en_0)
  );
  x505_reg x506_reg ( // @[m_x506_reg.scala 27:22:@7732.4]
    .clock(x506_reg_clock),
    .reset(x506_reg_reset),
    .io_rPort_0_output_0(x506_reg_io_rPort_0_output_0),
    .io_wPort_0_data_0(x506_reg_io_wPort_0_data_0),
    .io_wPort_0_reset(x506_reg_io_wPort_0_reset),
    .io_wPort_0_en_0(x506_reg_io_wPort_0_en_0)
  );
  x505_reg x507_reg ( // @[m_x507_reg.scala 27:22:@7749.4]
    .clock(x507_reg_clock),
    .reset(x507_reg_reset),
    .io_rPort_0_output_0(x507_reg_io_rPort_0_output_0),
    .io_wPort_0_data_0(x507_reg_io_wPort_0_data_0),
    .io_wPort_0_reset(x507_reg_io_wPort_0_reset),
    .io_wPort_0_en_0(x507_reg_io_wPort_0_en_0)
  );
  x516_inr_UnitPipe_sm x516_inr_UnitPipe_sm ( // @[sm_x516_inr_UnitPipe.scala 34:18:@7802.4]
    .clock(x516_inr_UnitPipe_sm_clock),
    .reset(x516_inr_UnitPipe_sm_reset),
    .io_enable(x516_inr_UnitPipe_sm_io_enable),
    .io_done(x516_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x516_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x516_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x516_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x516_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x516_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x516_inr_UnitPipe_sm_io_backpressure),
    .io_break(x516_inr_UnitPipe_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@7864.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@7872.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1 x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1 ( // @[sm_x516_inr_UnitPipe.scala 106:24:@7901.4]
    .io_in_x475_fifo_rPort_0_en_0(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x475_fifo_rPort_0_en_0),
    .io_in_x475_fifo_rPort_0_output_0(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x475_fifo_rPort_0_output_0),
    .io_in_x507_reg_wPort_0_data_0(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_data_0),
    .io_in_x507_reg_wPort_0_reset(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_reset),
    .io_in_x507_reg_wPort_0_en_0(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_en_0),
    .io_in_x507_reg_reset(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_reset),
    .io_in_x505_reg_wPort_0_data_0(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_data_0),
    .io_in_x505_reg_wPort_0_reset(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_reset),
    .io_in_x505_reg_wPort_0_en_0(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_en_0),
    .io_in_x505_reg_reset(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_reset),
    .io_in_x506_reg_wPort_0_data_0(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_data_0),
    .io_in_x506_reg_wPort_0_reset(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_reset),
    .io_in_x506_reg_wPort_0_en_0(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_en_0),
    .io_in_x506_reg_reset(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_reset),
    .io_sigsIn_forwardpressure(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_forwardpressure),
    .io_sigsIn_datapathEn(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_break),
    .io_rr(x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_rr)
  );
  x519_ctrchain x519_ctrchain ( // @[SpatialBlocks.scala 37:22:@8070.4]
    .clock(x519_ctrchain_clock),
    .reset(x519_ctrchain_reset),
    .io_setup_stops_0(x519_ctrchain_io_setup_stops_0),
    .io_input_reset(x519_ctrchain_io_input_reset),
    .io_input_enable(x519_ctrchain_io_input_enable),
    .io_output_counts_0(x519_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x519_ctrchain_io_output_oobs_0),
    .io_output_noop(x519_ctrchain_io_output_noop),
    .io_output_done(x519_ctrchain_io_output_done)
  );
  x536_inr_Foreach_sm x536_inr_Foreach_sm ( // @[sm_x536_inr_Foreach.scala 35:18:@8125.4]
    .clock(x536_inr_Foreach_sm_clock),
    .reset(x536_inr_Foreach_sm_reset),
    .io_enable(x536_inr_Foreach_sm_io_enable),
    .io_done(x536_inr_Foreach_sm_io_done),
    .io_doneLatch(x536_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x536_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x536_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x536_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x536_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x536_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x536_inr_Foreach_sm_io_backpressure),
    .io_break(x536_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@8154.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@8194.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@8202.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x536_inr_Foreach_kernelx536_inr_Foreach_concrete1 x536_inr_Foreach_kernelx536_inr_Foreach_concrete1 ( // @[sm_x536_inr_Foreach.scala 147:24:@8236.4]
    .clock(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_clock),
    .reset(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_reset),
    .io_in_x472_A_sram_1_wPort_0_ofs_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0),
    .io_in_x472_A_sram_1_wPort_0_data_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_data_0),
    .io_in_x472_A_sram_1_wPort_0_en_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_en_0),
    .io_in_b504(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_b504),
    .io_in_x471_A_sram_0_wPort_0_ofs_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0),
    .io_in_x471_A_sram_0_wPort_0_data_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_data_0),
    .io_in_x471_A_sram_0_wPort_0_en_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_en_0),
    .io_in_x476_ready(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x476_ready),
    .io_in_x476_bits_rdata_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x476_bits_rdata_0),
    .io_in_b503_number(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_b503_number),
    .io_in_x505_reg_rPort_0_output_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x505_reg_rPort_0_output_0),
    .io_in_x473_A_sram_2_wPort_0_ofs_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0),
    .io_in_x473_A_sram_2_wPort_0_data_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_data_0),
    .io_in_x473_A_sram_2_wPort_0_en_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_en_0),
    .io_in_x506_reg_rPort_0_output_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x506_reg_rPort_0_output_0),
    .io_sigsIn_datapathEn(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_rr)
  );
  assign b504 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x537_outr_Foreach.scala 75:18:@7714.4]
  assign _T_773 = x516_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@7830.4]
  assign _T_784 = ~ io_in_x475_fifo_empty; // @[sm_x537_outr_Foreach.scala 82:46:@7838.4]
  assign x516_inr_UnitPipe_mySignalsIn_forwardpressure = _T_784 | x516_inr_UnitPipe_sm_io_doneLatch; // @[sm_x537_outr_Foreach.scala 82:115:@7842.4]
  assign _T_797 = RetimeWrapper_io_out; // @[package.scala 96:25:@7869.4 package.scala 96:25:@7870.4]
  assign _T_803 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@7877.4 package.scala 96:25:@7878.4]
  assign _T_806 = ~ _T_803; // @[SpatialBlocks.scala 137:99:@7880.4]
  assign x516_inr_UnitPipe_mySignalsIn_baseEn = _T_797 & _T_806; // @[SpatialBlocks.scala 137:96:@7881.4]
  assign x734_rd_x507_number = x507_reg_io_rPort_0_output_0; // @[sm_x537_outr_Foreach.scala 88:30:@8056.4 sm_x537_outr_Foreach.scala 93:202:@8069.4]
  assign _T_894 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@8159.4 package.scala 96:25:@8160.4]
  assign x536_inr_Foreach_mySignalsIn_forwardpressure = io_in_x476_valid | x536_inr_Foreach_sm_io_doneLatch; // @[sm_x537_outr_Foreach.scala 101:68:@8166.4]
  assign _T_903 = ~ x519_ctrchain_io_output_noop; // @[sm_x537_outr_Foreach.scala 104:32:@8170.4]
  assign x536_inr_Foreach_mySignalsIn_mask = _T_903 & b504; // @[sm_x537_outr_Foreach.scala 104:74:@8171.4]
  assign _T_909 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@8199.4 package.scala 96:25:@8200.4]
  assign _T_915 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@8207.4 package.scala 96:25:@8208.4]
  assign _T_918 = ~ _T_915; // @[SpatialBlocks.scala 137:99:@8210.4]
  assign x536_inr_Foreach_mySignalsIn_baseEn = _T_909 & _T_918; // @[SpatialBlocks.scala 137:96:@8211.4]
  assign _T_920 = x536_inr_Foreach_sm_io_datapathEn & x536_inr_Foreach_mySignalsIn_mask; // @[SpatialBlocks.scala 156:36:@8219.4]
  assign _T_921 = ~ x536_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 156:78:@8220.4]
  assign _T_928 = x536_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 158:58:@8232.4]
  assign io_in_x472_A_sram_1_wPort_0_ofs_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@8342.4]
  assign io_in_x472_A_sram_1_wPort_0_data_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@8341.4]
  assign io_in_x472_A_sram_1_wPort_0_en_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@8337.4]
  assign io_in_x475_fifo_rPort_0_en_0 = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x475_fifo_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@8005.4]
  assign io_in_x471_A_sram_0_wPort_0_ofs_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@8350.4]
  assign io_in_x471_A_sram_0_wPort_0_data_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@8349.4]
  assign io_in_x471_A_sram_0_wPort_0_en_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@8345.4]
  assign io_in_x476_ready = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x476_ready; // @[sm_x536_inr_Foreach.scala 66:23:@8354.4]
  assign io_in_x473_A_sram_2_wPort_0_ofs_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@8366.4]
  assign io_in_x473_A_sram_2_wPort_0_data_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@8365.4]
  assign io_in_x473_A_sram_2_wPort_0_en_0 = x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@8361.4]
  assign io_sigsOut_smDoneIn_0 = x516_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 155:56:@7887.4]
  assign io_sigsOut_smDoneIn_1 = x536_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@8217.4]
  assign io_sigsOut_smMaskIn_0 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[SpatialBlocks.scala 155:86:@7888.4]
  assign io_sigsOut_smMaskIn_1 = _T_903 & b504; // @[SpatialBlocks.scala 155:86:@8218.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@7709.4]
  assign x505_reg_clock = clock; // @[:@7716.4]
  assign x505_reg_reset = reset; // @[:@7717.4]
  assign x505_reg_io_wPort_0_data_0 = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@8019.4]
  assign x505_reg_io_wPort_0_reset = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_reset; // @[MemInterfaceType.scala 67:44:@8018.4]
  assign x505_reg_io_wPort_0_en_0 = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x505_reg_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@8015.4]
  assign x506_reg_clock = clock; // @[:@7733.4]
  assign x506_reg_reset = reset; // @[:@7734.4]
  assign x506_reg_io_wPort_0_data_0 = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@8026.4]
  assign x506_reg_io_wPort_0_reset = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_reset; // @[MemInterfaceType.scala 67:44:@8025.4]
  assign x506_reg_io_wPort_0_en_0 = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x506_reg_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@8022.4]
  assign x507_reg_clock = clock; // @[:@7750.4]
  assign x507_reg_reset = reset; // @[:@7751.4]
  assign x507_reg_io_wPort_0_data_0 = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@8012.4]
  assign x507_reg_io_wPort_0_reset = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_reset; // @[MemInterfaceType.scala 67:44:@8011.4]
  assign x507_reg_io_wPort_0_en_0 = x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x507_reg_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@8008.4]
  assign x516_inr_UnitPipe_sm_clock = clock; // @[:@7803.4]
  assign x516_inr_UnitPipe_sm_reset = reset; // @[:@7804.4]
  assign x516_inr_UnitPipe_sm_io_enable = x516_inr_UnitPipe_mySignalsIn_baseEn & x516_inr_UnitPipe_mySignalsIn_forwardpressure; // @[SpatialBlocks.scala 139:18:@7884.4]
  assign x516_inr_UnitPipe_sm_io_ctrDone = x516_inr_UnitPipe_sm_io_ctrInc & _T_776; // @[sm_x537_outr_Foreach.scala 80:39:@7834.4]
  assign x516_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@7886.4]
  assign x516_inr_UnitPipe_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@7858.4]
  assign x516_inr_UnitPipe_sm_io_break = 1'h0; // @[sm_x537_outr_Foreach.scala 84:37:@7845.4]
  assign RetimeWrapper_clock = clock; // @[:@7865.4]
  assign RetimeWrapper_reset = reset; // @[:@7866.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@7868.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@7867.4]
  assign RetimeWrapper_1_clock = clock; // @[:@7873.4]
  assign RetimeWrapper_1_reset = reset; // @[:@7874.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@7876.4]
  assign RetimeWrapper_1_io_in = x516_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@7875.4]
  assign x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_in_x475_fifo_rPort_0_output_0 = io_in_x475_fifo_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@8003.4]
  assign x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_forwardpressure = _T_784 | x516_inr_UnitPipe_sm_io_doneLatch; // @[sm_x516_inr_UnitPipe.scala 111:22:@8042.4]
  assign x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x516_inr_UnitPipe_sm_io_datapathEn & b504; // @[sm_x516_inr_UnitPipe.scala 111:22:@8041.4]
  assign x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_sigsIn_break = x516_inr_UnitPipe_sm_io_break; // @[sm_x516_inr_UnitPipe.scala 111:22:@8039.4]
  assign x516_inr_UnitPipe_kernelx516_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x516_inr_UnitPipe.scala 110:18:@8029.4]
  assign x519_ctrchain_clock = clock; // @[:@8071.4]
  assign x519_ctrchain_reset = reset; // @[:@8072.4]
  assign x519_ctrchain_io_setup_stops_0 = $signed(x734_rd_x507_number); // @[SpatialBlocks.scala 40:87:@8086.4]
  assign x519_ctrchain_io_input_reset = x536_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@8235.4]
  assign x519_ctrchain_io_input_enable = _T_928 & x536_inr_Foreach_mySignalsIn_forwardpressure; // @[SpatialBlocks.scala 158:42:@8234.4]
  assign x536_inr_Foreach_sm_clock = clock; // @[:@8126.4]
  assign x536_inr_Foreach_sm_reset = reset; // @[:@8127.4]
  assign x536_inr_Foreach_sm_io_enable = x536_inr_Foreach_mySignalsIn_baseEn & x536_inr_Foreach_mySignalsIn_forwardpressure; // @[SpatialBlocks.scala 139:18:@8214.4]
  assign x536_inr_Foreach_sm_io_ctrDone = io_rr ? _T_894 : 1'h0; // @[sm_x537_outr_Foreach.scala 99:38:@8162.4]
  assign x536_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 141:21:@8216.4]
  assign x536_inr_Foreach_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@8188.4]
  assign x536_inr_Foreach_sm_io_break = 1'h0; // @[sm_x537_outr_Foreach.scala 103:36:@8169.4]
  assign RetimeWrapper_2_clock = clock; // @[:@8155.4]
  assign RetimeWrapper_2_reset = reset; // @[:@8156.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@8158.4]
  assign RetimeWrapper_2_io_in = x519_ctrchain_io_output_done; // @[package.scala 94:16:@8157.4]
  assign RetimeWrapper_3_clock = clock; // @[:@8195.4]
  assign RetimeWrapper_3_reset = reset; // @[:@8196.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@8198.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@8197.4]
  assign RetimeWrapper_4_clock = clock; // @[:@8203.4]
  assign RetimeWrapper_4_reset = reset; // @[:@8204.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@8206.4]
  assign RetimeWrapper_4_io_in = x536_inr_Foreach_sm_io_done; // @[package.scala 94:16:@8205.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_clock = clock; // @[:@8237.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_reset = reset; // @[:@8238.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_b504 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x536_inr_Foreach.scala 64:23:@8344.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x476_bits_rdata_0 = io_in_x476_bits_rdata_0; // @[sm_x536_inr_Foreach.scala 66:23:@8352.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_b503_number = __io_result; // @[sm_x536_inr_Foreach.scala 67:23:@8355.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x505_reg_rPort_0_output_0 = x505_reg_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@8356.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_in_x506_reg_rPort_0_output_0 = x506_reg_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@8368.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_920 & _T_921; // @[sm_x536_inr_Foreach.scala 152:22:@8385.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_break = x536_inr_Foreach_sm_io_break; // @[sm_x536_inr_Foreach.scala 152:22:@8383.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x519_ctrchain_io_output_counts_0; // @[sm_x536_inr_Foreach.scala 152:22:@8378.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x519_ctrchain_io_output_oobs_0; // @[sm_x536_inr_Foreach.scala 152:22:@8377.4]
  assign x536_inr_Foreach_kernelx536_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x536_inr_Foreach.scala 151:18:@8373.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_776 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_776 <= 1'h0;
    end else begin
      _T_776 <= _T_773;
    end
  end
endmodule
module x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1( // @[:@8401.2]
  input         clock, // @[:@8402.4]
  input         reset, // @[:@8403.4]
  input  [63:0] io_in_x468_A_dram_number, // @[:@8404.4]
  output [8:0]  io_in_x472_A_sram_1_wPort_0_ofs_0, // @[:@8404.4]
  output [31:0] io_in_x472_A_sram_1_wPort_0_data_0, // @[:@8404.4]
  output        io_in_x472_A_sram_1_wPort_0_en_0, // @[:@8404.4]
  output [8:0]  io_in_x471_A_sram_0_wPort_0_ofs_0, // @[:@8404.4]
  output [31:0] io_in_x471_A_sram_0_wPort_0_data_0, // @[:@8404.4]
  output        io_in_x471_A_sram_0_wPort_0_en_0, // @[:@8404.4]
  output        io_in_x476_ready, // @[:@8404.4]
  input         io_in_x476_valid, // @[:@8404.4]
  input  [31:0] io_in_x476_bits_rdata_0, // @[:@8404.4]
  output [8:0]  io_in_x473_A_sram_2_wPort_0_ofs_0, // @[:@8404.4]
  output [31:0] io_in_x473_A_sram_2_wPort_0_data_0, // @[:@8404.4]
  output        io_in_x473_A_sram_2_wPort_0_en_0, // @[:@8404.4]
  input         io_in_x474_ready, // @[:@8404.4]
  output        io_in_x474_valid, // @[:@8404.4]
  output [63:0] io_in_x474_bits_addr, // @[:@8404.4]
  output [31:0] io_in_x474_bits_size, // @[:@8404.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@8404.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@8404.4]
  input         io_sigsIn_smChildAcks_0, // @[:@8404.4]
  input         io_sigsIn_smChildAcks_1, // @[:@8404.4]
  output        io_sigsOut_smDoneIn_0, // @[:@8404.4]
  output        io_sigsOut_smDoneIn_1, // @[:@8404.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@8404.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@8404.4]
  input         io_rr // @[:@8404.4]
);
  wire  x475_fifo_clock; // @[m_x475_fifo.scala 27:22:@8457.4]
  wire  x475_fifo_reset; // @[m_x475_fifo.scala 27:22:@8457.4]
  wire  x475_fifo_io_rPort_0_en_0; // @[m_x475_fifo.scala 27:22:@8457.4]
  wire [95:0] x475_fifo_io_rPort_0_output_0; // @[m_x475_fifo.scala 27:22:@8457.4]
  wire [95:0] x475_fifo_io_wPort_0_data_0; // @[m_x475_fifo.scala 27:22:@8457.4]
  wire  x475_fifo_io_wPort_0_en_0; // @[m_x475_fifo.scala 27:22:@8457.4]
  wire  x475_fifo_io_full; // @[m_x475_fifo.scala 27:22:@8457.4]
  wire  x475_fifo_io_empty; // @[m_x475_fifo.scala 27:22:@8457.4]
  wire  x475_fifo_io_active_0_in; // @[m_x475_fifo.scala 27:22:@8457.4]
  wire  x475_fifo_io_active_0_out; // @[m_x475_fifo.scala 27:22:@8457.4]
  wire  x478_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@8483.4]
  wire  x478_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@8483.4]
  wire  x478_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@8483.4]
  wire  x478_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@8483.4]
  wire [8:0] x478_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@8483.4]
  wire  x478_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@8483.4]
  wire  x478_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@8483.4]
  wire  x499_inr_Foreach_sm_clock; // @[sm_x499_inr_Foreach.scala 34:18:@8536.4]
  wire  x499_inr_Foreach_sm_reset; // @[sm_x499_inr_Foreach.scala 34:18:@8536.4]
  wire  x499_inr_Foreach_sm_io_enable; // @[sm_x499_inr_Foreach.scala 34:18:@8536.4]
  wire  x499_inr_Foreach_sm_io_done; // @[sm_x499_inr_Foreach.scala 34:18:@8536.4]
  wire  x499_inr_Foreach_sm_io_doneLatch; // @[sm_x499_inr_Foreach.scala 34:18:@8536.4]
  wire  x499_inr_Foreach_sm_io_rst; // @[sm_x499_inr_Foreach.scala 34:18:@8536.4]
  wire  x499_inr_Foreach_sm_io_ctrDone; // @[sm_x499_inr_Foreach.scala 34:18:@8536.4]
  wire  x499_inr_Foreach_sm_io_datapathEn; // @[sm_x499_inr_Foreach.scala 34:18:@8536.4]
  wire  x499_inr_Foreach_sm_io_ctrInc; // @[sm_x499_inr_Foreach.scala 34:18:@8536.4]
  wire  x499_inr_Foreach_sm_io_ctrRst; // @[sm_x499_inr_Foreach.scala 34:18:@8536.4]
  wire  x499_inr_Foreach_sm_io_parentAck; // @[sm_x499_inr_Foreach.scala 34:18:@8536.4]
  wire  x499_inr_Foreach_sm_io_backpressure; // @[sm_x499_inr_Foreach.scala 34:18:@8536.4]
  wire  x499_inr_Foreach_sm_io_break; // @[sm_x499_inr_Foreach.scala 34:18:@8536.4]
  wire  x499_inr_Foreach_iiCtr_clock; // @[sm_x499_inr_Foreach.scala 35:21:@8561.4]
  wire  x499_inr_Foreach_iiCtr_reset; // @[sm_x499_inr_Foreach.scala 35:21:@8561.4]
  wire  x499_inr_Foreach_iiCtr_io_input_enable; // @[sm_x499_inr_Foreach.scala 35:21:@8561.4]
  wire  x499_inr_Foreach_iiCtr_io_input_reset; // @[sm_x499_inr_Foreach.scala 35:21:@8561.4]
  wire  x499_inr_Foreach_iiCtr_io_output_issue; // @[sm_x499_inr_Foreach.scala 35:21:@8561.4]
  wire  x499_inr_Foreach_iiCtr_io_output_done; // @[sm_x499_inr_Foreach.scala 35:21:@8561.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@8565.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@8565.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@8565.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@8565.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@8565.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@8574.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@8574.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@8574.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@8574.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@8574.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@8617.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@8617.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@8617.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@8617.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@8617.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@8625.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@8625.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@8625.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@8625.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@8625.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_clock; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_reset; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire [63:0] x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x468_A_dram_number; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire [95:0] x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_wPort_0_data_0; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_wPort_0_en_0; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_full; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_active_0_in; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_active_0_out; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_ready; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_valid; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire [63:0] x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_bits_addr; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire [31:0] x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_bits_size; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_iiIssue; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire [31:0] x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_rr; // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
  wire  x502_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@8765.4]
  wire  x502_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@8765.4]
  wire  x502_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@8765.4]
  wire  x502_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@8765.4]
  wire [8:0] x502_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@8765.4]
  wire  x502_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@8765.4]
  wire  x502_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@8765.4]
  wire  x537_outr_Foreach_sm_clock; // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
  wire  x537_outr_Foreach_sm_reset; // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
  wire  x537_outr_Foreach_sm_io_enable; // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
  wire  x537_outr_Foreach_sm_io_done; // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
  wire  x537_outr_Foreach_sm_io_ctrDone; // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
  wire  x537_outr_Foreach_sm_io_ctrInc; // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
  wire  x537_outr_Foreach_sm_io_ctrRst; // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
  wire  x537_outr_Foreach_sm_io_parentAck; // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
  wire  x537_outr_Foreach_sm_io_doneIn_0; // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
  wire  x537_outr_Foreach_sm_io_doneIn_1; // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
  wire  x537_outr_Foreach_sm_io_maskIn_0; // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
  wire  x537_outr_Foreach_sm_io_maskIn_1; // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
  wire  x537_outr_Foreach_sm_io_enableOut_0; // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
  wire  x537_outr_Foreach_sm_io_enableOut_1; // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
  wire  x537_outr_Foreach_sm_io_childAck_0; // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
  wire  x537_outr_Foreach_sm_io_childAck_1; // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@8857.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@8857.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@8857.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@8857.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@8857.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@8902.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@8902.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@8902.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@8902.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@8902.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@8910.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@8910.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@8910.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@8910.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@8910.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_clock; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_reset; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire [8:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire [31:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_data_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_en_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_rPort_0_en_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire [95:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_rPort_0_output_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_empty; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire [8:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire [31:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_data_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_en_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_ready; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_valid; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire [31:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_bits_rdata_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire [8:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire [31:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_data_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_en_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire [31:0] x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_rr; // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
  wire  _T_602; // @[package.scala 96:25:@8570.4 package.scala 96:25:@8571.4]
  wire  _T_608; // @[package.scala 96:25:@8579.4 package.scala 96:25:@8580.4]
  wire  _T_611; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 86:41:@8582.4]
  wire  _T_612; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 86:68:@8583.4]
  wire  _T_613; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 86:66:@8584.4]
  wire  _T_614; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 86:96:@8585.4]
  wire  _T_628; // @[package.scala 96:25:@8622.4 package.scala 96:25:@8623.4]
  wire  _T_634; // @[package.scala 96:25:@8630.4 package.scala 96:25:@8631.4]
  wire  _T_637; // @[SpatialBlocks.scala 137:99:@8633.4]
  wire  _T_639; // @[SpatialBlocks.scala 156:36:@8642.4]
  wire  _T_640; // @[SpatialBlocks.scala 156:78:@8643.4]
  wire  x499_inr_Foreach_mySignalsIn_iiDone; // @[SpatialBlocks.scala 157:126:@8650.4]
  wire  _T_711; // @[package.scala 96:25:@8862.4 package.scala 96:25:@8863.4]
  wire  _T_728; // @[package.scala 96:25:@8907.4 package.scala 96:25:@8908.4]
  wire  _T_734; // @[package.scala 96:25:@8915.4 package.scala 96:25:@8916.4]
  wire  _T_737; // @[SpatialBlocks.scala 137:99:@8918.4]
  x475_fifo x475_fifo ( // @[m_x475_fifo.scala 27:22:@8457.4]
    .clock(x475_fifo_clock),
    .reset(x475_fifo_reset),
    .io_rPort_0_en_0(x475_fifo_io_rPort_0_en_0),
    .io_rPort_0_output_0(x475_fifo_io_rPort_0_output_0),
    .io_wPort_0_data_0(x475_fifo_io_wPort_0_data_0),
    .io_wPort_0_en_0(x475_fifo_io_wPort_0_en_0),
    .io_full(x475_fifo_io_full),
    .io_empty(x475_fifo_io_empty),
    .io_active_0_in(x475_fifo_io_active_0_in),
    .io_active_0_out(x475_fifo_io_active_0_out)
  );
  x478_ctrchain x478_ctrchain ( // @[SpatialBlocks.scala 37:22:@8483.4]
    .clock(x478_ctrchain_clock),
    .reset(x478_ctrchain_reset),
    .io_input_reset(x478_ctrchain_io_input_reset),
    .io_input_enable(x478_ctrchain_io_input_enable),
    .io_output_counts_0(x478_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x478_ctrchain_io_output_oobs_0),
    .io_output_done(x478_ctrchain_io_output_done)
  );
  x499_inr_Foreach_sm x499_inr_Foreach_sm ( // @[sm_x499_inr_Foreach.scala 34:18:@8536.4]
    .clock(x499_inr_Foreach_sm_clock),
    .reset(x499_inr_Foreach_sm_reset),
    .io_enable(x499_inr_Foreach_sm_io_enable),
    .io_done(x499_inr_Foreach_sm_io_done),
    .io_doneLatch(x499_inr_Foreach_sm_io_doneLatch),
    .io_rst(x499_inr_Foreach_sm_io_rst),
    .io_ctrDone(x499_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x499_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x499_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x499_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x499_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x499_inr_Foreach_sm_io_backpressure),
    .io_break(x499_inr_Foreach_sm_io_break)
  );
  x499_inr_Foreach_iiCtr x499_inr_Foreach_iiCtr ( // @[sm_x499_inr_Foreach.scala 35:21:@8561.4]
    .clock(x499_inr_Foreach_iiCtr_clock),
    .reset(x499_inr_Foreach_iiCtr_reset),
    .io_input_enable(x499_inr_Foreach_iiCtr_io_input_enable),
    .io_input_reset(x499_inr_Foreach_iiCtr_io_input_reset),
    .io_output_issue(x499_inr_Foreach_iiCtr_io_output_issue),
    .io_output_done(x499_inr_Foreach_iiCtr_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@8565.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@8574.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@8617.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@8625.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x499_inr_Foreach_kernelx499_inr_Foreach_concrete1 x499_inr_Foreach_kernelx499_inr_Foreach_concrete1 ( // @[sm_x499_inr_Foreach.scala 124:24:@8660.4]
    .clock(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_clock),
    .reset(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_reset),
    .io_in_x468_A_dram_number(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x468_A_dram_number),
    .io_in_x475_fifo_wPort_0_data_0(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_wPort_0_data_0),
    .io_in_x475_fifo_wPort_0_en_0(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_wPort_0_en_0),
    .io_in_x475_fifo_full(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_full),
    .io_in_x475_fifo_active_0_in(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_active_0_in),
    .io_in_x475_fifo_active_0_out(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_active_0_out),
    .io_in_x474_ready(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_ready),
    .io_in_x474_valid(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_valid),
    .io_in_x474_bits_addr(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_bits_addr),
    .io_in_x474_bits_size(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_bits_size),
    .io_sigsIn_iiIssue(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_iiIssue),
    .io_sigsIn_backpressure(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_rr)
  );
  x478_ctrchain x502_ctrchain ( // @[SpatialBlocks.scala 37:22:@8765.4]
    .clock(x502_ctrchain_clock),
    .reset(x502_ctrchain_reset),
    .io_input_reset(x502_ctrchain_io_input_reset),
    .io_input_enable(x502_ctrchain_io_input_enable),
    .io_output_counts_0(x502_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x502_ctrchain_io_output_oobs_0),
    .io_output_done(x502_ctrchain_io_output_done)
  );
  x537_outr_Foreach_sm x537_outr_Foreach_sm ( // @[sm_x537_outr_Foreach.scala 34:18:@8823.4]
    .clock(x537_outr_Foreach_sm_clock),
    .reset(x537_outr_Foreach_sm_reset),
    .io_enable(x537_outr_Foreach_sm_io_enable),
    .io_done(x537_outr_Foreach_sm_io_done),
    .io_ctrDone(x537_outr_Foreach_sm_io_ctrDone),
    .io_ctrInc(x537_outr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x537_outr_Foreach_sm_io_ctrRst),
    .io_parentAck(x537_outr_Foreach_sm_io_parentAck),
    .io_doneIn_0(x537_outr_Foreach_sm_io_doneIn_0),
    .io_doneIn_1(x537_outr_Foreach_sm_io_doneIn_1),
    .io_maskIn_0(x537_outr_Foreach_sm_io_maskIn_0),
    .io_maskIn_1(x537_outr_Foreach_sm_io_maskIn_1),
    .io_enableOut_0(x537_outr_Foreach_sm_io_enableOut_0),
    .io_enableOut_1(x537_outr_Foreach_sm_io_enableOut_1),
    .io_childAck_0(x537_outr_Foreach_sm_io_childAck_0),
    .io_childAck_1(x537_outr_Foreach_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@8857.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@8902.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@8910.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x537_outr_Foreach_kernelx537_outr_Foreach_concrete1 x537_outr_Foreach_kernelx537_outr_Foreach_concrete1 ( // @[sm_x537_outr_Foreach.scala 108:24:@8945.4]
    .clock(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_clock),
    .reset(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_reset),
    .io_in_x472_A_sram_1_wPort_0_ofs_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0),
    .io_in_x472_A_sram_1_wPort_0_data_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_data_0),
    .io_in_x472_A_sram_1_wPort_0_en_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_en_0),
    .io_in_x475_fifo_rPort_0_en_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_rPort_0_en_0),
    .io_in_x475_fifo_rPort_0_output_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_rPort_0_output_0),
    .io_in_x475_fifo_empty(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_empty),
    .io_in_x471_A_sram_0_wPort_0_ofs_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0),
    .io_in_x471_A_sram_0_wPort_0_data_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_data_0),
    .io_in_x471_A_sram_0_wPort_0_en_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_en_0),
    .io_in_x476_ready(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_ready),
    .io_in_x476_valid(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_valid),
    .io_in_x476_bits_rdata_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_bits_rdata_0),
    .io_in_x473_A_sram_2_wPort_0_ofs_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0),
    .io_in_x473_A_sram_2_wPort_0_data_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_data_0),
    .io_in_x473_A_sram_2_wPort_0_en_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_en_0),
    .io_sigsIn_smEnableOuts_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsOut_smDoneIn_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smMaskIn_0(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0),
    .io_sigsOut_smMaskIn_1(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1),
    .io_rr(x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_rr)
  );
  assign _T_602 = RetimeWrapper_io_out; // @[package.scala 96:25:@8570.4 package.scala 96:25:@8571.4]
  assign _T_608 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@8579.4 package.scala 96:25:@8580.4]
  assign _T_611 = ~ _T_608; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 86:41:@8582.4]
  assign _T_612 = ~ x475_fifo_io_active_0_out; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 86:68:@8583.4]
  assign _T_613 = _T_611 | _T_612; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 86:66:@8584.4]
  assign _T_614 = _T_613 & io_in_x474_ready; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 86:96:@8585.4]
  assign _T_628 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@8622.4 package.scala 96:25:@8623.4]
  assign _T_634 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@8630.4 package.scala 96:25:@8631.4]
  assign _T_637 = ~ _T_634; // @[SpatialBlocks.scala 137:99:@8633.4]
  assign _T_639 = x499_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 156:36:@8642.4]
  assign _T_640 = ~ x499_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 156:78:@8643.4]
  assign x499_inr_Foreach_mySignalsIn_iiDone = x499_inr_Foreach_iiCtr_io_output_done; // @[SpatialBlocks.scala 157:126:@8650.4]
  assign _T_711 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@8862.4 package.scala 96:25:@8863.4]
  assign _T_728 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@8907.4 package.scala 96:25:@8908.4]
  assign _T_734 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@8915.4 package.scala 96:25:@8916.4]
  assign _T_737 = ~ _T_734; // @[SpatialBlocks.scala 137:99:@8918.4]
  assign io_in_x472_A_sram_1_wPort_0_ofs_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@9050.4]
  assign io_in_x472_A_sram_1_wPort_0_data_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@9049.4]
  assign io_in_x472_A_sram_1_wPort_0_en_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x472_A_sram_1_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@9045.4]
  assign io_in_x471_A_sram_0_wPort_0_ofs_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@9070.4]
  assign io_in_x471_A_sram_0_wPort_0_data_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@9069.4]
  assign io_in_x471_A_sram_0_wPort_0_en_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x471_A_sram_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@9065.4]
  assign io_in_x476_ready = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_ready; // @[sm_x537_outr_Foreach.scala 59:23:@9074.4]
  assign io_in_x473_A_sram_2_wPort_0_ofs_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@9080.4]
  assign io_in_x473_A_sram_2_wPort_0_data_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@9079.4]
  assign io_in_x473_A_sram_2_wPort_0_en_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x473_A_sram_2_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@9075.4]
  assign io_in_x474_valid = x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_valid; // @[sm_x499_inr_Foreach.scala 54:23:@8736.4]
  assign io_in_x474_bits_addr = x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_bits_addr; // @[sm_x499_inr_Foreach.scala 54:23:@8735.4]
  assign io_in_x474_bits_size = x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_bits_size; // @[sm_x499_inr_Foreach.scala 54:23:@8734.4]
  assign io_sigsOut_smDoneIn_0 = x499_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@8640.4]
  assign io_sigsOut_smDoneIn_1 = x537_outr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@8925.4]
  assign io_sigsOut_smCtrCopyDone_0 = x499_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 170:140:@8659.4]
  assign io_sigsOut_smCtrCopyDone_1 = x537_outr_Foreach_sm_io_done; // @[SpatialBlocks.scala 170:140:@8944.4]
  assign x475_fifo_clock = clock; // @[:@8458.4]
  assign x475_fifo_reset = reset; // @[:@8459.4]
  assign x475_fifo_io_rPort_0_en_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@9062.4]
  assign x475_fifo_io_wPort_0_data_0 = x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@8731.4]
  assign x475_fifo_io_wPort_0_en_0 = x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@8727.4]
  assign x475_fifo_io_active_0_in = x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_active_0_in; // @[MemInterfaceType.scala 167:86:@8726.4]
  assign x478_ctrchain_clock = clock; // @[:@8484.4]
  assign x478_ctrchain_reset = reset; // @[:@8485.4]
  assign x478_ctrchain_io_input_reset = x499_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@8658.4]
  assign x478_ctrchain_io_input_enable = x499_inr_Foreach_sm_io_ctrInc & x499_inr_Foreach_mySignalsIn_iiDone; // @[SpatialBlocks.scala 158:42:@8657.4]
  assign x499_inr_Foreach_sm_clock = clock; // @[:@8537.4]
  assign x499_inr_Foreach_sm_reset = reset; // @[:@8538.4]
  assign x499_inr_Foreach_sm_io_enable = _T_628 & _T_637; // @[SpatialBlocks.scala 139:18:@8637.4]
  assign x499_inr_Foreach_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 133:15:@8612.4]
  assign x499_inr_Foreach_sm_io_ctrDone = io_rr ? _T_602 : 1'h0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 85:38:@8573.4]
  assign x499_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@8639.4]
  assign x499_inr_Foreach_sm_io_backpressure = _T_614 | x499_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 132:24:@8611.4]
  assign x499_inr_Foreach_sm_io_break = 1'h0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 89:36:@8592.4]
  assign x499_inr_Foreach_iiCtr_clock = clock; // @[:@8562.4]
  assign x499_inr_Foreach_iiCtr_reset = reset; // @[:@8563.4]
  assign x499_inr_Foreach_iiCtr_io_input_enable = _T_639 & _T_640; // @[SpatialBlocks.scala 157:27:@8646.4]
  assign x499_inr_Foreach_iiCtr_io_input_reset = x499_inr_Foreach_sm_io_rst | x499_inr_Foreach_sm_io_parentAck; // @[SpatialBlocks.scala 157:63:@8648.4]
  assign RetimeWrapper_clock = clock; // @[:@8566.4]
  assign RetimeWrapper_reset = reset; // @[:@8567.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@8569.4]
  assign RetimeWrapper_io_in = x478_ctrchain_io_output_done; // @[package.scala 94:16:@8568.4]
  assign RetimeWrapper_1_clock = clock; // @[:@8575.4]
  assign RetimeWrapper_1_reset = reset; // @[:@8576.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@8578.4]
  assign RetimeWrapper_1_io_in = x475_fifo_io_full; // @[package.scala 94:16:@8577.4]
  assign RetimeWrapper_2_clock = clock; // @[:@8618.4]
  assign RetimeWrapper_2_reset = reset; // @[:@8619.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@8621.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@8620.4]
  assign RetimeWrapper_3_clock = clock; // @[:@8626.4]
  assign RetimeWrapper_3_reset = reset; // @[:@8627.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@8629.4]
  assign RetimeWrapper_3_io_in = x499_inr_Foreach_sm_io_done; // @[package.scala 94:16:@8628.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_clock = clock; // @[:@8661.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_reset = reset; // @[:@8662.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x468_A_dram_number = io_in_x468_A_dram_number; // @[sm_x499_inr_Foreach.scala 52:30:@8718.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_full = x475_fifo_io_full; // @[MemInterfaceType.scala 159:15:@8721.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x475_fifo_active_0_out = x475_fifo_io_active_0_out; // @[MemInterfaceType.scala 158:75:@8719.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_in_x474_ready = io_in_x474_ready; // @[sm_x499_inr_Foreach.scala 54:23:@8737.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_iiIssue = x499_inr_Foreach_iiCtr_io_output_issue; // @[sm_x499_inr_Foreach.scala 129:22:@8754.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_614 | x499_inr_Foreach_sm_io_doneLatch; // @[sm_x499_inr_Foreach.scala 129:22:@8752.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_639 & _T_640; // @[sm_x499_inr_Foreach.scala 129:22:@8750.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_break = x499_inr_Foreach_sm_io_break; // @[sm_x499_inr_Foreach.scala 129:22:@8748.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{23{x478_ctrchain_io_output_counts_0[8]}},x478_ctrchain_io_output_counts_0}; // @[sm_x499_inr_Foreach.scala 129:22:@8743.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x478_ctrchain_io_output_oobs_0; // @[sm_x499_inr_Foreach.scala 129:22:@8742.4]
  assign x499_inr_Foreach_kernelx499_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x499_inr_Foreach.scala 128:18:@8738.4]
  assign x502_ctrchain_clock = clock; // @[:@8766.4]
  assign x502_ctrchain_reset = reset; // @[:@8767.4]
  assign x502_ctrchain_io_input_reset = x537_outr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@8943.4]
  assign x502_ctrchain_io_input_enable = x537_outr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 158:42:@8942.4]
  assign x537_outr_Foreach_sm_clock = clock; // @[:@8824.4]
  assign x537_outr_Foreach_sm_reset = reset; // @[:@8825.4]
  assign x537_outr_Foreach_sm_io_enable = _T_728 & _T_737; // @[SpatialBlocks.scala 139:18:@8922.4]
  assign x537_outr_Foreach_sm_io_ctrDone = io_rr ? _T_711 : 1'h0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 98:39:@8865.4]
  assign x537_outr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 141:21:@8924.4]
  assign x537_outr_Foreach_sm_io_doneIn_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@8892.4]
  assign x537_outr_Foreach_sm_io_doneIn_1 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:72:@8893.4]
  assign x537_outr_Foreach_sm_io_maskIn_0 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0; // @[SpatialBlocks.scala 131:72:@8894.4]
  assign x537_outr_Foreach_sm_io_maskIn_1 = x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1; // @[SpatialBlocks.scala 131:72:@8895.4]
  assign RetimeWrapper_4_clock = clock; // @[:@8858.4]
  assign RetimeWrapper_4_reset = reset; // @[:@8859.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@8861.4]
  assign RetimeWrapper_4_io_in = x502_ctrchain_io_output_done; // @[package.scala 94:16:@8860.4]
  assign RetimeWrapper_5_clock = clock; // @[:@8903.4]
  assign RetimeWrapper_5_reset = reset; // @[:@8904.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@8906.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@8905.4]
  assign RetimeWrapper_6_clock = clock; // @[:@8911.4]
  assign RetimeWrapper_6_reset = reset; // @[:@8912.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@8914.4]
  assign RetimeWrapper_6_io_in = x537_outr_Foreach_sm_io_done; // @[package.scala 94:16:@8913.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_clock = clock; // @[:@8946.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_reset = reset; // @[:@8947.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_rPort_0_output_0 = x475_fifo_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@9060.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x475_fifo_empty = x475_fifo_io_empty; // @[MemInterfaceType.scala 161:16:@9056.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_valid = io_in_x476_valid; // @[sm_x537_outr_Foreach.scala 59:23:@9073.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_in_x476_bits_rdata_0 = io_in_x476_bits_rdata_0; // @[sm_x537_outr_Foreach.scala 59:23:@9072.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0 = x537_outr_Foreach_sm_io_enableOut_0; // @[sm_x537_outr_Foreach.scala 113:22:@9092.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1 = x537_outr_Foreach_sm_io_enableOut_1; // @[sm_x537_outr_Foreach.scala 113:22:@9093.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0 = x537_outr_Foreach_sm_io_childAck_0; // @[sm_x537_outr_Foreach.scala 113:22:@9088.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1 = x537_outr_Foreach_sm_io_childAck_1; // @[sm_x537_outr_Foreach.scala 113:22:@9089.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{23{x502_ctrchain_io_output_counts_0[8]}},x502_ctrchain_io_output_counts_0}; // @[sm_x537_outr_Foreach.scala 113:22:@9087.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x502_ctrchain_io_output_oobs_0; // @[sm_x537_outr_Foreach.scala 113:22:@9086.4]
  assign x537_outr_Foreach_kernelx537_outr_Foreach_concrete1_io_rr = io_rr; // @[sm_x537_outr_Foreach.scala 112:18:@9082.4]
endmodule
module x668_outr_Foreach_sm( // @[:@9761.2]
  input   clock, // @[:@9762.4]
  input   reset, // @[:@9763.4]
  input   io_enable, // @[:@9764.4]
  output  io_done, // @[:@9764.4]
  input   io_ctrDone, // @[:@9764.4]
  output  io_ctrInc, // @[:@9764.4]
  output  io_ctrRst, // @[:@9764.4]
  input   io_parentAck, // @[:@9764.4]
  input   io_doneIn_0, // @[:@9764.4]
  input   io_doneIn_1, // @[:@9764.4]
  input   io_maskIn_0, // @[:@9764.4]
  input   io_maskIn_1, // @[:@9764.4]
  output  io_enableOut_0, // @[:@9764.4]
  output  io_enableOut_1, // @[:@9764.4]
  output  io_childAck_0, // @[:@9764.4]
  output  io_childAck_1 // @[:@9764.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@9767.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@9767.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@9767.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@9767.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@9767.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@9767.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@9770.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@9770.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@9770.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@9770.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@9770.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@9770.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@9773.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@9773.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@9773.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@9773.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@9773.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@9773.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@9776.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@9776.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@9776.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@9776.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@9776.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@9776.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@9805.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@9805.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@9805.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@9805.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@9805.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@9805.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@9808.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@9808.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@9808.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@9808.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@9808.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@9808.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@9836.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@9836.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@9836.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@9836.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@9836.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@9849.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@9849.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@9849.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@9849.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@9849.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@9875.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@9875.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@9875.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@9875.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@9875.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@9895.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@9895.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@9895.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@9895.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@9895.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@9944.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@9944.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@9944.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@9944.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@9944.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@9961.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@9961.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@9961.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@9961.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@9961.4]
  wire  allDone; // @[Controllers.scala 80:47:@9779.4]
  wire  _T_128; // @[Controllers.scala 102:95:@9835.4]
  wire  _T_127; // @[Controllers.scala 101:55:@9834.4]
  wire  _T_132; // @[package.scala 96:25:@9841.4 package.scala 96:25:@9842.4]
  wire  _T_135; // @[Controllers.scala 102:142:@9844.4]
  wire  _T_136; // @[Controllers.scala 102:138:@9845.4]
  wire  _T_137; // @[Controllers.scala 102:123:@9846.4]
  wire  _T_138; // @[Controllers.scala 102:112:@9847.4]
  wire  _T_139; // @[Controllers.scala 102:95:@9848.4]
  wire  _T_143; // @[package.scala 96:25:@9854.4 package.scala 96:25:@9855.4]
  wire  _T_146; // @[Controllers.scala 102:142:@9857.4]
  wire  _T_147; // @[Controllers.scala 102:138:@9858.4]
  wire  _T_148; // @[Controllers.scala 102:123:@9859.4]
  wire  _T_149; // @[Controllers.scala 102:112:@9860.4]
  wire  synchronize; // @[Controllers.scala 102:164:@9861.4]
  wire  _T_152; // @[Controllers.scala 105:33:@9863.4]
  wire  _T_154; // @[Controllers.scala 105:54:@9864.4]
  wire  _T_155; // @[Controllers.scala 105:52:@9865.4]
  wire  _T_161; // @[Controllers.scala 107:51:@9872.4]
  wire  _T_164; // @[Controllers.scala 107:64:@9874.4]
  wire  _T_168; // @[package.scala 96:25:@9880.4 package.scala 96:25:@9881.4]
  wire  _T_172; // @[Controllers.scala 107:89:@9883.4]
  wire  _T_173; // @[Controllers.scala 107:86:@9884.4]
  wire  _T_174; // @[Controllers.scala 107:108:@9885.4]
  wire  _T_189; // @[Controllers.scala 114:49:@9903.4]
  wire  _T_192; // @[Controllers.scala 115:57:@9907.4]
  wire  _T_203; // @[Controllers.scala 213:68:@9922.4]
  wire  _T_204; // @[Controllers.scala 213:92:@9923.4]
  wire  _T_205; // @[Controllers.scala 213:90:@9924.4]
  wire  _T_206; // @[Controllers.scala 213:115:@9925.4]
  wire  _T_207; // @[Controllers.scala 213:132:@9926.4]
  wire  _T_208; // @[Controllers.scala 213:130:@9927.4]
  wire  _T_209; // @[Controllers.scala 213:156:@9928.4]
  wire  _T_211; // @[Controllers.scala 213:68:@9931.4]
  wire  _T_212; // @[Controllers.scala 213:92:@9932.4]
  wire  _T_213; // @[Controllers.scala 213:90:@9933.4]
  wire  _T_214; // @[Controllers.scala 213:115:@9934.4]
  wire  _T_220; // @[package.scala 100:49:@9939.4]
  reg  _T_223; // @[package.scala 48:56:@9940.4]
  reg [31:0] _RAND_0;
  wire  _T_224; // @[package.scala 100:41:@9942.4]
  reg  _T_237; // @[package.scala 48:56:@9958.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@9767.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@9770.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@9773.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@9776.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@9805.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@9808.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@9836.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@9849.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@9875.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@9895.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@9944.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@9961.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@9779.4]
  assign _T_128 = active_0_io_output == iterDone_0_io_output; // @[Controllers.scala 102:95:@9835.4]
  assign _T_127 = iterDone_0_io_output | iterDone_1_io_output; // @[Controllers.scala 101:55:@9834.4]
  assign _T_132 = RetimeWrapper_io_out; // @[package.scala 96:25:@9841.4 package.scala 96:25:@9842.4]
  assign _T_135 = ~ _T_132; // @[Controllers.scala 102:142:@9844.4]
  assign _T_136 = active_0_io_output == _T_135; // @[Controllers.scala 102:138:@9845.4]
  assign _T_137 = _T_127 & _T_136; // @[Controllers.scala 102:123:@9846.4]
  assign _T_138 = _T_128 | _T_137; // @[Controllers.scala 102:112:@9847.4]
  assign _T_139 = active_1_io_output == iterDone_1_io_output; // @[Controllers.scala 102:95:@9848.4]
  assign _T_143 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@9854.4 package.scala 96:25:@9855.4]
  assign _T_146 = ~ _T_143; // @[Controllers.scala 102:142:@9857.4]
  assign _T_147 = active_1_io_output == _T_146; // @[Controllers.scala 102:138:@9858.4]
  assign _T_148 = _T_127 & _T_147; // @[Controllers.scala 102:123:@9859.4]
  assign _T_149 = _T_139 | _T_148; // @[Controllers.scala 102:112:@9860.4]
  assign synchronize = _T_138 & _T_149; // @[Controllers.scala 102:164:@9861.4]
  assign _T_152 = done_0_io_output == 1'h0; // @[Controllers.scala 105:33:@9863.4]
  assign _T_154 = io_ctrDone == 1'h0; // @[Controllers.scala 105:54:@9864.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 105:52:@9865.4]
  assign _T_161 = synchronize == 1'h0; // @[Controllers.scala 107:51:@9872.4]
  assign _T_164 = _T_161 & _T_152; // @[Controllers.scala 107:64:@9874.4]
  assign _T_168 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@9880.4 package.scala 96:25:@9881.4]
  assign _T_172 = _T_168 == 1'h0; // @[Controllers.scala 107:89:@9883.4]
  assign _T_173 = _T_164 & _T_172; // @[Controllers.scala 107:86:@9884.4]
  assign _T_174 = _T_173 & io_enable; // @[Controllers.scala 107:108:@9885.4]
  assign _T_189 = synchronize & active_0_io_output; // @[Controllers.scala 114:49:@9903.4]
  assign _T_192 = done_0_io_output & synchronize; // @[Controllers.scala 115:57:@9907.4]
  assign _T_203 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@9922.4]
  assign _T_204 = ~ iterDone_0_io_output; // @[Controllers.scala 213:92:@9923.4]
  assign _T_205 = _T_203 & _T_204; // @[Controllers.scala 213:90:@9924.4]
  assign _T_206 = _T_205 & io_maskIn_0; // @[Controllers.scala 213:115:@9925.4]
  assign _T_207 = ~ allDone; // @[Controllers.scala 213:132:@9926.4]
  assign _T_208 = _T_206 & _T_207; // @[Controllers.scala 213:130:@9927.4]
  assign _T_209 = ~ io_ctrDone; // @[Controllers.scala 213:156:@9928.4]
  assign _T_211 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@9931.4]
  assign _T_212 = ~ iterDone_1_io_output; // @[Controllers.scala 213:92:@9932.4]
  assign _T_213 = _T_211 & _T_212; // @[Controllers.scala 213:90:@9933.4]
  assign _T_214 = _T_213 & io_maskIn_1; // @[Controllers.scala 213:115:@9934.4]
  assign _T_220 = allDone == 1'h0; // @[package.scala 100:49:@9939.4]
  assign _T_224 = allDone & _T_223; // @[package.scala 100:41:@9942.4]
  assign io_done = RetimeWrapper_5_io_out; // @[Controllers.scala 245:13:@9968.4]
  assign io_ctrInc = iterDone_0_io_output & synchronize; // @[Controllers.scala 98:17:@9833.4]
  assign io_ctrRst = RetimeWrapper_4_io_out; // @[Controllers.scala 215:13:@9951.4]
  assign io_enableOut_0 = _T_208 & _T_209; // @[Controllers.scala 213:55:@9930.4]
  assign io_enableOut_1 = _T_214 & _T_207; // @[Controllers.scala 213:55:@9938.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@9919.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@9921.4]
  assign active_0_clock = clock; // @[:@9768.4]
  assign active_0_reset = reset; // @[:@9769.4]
  assign active_0_io_input_set = _T_155 & io_enable; // @[Controllers.scala 105:30:@9868.4]
  assign active_0_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 106:32:@9871.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@9782.4]
  assign active_1_clock = clock; // @[:@9771.4]
  assign active_1_reset = reset; // @[:@9772.4]
  assign active_1_io_input_set = _T_189 & io_enable; // @[Controllers.scala 114:32:@9906.4]
  assign active_1_io_input_reset = _T_192 | io_parentAck; // @[Controllers.scala 115:34:@9910.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@9783.4]
  assign done_0_clock = clock; // @[:@9774.4]
  assign done_0_reset = reset; // @[:@9775.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 108:28:@9893.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@9794.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@9784.4]
  assign done_1_clock = clock; // @[:@9777.4]
  assign done_1_reset = reset; // @[:@9778.4]
  assign done_1_io_input_set = done_0_io_output & synchronize; // @[Controllers.scala 117:30:@9917.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@9803.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@9785.4]
  assign iterDone_0_clock = clock; // @[:@9806.4]
  assign iterDone_0_reset = reset; // @[:@9807.4]
  assign iterDone_0_io_input_set = io_doneIn_0 | _T_174; // @[Controllers.scala 107:32:@9889.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@9821.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@9811.4]
  assign iterDone_1_clock = clock; // @[:@9809.4]
  assign iterDone_1_reset = reset; // @[:@9810.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 116:34:@9912.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@9830.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@9812.4]
  assign RetimeWrapper_clock = clock; // @[:@9837.4]
  assign RetimeWrapper_reset = reset; // @[:@9838.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@9840.4]
  assign RetimeWrapper_io_in = io_maskIn_0; // @[package.scala 94:16:@9839.4]
  assign RetimeWrapper_1_clock = clock; // @[:@9850.4]
  assign RetimeWrapper_1_reset = reset; // @[:@9851.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@9853.4]
  assign RetimeWrapper_1_io_in = io_maskIn_1; // @[package.scala 94:16:@9852.4]
  assign RetimeWrapper_2_clock = clock; // @[:@9876.4]
  assign RetimeWrapper_2_reset = reset; // @[:@9877.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@9879.4]
  assign RetimeWrapper_2_io_in = io_maskIn_0; // @[package.scala 94:16:@9878.4]
  assign RetimeWrapper_3_clock = clock; // @[:@9896.4]
  assign RetimeWrapper_3_reset = reset; // @[:@9897.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@9899.4]
  assign RetimeWrapper_3_io_in = synchronize & iterDone_0_io_output; // @[package.scala 94:16:@9898.4]
  assign RetimeWrapper_4_clock = clock; // @[:@9945.4]
  assign RetimeWrapper_4_reset = reset; // @[:@9946.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@9948.4]
  assign RetimeWrapper_4_io_in = _T_224 | io_parentAck; // @[package.scala 94:16:@9947.4]
  assign RetimeWrapper_5_clock = clock; // @[:@9962.4]
  assign RetimeWrapper_5_reset = reset; // @[:@9963.4]
  assign RetimeWrapper_5_io_flow = io_enable; // @[package.scala 95:18:@9965.4]
  assign RetimeWrapper_5_io_in = allDone & _T_237; // @[package.scala 94:16:@9964.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_223 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_237 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_223 <= 1'h0;
    end else begin
      _T_223 <= _T_220;
    end
    if (reset) begin
      _T_237 <= 1'h0;
    end else begin
      _T_237 <= _T_220;
    end
  end
endmodule
module RetimeWrapper_96( // @[:@10439.2]
  input         clock, // @[:@10440.4]
  input         reset, // @[:@10441.4]
  input         io_flow, // @[:@10442.4]
  input  [31:0] io_in, // @[:@10442.4]
  output [31:0] io_out // @[:@10442.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@10444.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@10444.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@10444.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@10444.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@10444.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@10444.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@10444.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@10457.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@10456.4]
  assign sr_init = 32'h1; // @[RetimeShiftRegister.scala 19:16:@10455.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@10454.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@10453.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@10451.4]
endmodule
module NBufCtr( // @[:@10459.2]
  input         clock, // @[:@10460.4]
  input         reset, // @[:@10461.4]
  input         io_input_countUp, // @[:@10462.4]
  input         io_input_enable, // @[:@10462.4]
  output [31:0] io_output_count // @[:@10462.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@10499.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@10499.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@10499.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@10499.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@10499.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@10504.4 package.scala 96:25:@10505.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@10465.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@10466.4]
  wire  _T_21; // @[Counter.scala 49:55:@10467.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@10468.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@10469.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@10470.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@10471.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@10472.4]
  wire  _T_33; // @[Counter.scala 51:52:@10476.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@10477.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@10478.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@10479.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@10480.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@10481.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@10482.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@10483.4]
  wire  _T_45; // @[Counter.scala 52:70:@10484.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@10486.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@10487.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@10488.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@10489.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@10490.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@10491.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@10494.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@10495.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@10497.4]
  RetimeWrapper_96 RetimeWrapper ( // @[package.scala 93:22:@10499.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@10504.4 package.scala 96:25:@10505.4]
  assign _T_18 = {{1'd0}, _T_66}; // @[Counter.scala 49:32:@10465.4]
  assign _T_19 = _T_18[31:0]; // @[Counter.scala 49:32:@10466.4]
  assign _T_21 = _T_19 >= 32'h2; // @[Counter.scala 49:55:@10467.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@10468.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh2); // @[Counter.scala 49:91:@10469.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh2); // @[Counter.scala 49:91:@10470.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@10471.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@10472.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@10476.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@10477.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@10478.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@10479.4]
  assign _T_39 = _T_33 ? 32'h1 : _T_38; // @[Counter.scala 51:47:@10480.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@10481.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@10482.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@10483.4]
  assign _T_45 = _T_43 >= 32'h2; // @[Counter.scala 52:70:@10484.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 52:121:@10486.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 52:121:@10487.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@10488.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@10489.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@10490.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@10491.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@10494.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@10495.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@10497.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@10507.4]
  assign RetimeWrapper_clock = clock; // @[:@10500.4]
  assign RetimeWrapper_reset = reset; // @[:@10501.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@10503.4]
  assign RetimeWrapper_io_in = reset ? 32'h1 : _T_62; // @[package.scala 94:16:@10502.4]
endmodule
module NBufCtr_2( // @[:@10623.2]
  input         clock, // @[:@10624.4]
  input         reset, // @[:@10625.4]
  input         io_input_countUp, // @[:@10626.4]
  input         io_input_enable, // @[:@10626.4]
  output [31:0] io_output_count // @[:@10626.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@10663.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@10663.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@10663.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@10663.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@10663.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@10668.4 package.scala 96:25:@10669.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@10629.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@10630.4]
  wire  _T_21; // @[Counter.scala 49:55:@10631.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@10632.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@10633.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@10634.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@10635.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@10636.4]
  wire  _T_33; // @[Counter.scala 51:52:@10640.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@10641.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@10642.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@10643.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@10644.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@10645.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@10654.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@10655.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@10658.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@10659.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@10661.4]
  RetimeWrapper_96 RetimeWrapper ( // @[package.scala 93:22:@10663.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@10668.4 package.scala 96:25:@10669.4]
  assign _T_18 = _T_66 + 32'h1; // @[Counter.scala 49:32:@10629.4]
  assign _T_19 = _T_66 + 32'h1; // @[Counter.scala 49:32:@10630.4]
  assign _T_21 = _T_19 >= 32'h2; // @[Counter.scala 49:55:@10631.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@10632.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 49:91:@10633.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 49:91:@10634.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@10635.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@10636.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@10640.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@10641.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@10642.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@10643.4]
  assign _T_39 = _T_33 ? 32'h1 : _T_38; // @[Counter.scala 51:47:@10644.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@10645.4]
  assign _T_53 = {{1'd0}, _T_27}; // @[Counter.scala 52:107:@10654.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@10655.4]
  assign _T_58 = _T_21 ? _T_54 : _T_19; // @[Counter.scala 52:45:@10658.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@10659.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@10661.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@10671.4]
  assign RetimeWrapper_clock = clock; // @[:@10664.4]
  assign RetimeWrapper_reset = reset; // @[:@10665.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@10667.4]
  assign RetimeWrapper_io_in = reset ? 32'h1 : _T_62; // @[package.scala 94:16:@10666.4]
endmodule
module NBufController( // @[:@10673.2]
  input        clock, // @[:@10674.4]
  input        reset, // @[:@10675.4]
  input        io_sEn_0, // @[:@10676.4]
  input        io_sEn_1, // @[:@10676.4]
  input        io_sDone_0, // @[:@10676.4]
  input        io_sDone_1, // @[:@10676.4]
  output [2:0] io_statesInW_0, // @[:@10676.4]
  output [2:0] io_statesInR_1 // @[:@10676.4]
);
  wire  sEn_latch_0_clock; // @[NBuffers.scala 21:52:@10678.4]
  wire  sEn_latch_0_reset; // @[NBuffers.scala 21:52:@10678.4]
  wire  sEn_latch_0_io_input_set; // @[NBuffers.scala 21:52:@10678.4]
  wire  sEn_latch_0_io_input_reset; // @[NBuffers.scala 21:52:@10678.4]
  wire  sEn_latch_0_io_input_asyn_reset; // @[NBuffers.scala 21:52:@10678.4]
  wire  sEn_latch_0_io_output; // @[NBuffers.scala 21:52:@10678.4]
  wire  sEn_latch_1_clock; // @[NBuffers.scala 21:52:@10681.4]
  wire  sEn_latch_1_reset; // @[NBuffers.scala 21:52:@10681.4]
  wire  sEn_latch_1_io_input_set; // @[NBuffers.scala 21:52:@10681.4]
  wire  sEn_latch_1_io_input_reset; // @[NBuffers.scala 21:52:@10681.4]
  wire  sEn_latch_1_io_input_asyn_reset; // @[NBuffers.scala 21:52:@10681.4]
  wire  sEn_latch_1_io_output; // @[NBuffers.scala 21:52:@10681.4]
  wire  sDone_latch_0_clock; // @[NBuffers.scala 22:54:@10684.4]
  wire  sDone_latch_0_reset; // @[NBuffers.scala 22:54:@10684.4]
  wire  sDone_latch_0_io_input_set; // @[NBuffers.scala 22:54:@10684.4]
  wire  sDone_latch_0_io_input_reset; // @[NBuffers.scala 22:54:@10684.4]
  wire  sDone_latch_0_io_input_asyn_reset; // @[NBuffers.scala 22:54:@10684.4]
  wire  sDone_latch_0_io_output; // @[NBuffers.scala 22:54:@10684.4]
  wire  sDone_latch_1_clock; // @[NBuffers.scala 22:54:@10687.4]
  wire  sDone_latch_1_reset; // @[NBuffers.scala 22:54:@10687.4]
  wire  sDone_latch_1_io_input_set; // @[NBuffers.scala 22:54:@10687.4]
  wire  sDone_latch_1_io_input_reset; // @[NBuffers.scala 22:54:@10687.4]
  wire  sDone_latch_1_io_input_asyn_reset; // @[NBuffers.scala 22:54:@10687.4]
  wire  sDone_latch_1_io_output; // @[NBuffers.scala 22:54:@10687.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@10694.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@10694.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@10694.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@10694.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@10694.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@10702.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@10702.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@10702.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@10702.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@10702.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@10711.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@10711.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@10711.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@10711.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@10711.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@10719.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@10719.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@10719.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@10719.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@10719.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@10730.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@10730.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@10730.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@10730.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@10730.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@10738.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@10738.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@10738.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@10738.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@10738.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@10755.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@10755.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@10755.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@10755.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@10755.4]
  wire  NBufCtr_clock; // @[NBuffers.scala 40:19:@10776.4]
  wire  NBufCtr_reset; // @[NBuffers.scala 40:19:@10776.4]
  wire  NBufCtr_io_input_countUp; // @[NBuffers.scala 40:19:@10776.4]
  wire  NBufCtr_io_input_enable; // @[NBuffers.scala 40:19:@10776.4]
  wire [31:0] NBufCtr_io_output_count; // @[NBuffers.scala 40:19:@10776.4]
  wire  statesInR_0_clock; // @[NBuffers.scala 50:19:@10787.4]
  wire  statesInR_0_reset; // @[NBuffers.scala 50:19:@10787.4]
  wire  statesInR_0_io_input_countUp; // @[NBuffers.scala 50:19:@10787.4]
  wire  statesInR_0_io_input_enable; // @[NBuffers.scala 50:19:@10787.4]
  wire [31:0] statesInR_0_io_output_count; // @[NBuffers.scala 50:19:@10787.4]
  wire  statesInR_1_clock; // @[NBuffers.scala 50:19:@10798.4]
  wire  statesInR_1_reset; // @[NBuffers.scala 50:19:@10798.4]
  wire  statesInR_1_io_input_countUp; // @[NBuffers.scala 50:19:@10798.4]
  wire  statesInR_1_io_input_enable; // @[NBuffers.scala 50:19:@10798.4]
  wire [31:0] statesInR_1_io_output_count; // @[NBuffers.scala 50:19:@10798.4]
  wire  _T_33; // @[NBuffers.scala 26:46:@10691.4]
  wire  _T_48; // @[NBuffers.scala 26:46:@10727.4]
  wire  anyEnabled; // @[NBuffers.scala 33:64:@10763.4]
  wire  _T_62; // @[NBuffers.scala 34:124:@10764.4]
  wire  _T_63; // @[NBuffers.scala 34:104:@10765.4]
  wire  _T_64; // @[NBuffers.scala 34:124:@10766.4]
  wire  _T_65; // @[NBuffers.scala 34:104:@10767.4]
  wire  _T_66; // @[NBuffers.scala 34:150:@10768.4]
  wire  _T_67; // @[NBuffers.scala 34:154:@10769.4]
  wire  _T_69; // @[package.scala 100:49:@10770.4]
  reg  _T_72; // @[package.scala 48:56:@10771.4]
  reg [31:0] _RAND_0;
  SRFF sEn_latch_0 ( // @[NBuffers.scala 21:52:@10678.4]
    .clock(sEn_latch_0_clock),
    .reset(sEn_latch_0_reset),
    .io_input_set(sEn_latch_0_io_input_set),
    .io_input_reset(sEn_latch_0_io_input_reset),
    .io_input_asyn_reset(sEn_latch_0_io_input_asyn_reset),
    .io_output(sEn_latch_0_io_output)
  );
  SRFF sEn_latch_1 ( // @[NBuffers.scala 21:52:@10681.4]
    .clock(sEn_latch_1_clock),
    .reset(sEn_latch_1_reset),
    .io_input_set(sEn_latch_1_io_input_set),
    .io_input_reset(sEn_latch_1_io_input_reset),
    .io_input_asyn_reset(sEn_latch_1_io_input_asyn_reset),
    .io_output(sEn_latch_1_io_output)
  );
  SRFF sDone_latch_0 ( // @[NBuffers.scala 22:54:@10684.4]
    .clock(sDone_latch_0_clock),
    .reset(sDone_latch_0_reset),
    .io_input_set(sDone_latch_0_io_input_set),
    .io_input_reset(sDone_latch_0_io_input_reset),
    .io_input_asyn_reset(sDone_latch_0_io_input_asyn_reset),
    .io_output(sDone_latch_0_io_output)
  );
  SRFF sDone_latch_1 ( // @[NBuffers.scala 22:54:@10687.4]
    .clock(sDone_latch_1_clock),
    .reset(sDone_latch_1_reset),
    .io_input_set(sDone_latch_1_io_input_set),
    .io_input_reset(sDone_latch_1_io_input_reset),
    .io_input_asyn_reset(sDone_latch_1_io_input_asyn_reset),
    .io_output(sDone_latch_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@10694.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@10702.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@10711.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@10719.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@10730.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@10738.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@10747.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@10755.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  NBufCtr NBufCtr ( // @[NBuffers.scala 40:19:@10776.4]
    .clock(NBufCtr_clock),
    .reset(NBufCtr_reset),
    .io_input_countUp(NBufCtr_io_input_countUp),
    .io_input_enable(NBufCtr_io_input_enable),
    .io_output_count(NBufCtr_io_output_count)
  );
  NBufCtr statesInR_0 ( // @[NBuffers.scala 50:19:@10787.4]
    .clock(statesInR_0_clock),
    .reset(statesInR_0_reset),
    .io_input_countUp(statesInR_0_io_input_countUp),
    .io_input_enable(statesInR_0_io_input_enable),
    .io_output_count(statesInR_0_io_output_count)
  );
  NBufCtr_2 statesInR_1 ( // @[NBuffers.scala 50:19:@10798.4]
    .clock(statesInR_1_clock),
    .reset(statesInR_1_reset),
    .io_input_countUp(statesInR_1_io_input_countUp),
    .io_input_enable(statesInR_1_io_input_enable),
    .io_output_count(statesInR_1_io_output_count)
  );
  assign _T_33 = io_sDone_0 == 1'h0; // @[NBuffers.scala 26:46:@10691.4]
  assign _T_48 = io_sDone_1 == 1'h0; // @[NBuffers.scala 26:46:@10727.4]
  assign anyEnabled = sEn_latch_0_io_output | sEn_latch_1_io_output; // @[NBuffers.scala 33:64:@10763.4]
  assign _T_62 = sDone_latch_0_io_output | io_sDone_0; // @[NBuffers.scala 34:124:@10764.4]
  assign _T_63 = sEn_latch_0_io_output == _T_62; // @[NBuffers.scala 34:104:@10765.4]
  assign _T_64 = sDone_latch_1_io_output | io_sDone_1; // @[NBuffers.scala 34:124:@10766.4]
  assign _T_65 = sEn_latch_1_io_output == _T_64; // @[NBuffers.scala 34:104:@10767.4]
  assign _T_66 = _T_63 & _T_65; // @[NBuffers.scala 34:150:@10768.4]
  assign _T_67 = _T_66 & anyEnabled; // @[NBuffers.scala 34:154:@10769.4]
  assign _T_69 = _T_67 == 1'h0; // @[package.scala 100:49:@10770.4]
  assign io_statesInW_0 = NBufCtr_io_output_count[2:0]; // @[NBuffers.scala 44:21:@10786.4]
  assign io_statesInR_1 = statesInR_1_io_output_count[2:0]; // @[NBuffers.scala 54:21:@10808.4]
  assign sEn_latch_0_clock = clock; // @[:@10679.4]
  assign sEn_latch_0_reset = reset; // @[:@10680.4]
  assign sEn_latch_0_io_input_set = io_sEn_0 & _T_33; // @[NBuffers.scala 26:31:@10693.4]
  assign sEn_latch_0_io_input_reset = RetimeWrapper_io_out; // @[NBuffers.scala 27:33:@10701.4]
  assign sEn_latch_0_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[NBuffers.scala 28:38:@10709.4]
  assign sEn_latch_1_clock = clock; // @[:@10682.4]
  assign sEn_latch_1_reset = reset; // @[:@10683.4]
  assign sEn_latch_1_io_input_set = io_sEn_1 & _T_48; // @[NBuffers.scala 26:31:@10729.4]
  assign sEn_latch_1_io_input_reset = RetimeWrapper_4_io_out; // @[NBuffers.scala 27:33:@10737.4]
  assign sEn_latch_1_io_input_asyn_reset = RetimeWrapper_5_io_out; // @[NBuffers.scala 28:38:@10745.4]
  assign sDone_latch_0_clock = clock; // @[:@10685.4]
  assign sDone_latch_0_reset = reset; // @[:@10686.4]
  assign sDone_latch_0_io_input_set = io_sDone_0; // @[NBuffers.scala 29:33:@10710.4]
  assign sDone_latch_0_io_input_reset = RetimeWrapper_2_io_out; // @[NBuffers.scala 30:35:@10718.4]
  assign sDone_latch_0_io_input_asyn_reset = RetimeWrapper_3_io_out; // @[NBuffers.scala 31:40:@10726.4]
  assign sDone_latch_1_clock = clock; // @[:@10688.4]
  assign sDone_latch_1_reset = reset; // @[:@10689.4]
  assign sDone_latch_1_io_input_set = io_sDone_1; // @[NBuffers.scala 29:33:@10746.4]
  assign sDone_latch_1_io_input_reset = RetimeWrapper_6_io_out; // @[NBuffers.scala 30:35:@10754.4]
  assign sDone_latch_1_io_input_asyn_reset = RetimeWrapper_7_io_out; // @[NBuffers.scala 31:40:@10762.4]
  assign RetimeWrapper_clock = clock; // @[:@10695.4]
  assign RetimeWrapper_reset = reset; // @[:@10696.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@10698.4]
  assign RetimeWrapper_io_in = _T_67 & _T_72; // @[package.scala 94:16:@10697.4]
  assign RetimeWrapper_1_clock = clock; // @[:@10703.4]
  assign RetimeWrapper_1_reset = reset; // @[:@10704.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@10706.4]
  assign RetimeWrapper_1_io_in = reset; // @[package.scala 94:16:@10705.4]
  assign RetimeWrapper_2_clock = clock; // @[:@10712.4]
  assign RetimeWrapper_2_reset = reset; // @[:@10713.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@10715.4]
  assign RetimeWrapper_2_io_in = _T_67 & _T_72; // @[package.scala 94:16:@10714.4]
  assign RetimeWrapper_3_clock = clock; // @[:@10720.4]
  assign RetimeWrapper_3_reset = reset; // @[:@10721.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@10723.4]
  assign RetimeWrapper_3_io_in = reset; // @[package.scala 94:16:@10722.4]
  assign RetimeWrapper_4_clock = clock; // @[:@10731.4]
  assign RetimeWrapper_4_reset = reset; // @[:@10732.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@10734.4]
  assign RetimeWrapper_4_io_in = _T_67 & _T_72; // @[package.scala 94:16:@10733.4]
  assign RetimeWrapper_5_clock = clock; // @[:@10739.4]
  assign RetimeWrapper_5_reset = reset; // @[:@10740.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@10742.4]
  assign RetimeWrapper_5_io_in = reset; // @[package.scala 94:16:@10741.4]
  assign RetimeWrapper_6_clock = clock; // @[:@10748.4]
  assign RetimeWrapper_6_reset = reset; // @[:@10749.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@10751.4]
  assign RetimeWrapper_6_io_in = _T_67 & _T_72; // @[package.scala 94:16:@10750.4]
  assign RetimeWrapper_7_clock = clock; // @[:@10756.4]
  assign RetimeWrapper_7_reset = reset; // @[:@10757.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@10759.4]
  assign RetimeWrapper_7_io_in = reset; // @[package.scala 94:16:@10758.4]
  assign NBufCtr_clock = clock; // @[:@10777.4]
  assign NBufCtr_reset = reset; // @[:@10778.4]
  assign NBufCtr_io_input_countUp = 1'h0; // @[NBuffers.scala 43:24:@10785.4]
  assign NBufCtr_io_input_enable = _T_67 & _T_72; // @[NBuffers.scala 42:23:@10784.4]
  assign statesInR_0_clock = clock; // @[:@10788.4]
  assign statesInR_0_reset = reset; // @[:@10789.4]
  assign statesInR_0_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@10796.4]
  assign statesInR_0_io_input_enable = _T_67 & _T_72; // @[NBuffers.scala 52:23:@10795.4]
  assign statesInR_1_clock = clock; // @[:@10799.4]
  assign statesInR_1_reset = reset; // @[:@10800.4]
  assign statesInR_1_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@10807.4]
  assign statesInR_1_io_input_enable = _T_67 & _T_72; // @[NBuffers.scala 52:23:@10806.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_72 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_72 <= 1'h0;
    end else begin
      _T_72 <= _T_69;
    end
  end
endmodule
module NBuf( // @[:@10860.2]
  input         clock, // @[:@10861.4]
  input         reset, // @[:@10862.4]
  output [31:0] io_rPort_0_output_0, // @[:@10863.4]
  input  [31:0] io_wPort_0_data_0, // @[:@10863.4]
  input         io_wPort_0_reset, // @[:@10863.4]
  input         io_wPort_0_en_0, // @[:@10863.4]
  input         io_sEn_0, // @[:@10863.4]
  input         io_sEn_1, // @[:@10863.4]
  input         io_sDone_0, // @[:@10863.4]
  input         io_sDone_1 // @[:@10863.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@10871.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@10871.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@10871.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@10871.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@10871.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@10871.4]
  wire [2:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@10871.4]
  wire [2:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@10871.4]
  wire  FF_clock; // @[NBuffers.scala 146:23:@10878.4]
  wire  FF_reset; // @[NBuffers.scala 146:23:@10878.4]
  wire [31:0] FF_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@10878.4]
  wire [31:0] FF_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@10878.4]
  wire  FF_io_wPort_0_reset; // @[NBuffers.scala 146:23:@10878.4]
  wire  FF_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@10878.4]
  wire  FF_1_clock; // @[NBuffers.scala 146:23:@10894.4]
  wire  FF_1_reset; // @[NBuffers.scala 146:23:@10894.4]
  wire [31:0] FF_1_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@10894.4]
  wire [31:0] FF_1_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@10894.4]
  wire  FF_1_io_wPort_0_reset; // @[NBuffers.scala 146:23:@10894.4]
  wire  FF_1_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@10894.4]
  wire  _T_106; // @[NBuffers.scala 153:105:@10912.4]
  wire  _T_110; // @[NBuffers.scala 157:92:@10922.4]
  wire  _T_113; // @[NBuffers.scala 153:105:@10928.4]
  wire  _T_117; // @[NBuffers.scala 157:92:@10938.4]
  wire [31:0] _T_125; // @[Mux.scala 19:72:@10946.4]
  wire [31:0] _T_127; // @[Mux.scala 19:72:@10947.4]
  NBufController ctrl ( // @[NBuffers.scala 83:20:@10871.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1)
  );
  FF FF ( // @[NBuffers.scala 146:23:@10878.4]
    .clock(FF_clock),
    .reset(FF_reset),
    .io_rPort_0_output_0(FF_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_io_wPort_0_en_0)
  );
  FF FF_1 ( // @[NBuffers.scala 146:23:@10894.4]
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_rPort_0_output_0(FF_1_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_1_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_1_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_1_io_wPort_0_en_0)
  );
  assign _T_106 = ctrl_io_statesInW_0 == 3'h0; // @[NBuffers.scala 153:105:@10912.4]
  assign _T_110 = ctrl_io_statesInR_1 == 3'h0; // @[NBuffers.scala 157:92:@10922.4]
  assign _T_113 = ctrl_io_statesInW_0 == 3'h1; // @[NBuffers.scala 153:105:@10928.4]
  assign _T_117 = ctrl_io_statesInR_1 == 3'h1; // @[NBuffers.scala 157:92:@10938.4]
  assign _T_125 = _T_110 ? FF_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@10946.4]
  assign _T_127 = _T_117 ? FF_1_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@10947.4]
  assign io_rPort_0_output_0 = _T_125 | _T_127; // @[NBuffers.scala 163:66:@10951.4]
  assign ctrl_clock = clock; // @[:@10872.4]
  assign ctrl_reset = reset; // @[:@10873.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@10874.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@10876.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@10875.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@10877.4]
  assign FF_clock = clock; // @[:@10879.4]
  assign FF_reset = reset; // @[:@10880.4]
  assign FF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@10915.4]
  assign FF_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@10916.4]
  assign FF_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_106; // @[MemPrimitives.scala 37:29:@10921.4]
  assign FF_1_clock = clock; // @[:@10895.4]
  assign FF_1_reset = reset; // @[:@10896.4]
  assign FF_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@10931.4]
  assign FF_1_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@10932.4]
  assign FF_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_113; // @[MemPrimitives.scala 37:29:@10937.4]
endmodule
module b542_chain( // @[:@10953.2]
  input         clock, // @[:@10954.4]
  input         reset, // @[:@10955.4]
  output [31:0] io_rPort_0_output_0, // @[:@10956.4]
  input  [31:0] io_wPort_0_data_0, // @[:@10956.4]
  input         io_wPort_0_reset, // @[:@10956.4]
  input         io_wPort_0_en_0, // @[:@10956.4]
  input         io_sEn_0, // @[:@10956.4]
  input         io_sEn_1, // @[:@10956.4]
  input         io_sDone_0, // @[:@10956.4]
  input         io_sDone_1 // @[:@10956.4]
);
  wire  nbufFF_clock; // @[NBuffers.scala 298:22:@10964.4]
  wire  nbufFF_reset; // @[NBuffers.scala 298:22:@10964.4]
  wire [31:0] nbufFF_io_rPort_0_output_0; // @[NBuffers.scala 298:22:@10964.4]
  wire [31:0] nbufFF_io_wPort_0_data_0; // @[NBuffers.scala 298:22:@10964.4]
  wire  nbufFF_io_wPort_0_reset; // @[NBuffers.scala 298:22:@10964.4]
  wire  nbufFF_io_wPort_0_en_0; // @[NBuffers.scala 298:22:@10964.4]
  wire  nbufFF_io_sEn_0; // @[NBuffers.scala 298:22:@10964.4]
  wire  nbufFF_io_sEn_1; // @[NBuffers.scala 298:22:@10964.4]
  wire  nbufFF_io_sDone_0; // @[NBuffers.scala 298:22:@10964.4]
  wire  nbufFF_io_sDone_1; // @[NBuffers.scala 298:22:@10964.4]
  NBuf nbufFF ( // @[NBuffers.scala 298:22:@10964.4]
    .clock(nbufFF_clock),
    .reset(nbufFF_reset),
    .io_rPort_0_output_0(nbufFF_io_rPort_0_output_0),
    .io_wPort_0_data_0(nbufFF_io_wPort_0_data_0),
    .io_wPort_0_reset(nbufFF_io_wPort_0_reset),
    .io_wPort_0_en_0(nbufFF_io_wPort_0_en_0),
    .io_sEn_0(nbufFF_io_sEn_0),
    .io_sEn_1(nbufFF_io_sEn_1),
    .io_sDone_0(nbufFF_io_sDone_0),
    .io_sDone_1(nbufFF_io_sDone_1)
  );
  assign io_rPort_0_output_0 = nbufFF_io_rPort_0_output_0; // @[NBuffers.scala 299:6:@10986.4]
  assign nbufFF_clock = clock; // @[:@10965.4]
  assign nbufFF_reset = reset; // @[:@10966.4]
  assign nbufFF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[NBuffers.scala 299:6:@10983.4]
  assign nbufFF_io_wPort_0_reset = io_wPort_0_reset; // @[NBuffers.scala 299:6:@10982.4]
  assign nbufFF_io_wPort_0_en_0 = io_wPort_0_en_0; // @[NBuffers.scala 299:6:@10979.4]
  assign nbufFF_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 299:6:@10969.4]
  assign nbufFF_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 299:6:@10970.4]
  assign nbufFF_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 299:6:@10967.4]
  assign nbufFF_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 299:6:@10968.4]
endmodule
module FF_9( // @[:@11751.2]
  input   clock, // @[:@11752.4]
  input   reset, // @[:@11753.4]
  output  io_rPort_0_output_0, // @[:@11754.4]
  input   io_wPort_0_data_0, // @[:@11754.4]
  input   io_wPort_0_reset, // @[:@11754.4]
  input   io_wPort_0_en_0 // @[:@11754.4]
);
  reg  ff; // @[MemPrimitives.scala 321:19:@11769.4]
  reg [31:0] _RAND_0;
  wire  _T_68; // @[MemPrimitives.scala 325:32:@11771.4]
  wire  _T_69; // @[MemPrimitives.scala 325:12:@11772.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@11771.4]
  assign _T_69 = io_wPort_0_reset ? 1'h0 : _T_68; // @[MemPrimitives.scala 325:12:@11772.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@11774.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 1'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 1'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module NBuf_1( // @[:@11801.2]
  input   clock, // @[:@11802.4]
  input   reset, // @[:@11803.4]
  output  io_rPort_0_output_0, // @[:@11804.4]
  input   io_wPort_0_data_0, // @[:@11804.4]
  input   io_wPort_0_reset, // @[:@11804.4]
  input   io_wPort_0_en_0, // @[:@11804.4]
  input   io_sEn_0, // @[:@11804.4]
  input   io_sEn_1, // @[:@11804.4]
  input   io_sDone_0, // @[:@11804.4]
  input   io_sDone_1 // @[:@11804.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@11812.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@11812.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@11812.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@11812.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@11812.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@11812.4]
  wire [2:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@11812.4]
  wire [2:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@11812.4]
  wire  FF_clock; // @[NBuffers.scala 146:23:@11819.4]
  wire  FF_reset; // @[NBuffers.scala 146:23:@11819.4]
  wire  FF_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@11819.4]
  wire  FF_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@11819.4]
  wire  FF_io_wPort_0_reset; // @[NBuffers.scala 146:23:@11819.4]
  wire  FF_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@11819.4]
  wire  FF_1_clock; // @[NBuffers.scala 146:23:@11835.4]
  wire  FF_1_reset; // @[NBuffers.scala 146:23:@11835.4]
  wire  FF_1_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@11835.4]
  wire  FF_1_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@11835.4]
  wire  FF_1_io_wPort_0_reset; // @[NBuffers.scala 146:23:@11835.4]
  wire  FF_1_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@11835.4]
  wire  _T_106; // @[NBuffers.scala 153:105:@11853.4]
  wire  _T_110; // @[NBuffers.scala 157:92:@11863.4]
  wire  _T_113; // @[NBuffers.scala 153:105:@11869.4]
  wire  _T_117; // @[NBuffers.scala 157:92:@11879.4]
  wire  _T_125; // @[Mux.scala 19:72:@11887.4]
  wire  _T_127; // @[Mux.scala 19:72:@11888.4]
  NBufController ctrl ( // @[NBuffers.scala 83:20:@11812.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1)
  );
  FF_9 FF ( // @[NBuffers.scala 146:23:@11819.4]
    .clock(FF_clock),
    .reset(FF_reset),
    .io_rPort_0_output_0(FF_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_io_wPort_0_en_0)
  );
  FF_9 FF_1 ( // @[NBuffers.scala 146:23:@11835.4]
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_rPort_0_output_0(FF_1_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_1_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_1_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_1_io_wPort_0_en_0)
  );
  assign _T_106 = ctrl_io_statesInW_0 == 3'h0; // @[NBuffers.scala 153:105:@11853.4]
  assign _T_110 = ctrl_io_statesInR_1 == 3'h0; // @[NBuffers.scala 157:92:@11863.4]
  assign _T_113 = ctrl_io_statesInW_0 == 3'h1; // @[NBuffers.scala 153:105:@11869.4]
  assign _T_117 = ctrl_io_statesInR_1 == 3'h1; // @[NBuffers.scala 157:92:@11879.4]
  assign _T_125 = _T_110 ? FF_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@11887.4]
  assign _T_127 = _T_117 ? FF_1_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@11888.4]
  assign io_rPort_0_output_0 = _T_125 | _T_127; // @[NBuffers.scala 163:66:@11892.4]
  assign ctrl_clock = clock; // @[:@11813.4]
  assign ctrl_reset = reset; // @[:@11814.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@11815.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@11817.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@11816.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@11818.4]
  assign FF_clock = clock; // @[:@11820.4]
  assign FF_reset = reset; // @[:@11821.4]
  assign FF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@11856.4]
  assign FF_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@11857.4]
  assign FF_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_106; // @[MemPrimitives.scala 37:29:@11862.4]
  assign FF_1_clock = clock; // @[:@11836.4]
  assign FF_1_reset = reset; // @[:@11837.4]
  assign FF_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@11872.4]
  assign FF_1_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@11873.4]
  assign FF_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_113; // @[MemPrimitives.scala 37:29:@11878.4]
endmodule
module b543_chain( // @[:@11894.2]
  input   clock, // @[:@11895.4]
  input   reset, // @[:@11896.4]
  output  io_rPort_0_output_0, // @[:@11897.4]
  input   io_wPort_0_data_0, // @[:@11897.4]
  input   io_wPort_0_reset, // @[:@11897.4]
  input   io_wPort_0_en_0, // @[:@11897.4]
  input   io_sEn_0, // @[:@11897.4]
  input   io_sEn_1, // @[:@11897.4]
  input   io_sDone_0, // @[:@11897.4]
  input   io_sDone_1 // @[:@11897.4]
);
  wire  nbufFF_clock; // @[NBuffers.scala 298:22:@11905.4]
  wire  nbufFF_reset; // @[NBuffers.scala 298:22:@11905.4]
  wire  nbufFF_io_rPort_0_output_0; // @[NBuffers.scala 298:22:@11905.4]
  wire  nbufFF_io_wPort_0_data_0; // @[NBuffers.scala 298:22:@11905.4]
  wire  nbufFF_io_wPort_0_reset; // @[NBuffers.scala 298:22:@11905.4]
  wire  nbufFF_io_wPort_0_en_0; // @[NBuffers.scala 298:22:@11905.4]
  wire  nbufFF_io_sEn_0; // @[NBuffers.scala 298:22:@11905.4]
  wire  nbufFF_io_sEn_1; // @[NBuffers.scala 298:22:@11905.4]
  wire  nbufFF_io_sDone_0; // @[NBuffers.scala 298:22:@11905.4]
  wire  nbufFF_io_sDone_1; // @[NBuffers.scala 298:22:@11905.4]
  NBuf_1 nbufFF ( // @[NBuffers.scala 298:22:@11905.4]
    .clock(nbufFF_clock),
    .reset(nbufFF_reset),
    .io_rPort_0_output_0(nbufFF_io_rPort_0_output_0),
    .io_wPort_0_data_0(nbufFF_io_wPort_0_data_0),
    .io_wPort_0_reset(nbufFF_io_wPort_0_reset),
    .io_wPort_0_en_0(nbufFF_io_wPort_0_en_0),
    .io_sEn_0(nbufFF_io_sEn_0),
    .io_sEn_1(nbufFF_io_sEn_1),
    .io_sDone_0(nbufFF_io_sDone_0),
    .io_sDone_1(nbufFF_io_sDone_1)
  );
  assign io_rPort_0_output_0 = nbufFF_io_rPort_0_output_0; // @[NBuffers.scala 299:6:@11927.4]
  assign nbufFF_clock = clock; // @[:@11906.4]
  assign nbufFF_reset = reset; // @[:@11907.4]
  assign nbufFF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[NBuffers.scala 299:6:@11924.4]
  assign nbufFF_io_wPort_0_reset = io_wPort_0_reset; // @[NBuffers.scala 299:6:@11923.4]
  assign nbufFF_io_wPort_0_en_0 = io_wPort_0_en_0; // @[NBuffers.scala 299:6:@11920.4]
  assign nbufFF_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 299:6:@11910.4]
  assign nbufFF_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 299:6:@11911.4]
  assign nbufFF_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 299:6:@11908.4]
  assign nbufFF_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 299:6:@11909.4]
endmodule
module SRAM_4( // @[:@11981.2]
  input         clock, // @[:@11982.4]
  input         reset, // @[:@11983.4]
  input  [1:0]  io_raddr, // @[:@11984.4]
  input         io_wen, // @[:@11984.4]
  input  [1:0]  io_waddr, // @[:@11984.4]
  input  [31:0] io_wdata, // @[:@11984.4]
  output [31:0] io_rdata, // @[:@11984.4]
  input         io_backpressure // @[:@11984.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@11986.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@11986.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@11986.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@11986.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@11986.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@11986.4]
  wire [1:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@11986.4]
  wire [1:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@11986.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@11986.4]
  wire  _T_19; // @[SRAM.scala 182:49:@12004.4]
  wire  _T_20; // @[SRAM.scala 182:37:@12005.4]
  reg  _T_23; // @[SRAM.scala 182:29:@12006.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@12008.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(3), .AWIDTH(2)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@11986.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@12004.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@12005.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@12013.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@12000.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@12001.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@11998.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@12003.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@12002.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@11999.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@11997.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@11996.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_112( // @[:@12027.2]
  input        clock, // @[:@12028.4]
  input        reset, // @[:@12029.4]
  input        io_flow, // @[:@12030.4]
  input  [1:0] io_in, // @[:@12030.4]
  output [1:0] io_out // @[:@12030.4]
);
  wire [1:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12032.4]
  wire [1:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12032.4]
  wire [1:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12032.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12032.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12032.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12032.4]
  RetimeShiftRegister #(.WIDTH(2), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@12032.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12045.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12044.4]
  assign sr_init = 2'h0; // @[RetimeShiftRegister.scala 19:16:@12043.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12042.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12041.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12039.4]
endmodule
module Mem1D_5( // @[:@12047.2]
  input         clock, // @[:@12048.4]
  input         reset, // @[:@12049.4]
  input  [1:0]  io_r_ofs_0, // @[:@12050.4]
  input         io_r_backpressure, // @[:@12050.4]
  input  [1:0]  io_w_ofs_0, // @[:@12050.4]
  input  [31:0] io_w_data_0, // @[:@12050.4]
  input         io_w_en_0, // @[:@12050.4]
  output [31:0] io_output // @[:@12050.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 753:21:@12054.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 753:21:@12054.4]
  wire [1:0] SRAM_io_raddr; // @[MemPrimitives.scala 753:21:@12054.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 753:21:@12054.4]
  wire [1:0] SRAM_io_waddr; // @[MemPrimitives.scala 753:21:@12054.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 753:21:@12054.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 753:21:@12054.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 753:21:@12054.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@12057.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@12057.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@12057.4]
  wire [1:0] RetimeWrapper_io_in; // @[package.scala 93:22:@12057.4]
  wire [1:0] RetimeWrapper_io_out; // @[package.scala 93:22:@12057.4]
  SRAM_4 SRAM ( // @[MemPrimitives.scala 753:21:@12054.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_112 RetimeWrapper ( // @[package.scala 93:22:@12057.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 760:17:@12070.4]
  assign SRAM_clock = clock; // @[:@12055.4]
  assign SRAM_reset = reset; // @[:@12056.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 754:37:@12064.4]
  assign SRAM_io_wen = io_w_en_0; // @[MemPrimitives.scala 757:22:@12067.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 756:22:@12065.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 758:22:@12068.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 759:30:@12069.4]
  assign RetimeWrapper_clock = clock; // @[:@12058.4]
  assign RetimeWrapper_reset = reset; // @[:@12059.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@12061.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@12060.4]
endmodule
module x544_accum_0( // @[:@12111.2]
  input         clock, // @[:@12112.4]
  input         reset, // @[:@12113.4]
  input  [1:0]  io_rPort_0_ofs_0, // @[:@12114.4]
  input         io_rPort_0_en_0, // @[:@12114.4]
  output [31:0] io_rPort_0_output_0, // @[:@12114.4]
  input  [1:0]  io_wPort_0_ofs_0, // @[:@12114.4]
  input  [31:0] io_wPort_0_data_0, // @[:@12114.4]
  input         io_wPort_0_en_0 // @[:@12114.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@12129.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@12129.4]
  wire [1:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12129.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12129.4]
  wire [1:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12129.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@12129.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@12129.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@12129.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@12155.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@12155.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@12169.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@12169.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@12169.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@12169.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@12169.4]
  wire [34:0] _T_70; // @[Cat.scala 30:58:@12147.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@12159.4]
  wire [3:0] _T_78; // @[Cat.scala 30:58:@12161.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@12129.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@12155.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@12169.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_70 = {io_wPort_0_en_0,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12147.4]
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@12159.4]
  assign _T_78 = {_T_76,1'h1,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12161.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@12176.4]
  assign Mem1D_clock = clock; // @[:@12130.4]
  assign Mem1D_reset = reset; // @[:@12131.4]
  assign Mem1D_io_r_ofs_0 = _T_78[1:0]; // @[MemPrimitives.scala 131:28:@12165.4]
  assign Mem1D_io_r_backpressure = _T_78[2]; // @[MemPrimitives.scala 132:32:@12166.4]
  assign Mem1D_io_w_ofs_0 = _T_70[1:0]; // @[MemPrimitives.scala 94:28:@12151.4]
  assign Mem1D_io_w_data_0 = _T_70[33:2]; // @[MemPrimitives.scala 95:29:@12152.4]
  assign Mem1D_io_w_en_0 = _T_70[34]; // @[MemPrimitives.scala 96:27:@12153.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@12158.4]
  assign RetimeWrapper_clock = clock; // @[:@12170.4]
  assign RetimeWrapper_reset = reset; // @[:@12171.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@12173.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@12172.4]
endmodule
module x545_accum_1( // @[:@13295.2]
  input         clock, // @[:@13296.4]
  input         reset, // @[:@13297.4]
  input  [1:0]  io_rPort_0_ofs_0, // @[:@13298.4]
  input         io_rPort_0_en_0, // @[:@13298.4]
  output [31:0] io_rPort_0_output_0, // @[:@13298.4]
  input  [1:0]  io_wPort_0_ofs_0, // @[:@13298.4]
  input  [31:0] io_wPort_0_data_0, // @[:@13298.4]
  input         io_wPort_0_en_0, // @[:@13298.4]
  input         io_sEn_0, // @[:@13298.4]
  input         io_sEn_1, // @[:@13298.4]
  input         io_sDone_0, // @[:@13298.4]
  input         io_sDone_1 // @[:@13298.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@13307.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@13307.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@13307.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@13307.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@13307.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@13307.4]
  wire [2:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@13307.4]
  wire [2:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@13307.4]
  wire  SRAM_clock; // @[NBuffers.scala 94:23:@13314.4]
  wire  SRAM_reset; // @[NBuffers.scala 94:23:@13314.4]
  wire [1:0] SRAM_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@13314.4]
  wire  SRAM_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@13314.4]
  wire [31:0] SRAM_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@13314.4]
  wire [1:0] SRAM_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@13314.4]
  wire [31:0] SRAM_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@13314.4]
  wire  SRAM_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@13314.4]
  wire  SRAM_1_clock; // @[NBuffers.scala 94:23:@13330.4]
  wire  SRAM_1_reset; // @[NBuffers.scala 94:23:@13330.4]
  wire [1:0] SRAM_1_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@13330.4]
  wire  SRAM_1_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@13330.4]
  wire [31:0] SRAM_1_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@13330.4]
  wire [1:0] SRAM_1_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@13330.4]
  wire [31:0] SRAM_1_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@13330.4]
  wire  SRAM_1_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@13330.4]
  wire  _T_110; // @[NBuffers.scala 104:105:@13346.4]
  wire  _T_114; // @[NBuffers.scala 108:92:@13356.4]
  wire  _T_117; // @[NBuffers.scala 104:105:@13362.4]
  wire  _T_121; // @[NBuffers.scala 108:92:@13372.4]
  wire [31:0] _T_129; // @[Mux.scala 19:72:@13380.4]
  wire [31:0] _T_131; // @[Mux.scala 19:72:@13381.4]
  NBufController ctrl ( // @[NBuffers.scala 83:20:@13307.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1)
  );
  x544_accum_0 SRAM ( // @[NBuffers.scala 94:23:@13314.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_rPort_0_ofs_0(SRAM_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_io_rPort_0_en_0),
    .io_rPort_0_output_0(SRAM_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(SRAM_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_io_wPort_0_en_0)
  );
  x544_accum_0 SRAM_1 ( // @[NBuffers.scala 94:23:@13330.4]
    .clock(SRAM_1_clock),
    .reset(SRAM_1_reset),
    .io_rPort_0_ofs_0(SRAM_1_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_1_io_rPort_0_en_0),
    .io_rPort_0_output_0(SRAM_1_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(SRAM_1_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_1_io_wPort_0_en_0)
  );
  assign _T_110 = ctrl_io_statesInW_0 == 3'h0; // @[NBuffers.scala 104:105:@13346.4]
  assign _T_114 = ctrl_io_statesInR_1 == 3'h0; // @[NBuffers.scala 108:92:@13356.4]
  assign _T_117 = ctrl_io_statesInW_0 == 3'h1; // @[NBuffers.scala 104:105:@13362.4]
  assign _T_121 = ctrl_io_statesInR_1 == 3'h1; // @[NBuffers.scala 108:92:@13372.4]
  assign _T_129 = _T_114 ? SRAM_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@13380.4]
  assign _T_131 = _T_121 ? SRAM_1_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@13381.4]
  assign io_rPort_0_output_0 = _T_129 | _T_131; // @[NBuffers.scala 115:66:@13385.4]
  assign ctrl_clock = clock; // @[:@13308.4]
  assign ctrl_reset = reset; // @[:@13309.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@13310.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@13312.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@13311.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@13313.4]
  assign SRAM_clock = clock; // @[:@13315.4]
  assign SRAM_reset = reset; // @[:@13316.4]
  assign SRAM_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@13358.4]
  assign SRAM_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_114; // @[MemPrimitives.scala 43:33:@13360.4]
  assign SRAM_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@13348.4]
  assign SRAM_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@13349.4]
  assign SRAM_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_110; // @[MemPrimitives.scala 37:29:@13355.4]
  assign SRAM_1_clock = clock; // @[:@13331.4]
  assign SRAM_1_reset = reset; // @[:@13332.4]
  assign SRAM_1_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@13374.4]
  assign SRAM_1_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_121; // @[MemPrimitives.scala 43:33:@13376.4]
  assign SRAM_1_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@13364.4]
  assign SRAM_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@13365.4]
  assign SRAM_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_117; // @[MemPrimitives.scala 37:29:@13371.4]
endmodule
module FF_12( // @[:@13550.2]
  input        clock, // @[:@13551.4]
  input        reset, // @[:@13552.4]
  output [3:0] io_rPort_0_output_0, // @[:@13553.4]
  input  [3:0] io_wPort_0_data_0, // @[:@13553.4]
  input        io_wPort_0_reset, // @[:@13553.4]
  input        io_wPort_0_en_0 // @[:@13553.4]
);
  reg [3:0] ff; // @[MemPrimitives.scala 321:19:@13568.4]
  reg [31:0] _RAND_0;
  wire [3:0] _T_68; // @[MemPrimitives.scala 325:32:@13570.4]
  wire [3:0] _T_69; // @[MemPrimitives.scala 325:12:@13571.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@13570.4]
  assign _T_69 = io_wPort_0_reset ? 4'h0 : _T_68; // @[MemPrimitives.scala 325:12:@13571.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@13573.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 4'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 4'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_6( // @[:@13588.2]
  input        clock, // @[:@13589.4]
  input        reset, // @[:@13590.4]
  input        io_setup_saturate, // @[:@13591.4]
  input        io_input_reset, // @[:@13591.4]
  input        io_input_enable, // @[:@13591.4]
  output [3:0] io_output_count_0, // @[:@13591.4]
  output       io_output_oobs_0, // @[:@13591.4]
  output       io_output_done // @[:@13591.4]
);
  wire  bases_0_clock; // @[Counter.scala 262:53:@13604.4]
  wire  bases_0_reset; // @[Counter.scala 262:53:@13604.4]
  wire [3:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 262:53:@13604.4]
  wire [3:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 262:53:@13604.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 262:53:@13604.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 262:53:@13604.4]
  wire  SRFF_clock; // @[Counter.scala 264:22:@13620.4]
  wire  SRFF_reset; // @[Counter.scala 264:22:@13620.4]
  wire  SRFF_io_input_set; // @[Counter.scala 264:22:@13620.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 264:22:@13620.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 264:22:@13620.4]
  wire  SRFF_io_output; // @[Counter.scala 264:22:@13620.4]
  wire  _T_36; // @[Counter.scala 265:45:@13623.4]
  wire [3:0] _T_48; // @[Counter.scala 288:52:@13648.4]
  wire [4:0] _T_50; // @[Counter.scala 292:33:@13649.4]
  wire [3:0] _T_51; // @[Counter.scala 292:33:@13650.4]
  wire [3:0] _T_52; // @[Counter.scala 292:33:@13651.4]
  wire  _T_57; // @[Counter.scala 294:18:@13653.4]
  wire [3:0] _T_68; // @[Counter.scala 300:115:@13661.4]
  wire [3:0] _T_70; // @[Counter.scala 300:85:@13663.4]
  wire [3:0] _T_71; // @[Counter.scala 300:152:@13664.4]
  wire [3:0] _T_72; // @[Counter.scala 300:74:@13665.4]
  wire  _T_75; // @[Counter.scala 323:102:@13669.4]
  wire  _T_77; // @[Counter.scala 323:130:@13670.4]
  FF_12 bases_0 ( // @[Counter.scala 262:53:@13604.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 264:22:@13620.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 265:45:@13623.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 288:52:@13648.4]
  assign _T_50 = $signed(_T_48) + $signed(4'sh1); // @[Counter.scala 292:33:@13649.4]
  assign _T_51 = $signed(_T_48) + $signed(4'sh1); // @[Counter.scala 292:33:@13650.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 292:33:@13651.4]
  assign _T_57 = $signed(_T_52) >= $signed(4'sh3); // @[Counter.scala 294:18:@13653.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 300:115:@13661.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 4'h0; // @[Counter.scala 300:85:@13663.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 300:152:@13664.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 300:74:@13665.4]
  assign _T_75 = $signed(_T_48) < $signed(4'sh0); // @[Counter.scala 323:102:@13669.4]
  assign _T_77 = $signed(_T_48) >= $signed(4'sh3); // @[Counter.scala 323:130:@13670.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 305:28:@13668.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 323:60:@13672.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 334:20:@13674.4]
  assign bases_0_clock = clock; // @[:@13605.4]
  assign bases_0_reset = reset; // @[:@13606.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 4'h0 : _T_72; // @[Counter.scala 300:31:@13667.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 282:27:@13646.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 285:29:@13647.4]
  assign SRFF_clock = clock; // @[:@13621.4]
  assign SRFF_reset = reset; // @[:@13622.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 265:23:@13625.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 266:25:@13627.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 267:30:@13628.4]
endmodule
module x549_ctrchain( // @[:@13679.2]
  input        clock, // @[:@13680.4]
  input        reset, // @[:@13681.4]
  input        io_input_reset, // @[:@13682.4]
  input        io_input_enable, // @[:@13682.4]
  output [3:0] io_output_counts_0, // @[:@13682.4]
  output       io_output_oobs_0, // @[:@13682.4]
  output       io_output_done // @[:@13682.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 514:46:@13684.4]
  wire  ctrs_0_reset; // @[Counter.scala 514:46:@13684.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 514:46:@13684.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 514:46:@13684.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 514:46:@13684.4]
  wire [3:0] ctrs_0_io_output_count_0; // @[Counter.scala 514:46:@13684.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 514:46:@13684.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 514:46:@13684.4]
  reg  wasDone; // @[Counter.scala 543:24:@13693.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 547:69:@13699.4]
  wire  _T_47; // @[Counter.scala 547:80:@13700.4]
  reg  doneLatch; // @[Counter.scala 551:26:@13705.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 552:48:@13706.4]
  wire  _T_55; // @[Counter.scala 552:19:@13707.4]
  SingleCounter_6 ctrs_0 ( // @[Counter.scala 514:46:@13684.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 547:69:@13699.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 547:80:@13700.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 552:48:@13706.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 552:19:@13707.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 558:32:@13709.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 559:30:@13711.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 547:18:@13702.4]
  assign ctrs_0_clock = clock; // @[:@13685.4]
  assign ctrs_0_reset = reset; // @[:@13686.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 531:29:@13692.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 521:24:@13690.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 525:33:@13691.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x653_outr_Reduce_sm( // @[:@14498.2]
  input   clock, // @[:@14499.4]
  input   reset, // @[:@14500.4]
  input   io_enable, // @[:@14501.4]
  output  io_done, // @[:@14501.4]
  input   io_ctrDone, // @[:@14501.4]
  output  io_ctrInc, // @[:@14501.4]
  output  io_ctrRst, // @[:@14501.4]
  input   io_parentAck, // @[:@14501.4]
  input   io_backpressure, // @[:@14501.4]
  input   io_doneIn_0, // @[:@14501.4]
  input   io_doneIn_1, // @[:@14501.4]
  input   io_doneIn_2, // @[:@14501.4]
  input   io_doneIn_3, // @[:@14501.4]
  input   io_doneIn_4, // @[:@14501.4]
  input   io_doneIn_5, // @[:@14501.4]
  input   io_doneIn_6, // @[:@14501.4]
  input   io_maskIn_0, // @[:@14501.4]
  input   io_maskIn_1, // @[:@14501.4]
  input   io_maskIn_2, // @[:@14501.4]
  input   io_maskIn_4, // @[:@14501.4]
  input   io_maskIn_5, // @[:@14501.4]
  output  io_enableOut_0, // @[:@14501.4]
  output  io_enableOut_1, // @[:@14501.4]
  output  io_enableOut_2, // @[:@14501.4]
  output  io_enableOut_3, // @[:@14501.4]
  output  io_enableOut_4, // @[:@14501.4]
  output  io_enableOut_5, // @[:@14501.4]
  output  io_enableOut_6, // @[:@14501.4]
  output  io_childAck_0, // @[:@14501.4]
  output  io_childAck_1, // @[:@14501.4]
  output  io_childAck_2, // @[:@14501.4]
  output  io_childAck_3, // @[:@14501.4]
  output  io_childAck_4, // @[:@14501.4]
  output  io_childAck_5, // @[:@14501.4]
  output  io_childAck_6 // @[:@14501.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@14504.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@14504.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@14504.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@14504.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@14504.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@14504.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@14507.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@14507.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@14507.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@14507.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@14507.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@14507.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@14510.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@14510.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@14510.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@14510.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@14510.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@14510.4]
  wire  active_3_clock; // @[Controllers.scala 76:50:@14513.4]
  wire  active_3_reset; // @[Controllers.scala 76:50:@14513.4]
  wire  active_3_io_input_set; // @[Controllers.scala 76:50:@14513.4]
  wire  active_3_io_input_reset; // @[Controllers.scala 76:50:@14513.4]
  wire  active_3_io_input_asyn_reset; // @[Controllers.scala 76:50:@14513.4]
  wire  active_3_io_output; // @[Controllers.scala 76:50:@14513.4]
  wire  active_4_clock; // @[Controllers.scala 76:50:@14516.4]
  wire  active_4_reset; // @[Controllers.scala 76:50:@14516.4]
  wire  active_4_io_input_set; // @[Controllers.scala 76:50:@14516.4]
  wire  active_4_io_input_reset; // @[Controllers.scala 76:50:@14516.4]
  wire  active_4_io_input_asyn_reset; // @[Controllers.scala 76:50:@14516.4]
  wire  active_4_io_output; // @[Controllers.scala 76:50:@14516.4]
  wire  active_5_clock; // @[Controllers.scala 76:50:@14519.4]
  wire  active_5_reset; // @[Controllers.scala 76:50:@14519.4]
  wire  active_5_io_input_set; // @[Controllers.scala 76:50:@14519.4]
  wire  active_5_io_input_reset; // @[Controllers.scala 76:50:@14519.4]
  wire  active_5_io_input_asyn_reset; // @[Controllers.scala 76:50:@14519.4]
  wire  active_5_io_output; // @[Controllers.scala 76:50:@14519.4]
  wire  active_6_clock; // @[Controllers.scala 76:50:@14522.4]
  wire  active_6_reset; // @[Controllers.scala 76:50:@14522.4]
  wire  active_6_io_input_set; // @[Controllers.scala 76:50:@14522.4]
  wire  active_6_io_input_reset; // @[Controllers.scala 76:50:@14522.4]
  wire  active_6_io_input_asyn_reset; // @[Controllers.scala 76:50:@14522.4]
  wire  active_6_io_output; // @[Controllers.scala 76:50:@14522.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@14525.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@14525.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@14525.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@14525.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@14525.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@14525.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@14528.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@14528.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@14528.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@14528.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@14528.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@14528.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@14531.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@14531.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@14531.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@14531.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@14531.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@14531.4]
  wire  done_3_clock; // @[Controllers.scala 77:48:@14534.4]
  wire  done_3_reset; // @[Controllers.scala 77:48:@14534.4]
  wire  done_3_io_input_set; // @[Controllers.scala 77:48:@14534.4]
  wire  done_3_io_input_reset; // @[Controllers.scala 77:48:@14534.4]
  wire  done_3_io_input_asyn_reset; // @[Controllers.scala 77:48:@14534.4]
  wire  done_3_io_output; // @[Controllers.scala 77:48:@14534.4]
  wire  done_4_clock; // @[Controllers.scala 77:48:@14537.4]
  wire  done_4_reset; // @[Controllers.scala 77:48:@14537.4]
  wire  done_4_io_input_set; // @[Controllers.scala 77:48:@14537.4]
  wire  done_4_io_input_reset; // @[Controllers.scala 77:48:@14537.4]
  wire  done_4_io_input_asyn_reset; // @[Controllers.scala 77:48:@14537.4]
  wire  done_4_io_output; // @[Controllers.scala 77:48:@14537.4]
  wire  done_5_clock; // @[Controllers.scala 77:48:@14540.4]
  wire  done_5_reset; // @[Controllers.scala 77:48:@14540.4]
  wire  done_5_io_input_set; // @[Controllers.scala 77:48:@14540.4]
  wire  done_5_io_input_reset; // @[Controllers.scala 77:48:@14540.4]
  wire  done_5_io_input_asyn_reset; // @[Controllers.scala 77:48:@14540.4]
  wire  done_5_io_output; // @[Controllers.scala 77:48:@14540.4]
  wire  done_6_clock; // @[Controllers.scala 77:48:@14543.4]
  wire  done_6_reset; // @[Controllers.scala 77:48:@14543.4]
  wire  done_6_io_input_set; // @[Controllers.scala 77:48:@14543.4]
  wire  done_6_io_input_reset; // @[Controllers.scala 77:48:@14543.4]
  wire  done_6_io_input_asyn_reset; // @[Controllers.scala 77:48:@14543.4]
  wire  done_6_io_output; // @[Controllers.scala 77:48:@14543.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@14632.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@14632.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@14632.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@14632.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@14632.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@14632.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@14635.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@14635.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@14635.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@14635.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@14635.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@14635.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@14638.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@14638.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@14638.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@14638.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@14638.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@14638.4]
  wire  iterDone_3_clock; // @[Controllers.scala 90:52:@14641.4]
  wire  iterDone_3_reset; // @[Controllers.scala 90:52:@14641.4]
  wire  iterDone_3_io_input_set; // @[Controllers.scala 90:52:@14641.4]
  wire  iterDone_3_io_input_reset; // @[Controllers.scala 90:52:@14641.4]
  wire  iterDone_3_io_input_asyn_reset; // @[Controllers.scala 90:52:@14641.4]
  wire  iterDone_3_io_output; // @[Controllers.scala 90:52:@14641.4]
  wire  iterDone_4_clock; // @[Controllers.scala 90:52:@14644.4]
  wire  iterDone_4_reset; // @[Controllers.scala 90:52:@14644.4]
  wire  iterDone_4_io_input_set; // @[Controllers.scala 90:52:@14644.4]
  wire  iterDone_4_io_input_reset; // @[Controllers.scala 90:52:@14644.4]
  wire  iterDone_4_io_input_asyn_reset; // @[Controllers.scala 90:52:@14644.4]
  wire  iterDone_4_io_output; // @[Controllers.scala 90:52:@14644.4]
  wire  iterDone_5_clock; // @[Controllers.scala 90:52:@14647.4]
  wire  iterDone_5_reset; // @[Controllers.scala 90:52:@14647.4]
  wire  iterDone_5_io_input_set; // @[Controllers.scala 90:52:@14647.4]
  wire  iterDone_5_io_input_reset; // @[Controllers.scala 90:52:@14647.4]
  wire  iterDone_5_io_input_asyn_reset; // @[Controllers.scala 90:52:@14647.4]
  wire  iterDone_5_io_output; // @[Controllers.scala 90:52:@14647.4]
  wire  iterDone_6_clock; // @[Controllers.scala 90:52:@14650.4]
  wire  iterDone_6_reset; // @[Controllers.scala 90:52:@14650.4]
  wire  iterDone_6_io_input_set; // @[Controllers.scala 90:52:@14650.4]
  wire  iterDone_6_io_input_reset; // @[Controllers.scala 90:52:@14650.4]
  wire  iterDone_6_io_input_asyn_reset; // @[Controllers.scala 90:52:@14650.4]
  wire  iterDone_6_io_output; // @[Controllers.scala 90:52:@14650.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@14746.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@14746.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@14746.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@14746.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@14746.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@14759.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@14759.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@14759.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@14759.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@14759.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@14772.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@14772.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@14772.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@14772.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@14772.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@14785.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@14785.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@14785.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@14785.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@14785.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@14798.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@14798.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@14798.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@14798.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@14798.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@14811.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@14811.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@14811.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@14811.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@14811.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@14842.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@14842.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@14842.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@14842.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@14842.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@14886.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@14886.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@14886.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@14886.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@14886.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@14910.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@14910.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@14910.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@14910.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@14910.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@14934.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@14934.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@14934.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@14934.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@14934.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@15081.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@15081.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@15081.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@15081.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@15081.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@15098.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@15098.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@15098.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@15098.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@15098.4]
  wire  _T_77; // @[Controllers.scala 80:47:@14546.4]
  wire  _T_78; // @[Controllers.scala 80:47:@14547.4]
  wire  _T_79; // @[Controllers.scala 80:47:@14548.4]
  wire  _T_80; // @[Controllers.scala 80:47:@14549.4]
  wire  _T_81; // @[Controllers.scala 80:47:@14550.4]
  wire  allDone; // @[Controllers.scala 80:47:@14551.4]
  wire  _T_253; // @[Controllers.scala 102:95:@14732.4]
  wire  _T_247; // @[Controllers.scala 101:55:@14726.4]
  wire  _T_248; // @[Controllers.scala 101:55:@14727.4]
  wire  _T_249; // @[Controllers.scala 101:55:@14728.4]
  wire  _T_250; // @[Controllers.scala 101:55:@14729.4]
  wire  _T_251; // @[Controllers.scala 101:55:@14730.4]
  wire  _T_252; // @[Controllers.scala 101:55:@14731.4]
  wire  _T_257; // @[package.scala 96:25:@14738.4 package.scala 96:25:@14739.4]
  wire  _T_260; // @[Controllers.scala 102:142:@14741.4]
  wire  _T_261; // @[Controllers.scala 102:138:@14742.4]
  wire  _T_262; // @[Controllers.scala 102:123:@14743.4]
  wire  _T_263; // @[Controllers.scala 102:112:@14744.4]
  wire  _T_264; // @[Controllers.scala 102:95:@14745.4]
  wire  _T_268; // @[package.scala 96:25:@14751.4 package.scala 96:25:@14752.4]
  wire  _T_271; // @[Controllers.scala 102:142:@14754.4]
  wire  _T_272; // @[Controllers.scala 102:138:@14755.4]
  wire  _T_273; // @[Controllers.scala 102:123:@14756.4]
  wire  _T_274; // @[Controllers.scala 102:112:@14757.4]
  wire  _T_330; // @[Controllers.scala 102:164:@14823.4]
  wire  _T_275; // @[Controllers.scala 102:95:@14758.4]
  wire  _T_279; // @[package.scala 96:25:@14764.4 package.scala 96:25:@14765.4]
  wire  _T_282; // @[Controllers.scala 102:142:@14767.4]
  wire  _T_283; // @[Controllers.scala 102:138:@14768.4]
  wire  _T_284; // @[Controllers.scala 102:123:@14769.4]
  wire  _T_285; // @[Controllers.scala 102:112:@14770.4]
  wire  _T_331; // @[Controllers.scala 102:164:@14824.4]
  wire  _T_286; // @[Controllers.scala 102:95:@14771.4]
  wire  _T_290; // @[package.scala 96:25:@14777.4 package.scala 96:25:@14778.4]
  wire  _T_293; // @[Controllers.scala 102:142:@14780.4]
  wire  _T_294; // @[Controllers.scala 102:138:@14781.4]
  wire  _T_295; // @[Controllers.scala 102:123:@14782.4]
  wire  _T_296; // @[Controllers.scala 102:112:@14783.4]
  wire  _T_332; // @[Controllers.scala 102:164:@14825.4]
  wire  _T_297; // @[Controllers.scala 102:95:@14784.4]
  wire  _T_301; // @[package.scala 96:25:@14790.4 package.scala 96:25:@14791.4]
  wire  _T_304; // @[Controllers.scala 102:142:@14793.4]
  wire  _T_305; // @[Controllers.scala 102:138:@14794.4]
  wire  _T_306; // @[Controllers.scala 102:123:@14795.4]
  wire  _T_307; // @[Controllers.scala 102:112:@14796.4]
  wire  _T_333; // @[Controllers.scala 102:164:@14826.4]
  wire  _T_308; // @[Controllers.scala 102:95:@14797.4]
  wire  _T_312; // @[package.scala 96:25:@14803.4 package.scala 96:25:@14804.4]
  wire  _T_315; // @[Controllers.scala 102:142:@14806.4]
  wire  _T_316; // @[Controllers.scala 102:138:@14807.4]
  wire  _T_317; // @[Controllers.scala 102:123:@14808.4]
  wire  _T_318; // @[Controllers.scala 102:112:@14809.4]
  wire  _T_334; // @[Controllers.scala 102:164:@14827.4]
  wire  _T_319; // @[Controllers.scala 102:95:@14810.4]
  wire  _T_323; // @[package.scala 96:25:@14816.4 package.scala 96:25:@14817.4]
  wire  _T_326; // @[Controllers.scala 102:142:@14819.4]
  wire  _T_327; // @[Controllers.scala 102:138:@14820.4]
  wire  _T_328; // @[Controllers.scala 102:123:@14821.4]
  wire  _T_329; // @[Controllers.scala 102:112:@14822.4]
  wire  synchronize; // @[Controllers.scala 102:164:@14828.4]
  wire  _T_337; // @[Controllers.scala 105:33:@14830.4]
  wire  _T_339; // @[Controllers.scala 105:54:@14831.4]
  wire  _T_340; // @[Controllers.scala 105:52:@14832.4]
  wire  _T_346; // @[Controllers.scala 107:51:@14839.4]
  wire  _T_349; // @[Controllers.scala 107:64:@14841.4]
  wire  _T_353; // @[package.scala 96:25:@14847.4 package.scala 96:25:@14848.4]
  wire  _T_357; // @[Controllers.scala 107:89:@14850.4]
  wire  _T_358; // @[Controllers.scala 107:86:@14851.4]
  wire  _T_359; // @[Controllers.scala 107:108:@14852.4]
  wire  _T_374; // @[Controllers.scala 114:49:@14870.4]
  wire  _T_377; // @[Controllers.scala 115:57:@14874.4]
  wire  _T_393; // @[Controllers.scala 114:49:@14894.4]
  wire  _T_396; // @[Controllers.scala 115:57:@14898.4]
  wire  _T_412; // @[Controllers.scala 114:49:@14918.4]
  wire  _T_415; // @[Controllers.scala 115:57:@14922.4]
  wire  _T_431; // @[Controllers.scala 114:49:@14942.4]
  wire  _T_434; // @[Controllers.scala 115:57:@14946.4]
  wire  _T_450; // @[Controllers.scala 114:49:@14966.4]
  wire  _T_453; // @[Controllers.scala 115:57:@14970.4]
  wire  _T_469; // @[Controllers.scala 114:49:@14990.4]
  wire  _T_472; // @[Controllers.scala 115:57:@14994.4]
  wire  _T_488; // @[Controllers.scala 213:68:@15019.4]
  wire  _T_489; // @[Controllers.scala 213:92:@15020.4]
  wire  _T_490; // @[Controllers.scala 213:90:@15021.4]
  wire  _T_491; // @[Controllers.scala 213:115:@15022.4]
  wire  _T_492; // @[Controllers.scala 213:132:@15023.4]
  wire  _T_493; // @[Controllers.scala 213:130:@15024.4]
  wire  _T_494; // @[Controllers.scala 213:156:@15025.4]
  wire  _T_496; // @[Controllers.scala 213:68:@15028.4]
  wire  _T_497; // @[Controllers.scala 213:92:@15029.4]
  wire  _T_498; // @[Controllers.scala 213:90:@15030.4]
  wire  _T_499; // @[Controllers.scala 213:115:@15031.4]
  wire  _T_504; // @[Controllers.scala 213:68:@15036.4]
  wire  _T_505; // @[Controllers.scala 213:92:@15037.4]
  wire  _T_506; // @[Controllers.scala 213:90:@15038.4]
  wire  _T_507; // @[Controllers.scala 213:115:@15039.4]
  wire  _T_512; // @[Controllers.scala 213:68:@15044.4]
  wire  _T_513; // @[Controllers.scala 213:92:@15045.4]
  wire  _T_514; // @[Controllers.scala 213:90:@15046.4]
  wire  _T_520; // @[Controllers.scala 213:68:@15052.4]
  wire  _T_521; // @[Controllers.scala 213:92:@15053.4]
  wire  _T_522; // @[Controllers.scala 213:90:@15054.4]
  wire  _T_523; // @[Controllers.scala 213:115:@15055.4]
  wire  _T_528; // @[Controllers.scala 213:68:@15060.4]
  wire  _T_529; // @[Controllers.scala 213:92:@15061.4]
  wire  _T_530; // @[Controllers.scala 213:90:@15062.4]
  wire  _T_531; // @[Controllers.scala 213:115:@15063.4]
  wire  _T_536; // @[Controllers.scala 213:68:@15068.4]
  wire  _T_537; // @[Controllers.scala 213:92:@15069.4]
  wire  _T_538; // @[Controllers.scala 213:90:@15070.4]
  wire  _T_545; // @[package.scala 100:49:@15076.4]
  reg  _T_548; // @[package.scala 48:56:@15077.4]
  reg [31:0] _RAND_0;
  wire  _T_549; // @[package.scala 100:41:@15079.4]
  reg  _T_562; // @[package.scala 48:56:@15095.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@14504.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@14507.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@14510.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF active_3 ( // @[Controllers.scala 76:50:@14513.4]
    .clock(active_3_clock),
    .reset(active_3_reset),
    .io_input_set(active_3_io_input_set),
    .io_input_reset(active_3_io_input_reset),
    .io_input_asyn_reset(active_3_io_input_asyn_reset),
    .io_output(active_3_io_output)
  );
  SRFF active_4 ( // @[Controllers.scala 76:50:@14516.4]
    .clock(active_4_clock),
    .reset(active_4_reset),
    .io_input_set(active_4_io_input_set),
    .io_input_reset(active_4_io_input_reset),
    .io_input_asyn_reset(active_4_io_input_asyn_reset),
    .io_output(active_4_io_output)
  );
  SRFF active_5 ( // @[Controllers.scala 76:50:@14519.4]
    .clock(active_5_clock),
    .reset(active_5_reset),
    .io_input_set(active_5_io_input_set),
    .io_input_reset(active_5_io_input_reset),
    .io_input_asyn_reset(active_5_io_input_asyn_reset),
    .io_output(active_5_io_output)
  );
  SRFF active_6 ( // @[Controllers.scala 76:50:@14522.4]
    .clock(active_6_clock),
    .reset(active_6_reset),
    .io_input_set(active_6_io_input_set),
    .io_input_reset(active_6_io_input_reset),
    .io_input_asyn_reset(active_6_io_input_asyn_reset),
    .io_output(active_6_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@14525.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@14528.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@14531.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF done_3 ( // @[Controllers.scala 77:48:@14534.4]
    .clock(done_3_clock),
    .reset(done_3_reset),
    .io_input_set(done_3_io_input_set),
    .io_input_reset(done_3_io_input_reset),
    .io_input_asyn_reset(done_3_io_input_asyn_reset),
    .io_output(done_3_io_output)
  );
  SRFF done_4 ( // @[Controllers.scala 77:48:@14537.4]
    .clock(done_4_clock),
    .reset(done_4_reset),
    .io_input_set(done_4_io_input_set),
    .io_input_reset(done_4_io_input_reset),
    .io_input_asyn_reset(done_4_io_input_asyn_reset),
    .io_output(done_4_io_output)
  );
  SRFF done_5 ( // @[Controllers.scala 77:48:@14540.4]
    .clock(done_5_clock),
    .reset(done_5_reset),
    .io_input_set(done_5_io_input_set),
    .io_input_reset(done_5_io_input_reset),
    .io_input_asyn_reset(done_5_io_input_asyn_reset),
    .io_output(done_5_io_output)
  );
  SRFF done_6 ( // @[Controllers.scala 77:48:@14543.4]
    .clock(done_6_clock),
    .reset(done_6_reset),
    .io_input_set(done_6_io_input_set),
    .io_input_reset(done_6_io_input_reset),
    .io_input_asyn_reset(done_6_io_input_asyn_reset),
    .io_output(done_6_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@14632.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@14635.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@14638.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  SRFF iterDone_3 ( // @[Controllers.scala 90:52:@14641.4]
    .clock(iterDone_3_clock),
    .reset(iterDone_3_reset),
    .io_input_set(iterDone_3_io_input_set),
    .io_input_reset(iterDone_3_io_input_reset),
    .io_input_asyn_reset(iterDone_3_io_input_asyn_reset),
    .io_output(iterDone_3_io_output)
  );
  SRFF iterDone_4 ( // @[Controllers.scala 90:52:@14644.4]
    .clock(iterDone_4_clock),
    .reset(iterDone_4_reset),
    .io_input_set(iterDone_4_io_input_set),
    .io_input_reset(iterDone_4_io_input_reset),
    .io_input_asyn_reset(iterDone_4_io_input_asyn_reset),
    .io_output(iterDone_4_io_output)
  );
  SRFF iterDone_5 ( // @[Controllers.scala 90:52:@14647.4]
    .clock(iterDone_5_clock),
    .reset(iterDone_5_reset),
    .io_input_set(iterDone_5_io_input_set),
    .io_input_reset(iterDone_5_io_input_reset),
    .io_input_asyn_reset(iterDone_5_io_input_asyn_reset),
    .io_output(iterDone_5_io_output)
  );
  SRFF iterDone_6 ( // @[Controllers.scala 90:52:@14650.4]
    .clock(iterDone_6_clock),
    .reset(iterDone_6_reset),
    .io_input_set(iterDone_6_io_input_set),
    .io_input_reset(iterDone_6_io_input_reset),
    .io_input_asyn_reset(iterDone_6_io_input_asyn_reset),
    .io_output(iterDone_6_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@14733.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@14746.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@14759.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@14772.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@14785.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@14798.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@14811.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@14842.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@14862.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@14886.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@14910.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 ( // @[package.scala 93:22:@14934.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper RetimeWrapper_12 ( // @[package.scala 93:22:@14958.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 ( // @[package.scala 93:22:@14982.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@15081.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@15098.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@14546.4]
  assign _T_78 = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@14547.4]
  assign _T_79 = _T_78 & done_3_io_output; // @[Controllers.scala 80:47:@14548.4]
  assign _T_80 = _T_79 & done_4_io_output; // @[Controllers.scala 80:47:@14549.4]
  assign _T_81 = _T_80 & done_5_io_output; // @[Controllers.scala 80:47:@14550.4]
  assign allDone = _T_81 & done_6_io_output; // @[Controllers.scala 80:47:@14551.4]
  assign _T_253 = active_0_io_output == iterDone_0_io_output; // @[Controllers.scala 102:95:@14732.4]
  assign _T_247 = iterDone_0_io_output | iterDone_1_io_output; // @[Controllers.scala 101:55:@14726.4]
  assign _T_248 = _T_247 | iterDone_2_io_output; // @[Controllers.scala 101:55:@14727.4]
  assign _T_249 = _T_248 | iterDone_3_io_output; // @[Controllers.scala 101:55:@14728.4]
  assign _T_250 = _T_249 | iterDone_4_io_output; // @[Controllers.scala 101:55:@14729.4]
  assign _T_251 = _T_250 | iterDone_5_io_output; // @[Controllers.scala 101:55:@14730.4]
  assign _T_252 = _T_251 | iterDone_6_io_output; // @[Controllers.scala 101:55:@14731.4]
  assign _T_257 = RetimeWrapper_io_out; // @[package.scala 96:25:@14738.4 package.scala 96:25:@14739.4]
  assign _T_260 = ~ _T_257; // @[Controllers.scala 102:142:@14741.4]
  assign _T_261 = active_0_io_output == _T_260; // @[Controllers.scala 102:138:@14742.4]
  assign _T_262 = _T_252 & _T_261; // @[Controllers.scala 102:123:@14743.4]
  assign _T_263 = _T_253 | _T_262; // @[Controllers.scala 102:112:@14744.4]
  assign _T_264 = active_1_io_output == iterDone_1_io_output; // @[Controllers.scala 102:95:@14745.4]
  assign _T_268 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@14751.4 package.scala 96:25:@14752.4]
  assign _T_271 = ~ _T_268; // @[Controllers.scala 102:142:@14754.4]
  assign _T_272 = active_1_io_output == _T_271; // @[Controllers.scala 102:138:@14755.4]
  assign _T_273 = _T_252 & _T_272; // @[Controllers.scala 102:123:@14756.4]
  assign _T_274 = _T_264 | _T_273; // @[Controllers.scala 102:112:@14757.4]
  assign _T_330 = _T_263 & _T_274; // @[Controllers.scala 102:164:@14823.4]
  assign _T_275 = active_2_io_output == iterDone_2_io_output; // @[Controllers.scala 102:95:@14758.4]
  assign _T_279 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@14764.4 package.scala 96:25:@14765.4]
  assign _T_282 = ~ _T_279; // @[Controllers.scala 102:142:@14767.4]
  assign _T_283 = active_2_io_output == _T_282; // @[Controllers.scala 102:138:@14768.4]
  assign _T_284 = _T_252 & _T_283; // @[Controllers.scala 102:123:@14769.4]
  assign _T_285 = _T_275 | _T_284; // @[Controllers.scala 102:112:@14770.4]
  assign _T_331 = _T_330 & _T_285; // @[Controllers.scala 102:164:@14824.4]
  assign _T_286 = active_3_io_output == iterDone_3_io_output; // @[Controllers.scala 102:95:@14771.4]
  assign _T_290 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@14777.4 package.scala 96:25:@14778.4]
  assign _T_293 = ~ _T_290; // @[Controllers.scala 102:142:@14780.4]
  assign _T_294 = active_3_io_output == _T_293; // @[Controllers.scala 102:138:@14781.4]
  assign _T_295 = _T_252 & _T_294; // @[Controllers.scala 102:123:@14782.4]
  assign _T_296 = _T_286 | _T_295; // @[Controllers.scala 102:112:@14783.4]
  assign _T_332 = _T_331 & _T_296; // @[Controllers.scala 102:164:@14825.4]
  assign _T_297 = active_4_io_output == iterDone_4_io_output; // @[Controllers.scala 102:95:@14784.4]
  assign _T_301 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@14790.4 package.scala 96:25:@14791.4]
  assign _T_304 = ~ _T_301; // @[Controllers.scala 102:142:@14793.4]
  assign _T_305 = active_4_io_output == _T_304; // @[Controllers.scala 102:138:@14794.4]
  assign _T_306 = _T_252 & _T_305; // @[Controllers.scala 102:123:@14795.4]
  assign _T_307 = _T_297 | _T_306; // @[Controllers.scala 102:112:@14796.4]
  assign _T_333 = _T_332 & _T_307; // @[Controllers.scala 102:164:@14826.4]
  assign _T_308 = active_5_io_output == iterDone_5_io_output; // @[Controllers.scala 102:95:@14797.4]
  assign _T_312 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@14803.4 package.scala 96:25:@14804.4]
  assign _T_315 = ~ _T_312; // @[Controllers.scala 102:142:@14806.4]
  assign _T_316 = active_5_io_output == _T_315; // @[Controllers.scala 102:138:@14807.4]
  assign _T_317 = _T_252 & _T_316; // @[Controllers.scala 102:123:@14808.4]
  assign _T_318 = _T_308 | _T_317; // @[Controllers.scala 102:112:@14809.4]
  assign _T_334 = _T_333 & _T_318; // @[Controllers.scala 102:164:@14827.4]
  assign _T_319 = active_6_io_output == iterDone_6_io_output; // @[Controllers.scala 102:95:@14810.4]
  assign _T_323 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@14816.4 package.scala 96:25:@14817.4]
  assign _T_326 = ~ _T_323; // @[Controllers.scala 102:142:@14819.4]
  assign _T_327 = active_6_io_output == _T_326; // @[Controllers.scala 102:138:@14820.4]
  assign _T_328 = _T_252 & _T_327; // @[Controllers.scala 102:123:@14821.4]
  assign _T_329 = _T_319 | _T_328; // @[Controllers.scala 102:112:@14822.4]
  assign synchronize = _T_334 & _T_329; // @[Controllers.scala 102:164:@14828.4]
  assign _T_337 = done_0_io_output == 1'h0; // @[Controllers.scala 105:33:@14830.4]
  assign _T_339 = io_ctrDone == 1'h0; // @[Controllers.scala 105:54:@14831.4]
  assign _T_340 = _T_337 & _T_339; // @[Controllers.scala 105:52:@14832.4]
  assign _T_346 = synchronize == 1'h0; // @[Controllers.scala 107:51:@14839.4]
  assign _T_349 = _T_346 & _T_337; // @[Controllers.scala 107:64:@14841.4]
  assign _T_353 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@14847.4 package.scala 96:25:@14848.4]
  assign _T_357 = _T_353 == 1'h0; // @[Controllers.scala 107:89:@14850.4]
  assign _T_358 = _T_349 & _T_357; // @[Controllers.scala 107:86:@14851.4]
  assign _T_359 = _T_358 & io_enable; // @[Controllers.scala 107:108:@14852.4]
  assign _T_374 = synchronize & active_0_io_output; // @[Controllers.scala 114:49:@14870.4]
  assign _T_377 = done_0_io_output & synchronize; // @[Controllers.scala 115:57:@14874.4]
  assign _T_393 = synchronize & active_1_io_output; // @[Controllers.scala 114:49:@14894.4]
  assign _T_396 = done_1_io_output & synchronize; // @[Controllers.scala 115:57:@14898.4]
  assign _T_412 = synchronize & active_2_io_output; // @[Controllers.scala 114:49:@14918.4]
  assign _T_415 = done_2_io_output & synchronize; // @[Controllers.scala 115:57:@14922.4]
  assign _T_431 = synchronize & active_3_io_output; // @[Controllers.scala 114:49:@14942.4]
  assign _T_434 = done_3_io_output & synchronize; // @[Controllers.scala 115:57:@14946.4]
  assign _T_450 = synchronize & active_4_io_output; // @[Controllers.scala 114:49:@14966.4]
  assign _T_453 = done_4_io_output & synchronize; // @[Controllers.scala 115:57:@14970.4]
  assign _T_469 = synchronize & active_5_io_output; // @[Controllers.scala 114:49:@14990.4]
  assign _T_472 = done_5_io_output & synchronize; // @[Controllers.scala 115:57:@14994.4]
  assign _T_488 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@15019.4]
  assign _T_489 = ~ iterDone_0_io_output; // @[Controllers.scala 213:92:@15020.4]
  assign _T_490 = _T_488 & _T_489; // @[Controllers.scala 213:90:@15021.4]
  assign _T_491 = _T_490 & io_maskIn_0; // @[Controllers.scala 213:115:@15022.4]
  assign _T_492 = ~ allDone; // @[Controllers.scala 213:132:@15023.4]
  assign _T_493 = _T_491 & _T_492; // @[Controllers.scala 213:130:@15024.4]
  assign _T_494 = ~ io_ctrDone; // @[Controllers.scala 213:156:@15025.4]
  assign _T_496 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@15028.4]
  assign _T_497 = ~ iterDone_1_io_output; // @[Controllers.scala 213:92:@15029.4]
  assign _T_498 = _T_496 & _T_497; // @[Controllers.scala 213:90:@15030.4]
  assign _T_499 = _T_498 & io_maskIn_1; // @[Controllers.scala 213:115:@15031.4]
  assign _T_504 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@15036.4]
  assign _T_505 = ~ iterDone_2_io_output; // @[Controllers.scala 213:92:@15037.4]
  assign _T_506 = _T_504 & _T_505; // @[Controllers.scala 213:90:@15038.4]
  assign _T_507 = _T_506 & io_maskIn_2; // @[Controllers.scala 213:115:@15039.4]
  assign _T_512 = io_enable & active_3_io_output; // @[Controllers.scala 213:68:@15044.4]
  assign _T_513 = ~ iterDone_3_io_output; // @[Controllers.scala 213:92:@15045.4]
  assign _T_514 = _T_512 & _T_513; // @[Controllers.scala 213:90:@15046.4]
  assign _T_520 = io_enable & active_4_io_output; // @[Controllers.scala 213:68:@15052.4]
  assign _T_521 = ~ iterDone_4_io_output; // @[Controllers.scala 213:92:@15053.4]
  assign _T_522 = _T_520 & _T_521; // @[Controllers.scala 213:90:@15054.4]
  assign _T_523 = _T_522 & io_maskIn_4; // @[Controllers.scala 213:115:@15055.4]
  assign _T_528 = io_enable & active_5_io_output; // @[Controllers.scala 213:68:@15060.4]
  assign _T_529 = ~ iterDone_5_io_output; // @[Controllers.scala 213:92:@15061.4]
  assign _T_530 = _T_528 & _T_529; // @[Controllers.scala 213:90:@15062.4]
  assign _T_531 = _T_530 & io_maskIn_5; // @[Controllers.scala 213:115:@15063.4]
  assign _T_536 = io_enable & active_6_io_output; // @[Controllers.scala 213:68:@15068.4]
  assign _T_537 = ~ iterDone_6_io_output; // @[Controllers.scala 213:92:@15069.4]
  assign _T_538 = _T_536 & _T_537; // @[Controllers.scala 213:90:@15070.4]
  assign _T_545 = allDone == 1'h0; // @[package.scala 100:49:@15076.4]
  assign _T_549 = allDone & _T_548; // @[package.scala 100:41:@15079.4]
  assign io_done = RetimeWrapper_15_io_out; // @[Controllers.scala 245:13:@15105.4]
  assign io_ctrInc = iterDone_0_io_output & synchronize; // @[Controllers.scala 98:17:@14725.4]
  assign io_ctrRst = RetimeWrapper_14_io_out; // @[Controllers.scala 215:13:@15088.4]
  assign io_enableOut_0 = _T_493 & _T_494; // @[Controllers.scala 213:55:@15027.4]
  assign io_enableOut_1 = _T_499 & _T_492; // @[Controllers.scala 213:55:@15035.4]
  assign io_enableOut_2 = _T_507 & _T_492; // @[Controllers.scala 213:55:@15043.4]
  assign io_enableOut_3 = _T_514 & _T_492; // @[Controllers.scala 213:55:@15051.4]
  assign io_enableOut_4 = _T_523 & _T_492; // @[Controllers.scala 213:55:@15059.4]
  assign io_enableOut_5 = _T_531 & _T_492; // @[Controllers.scala 213:55:@15067.4]
  assign io_enableOut_6 = _T_538 & _T_492; // @[Controllers.scala 213:55:@15075.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@15006.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@15008.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@15010.4]
  assign io_childAck_3 = iterDone_3_io_output; // @[Controllers.scala 212:58:@15012.4]
  assign io_childAck_4 = iterDone_4_io_output; // @[Controllers.scala 212:58:@15014.4]
  assign io_childAck_5 = iterDone_5_io_output; // @[Controllers.scala 212:58:@15016.4]
  assign io_childAck_6 = iterDone_6_io_output; // @[Controllers.scala 212:58:@15018.4]
  assign active_0_clock = clock; // @[:@14505.4]
  assign active_0_reset = reset; // @[:@14506.4]
  assign active_0_io_input_set = _T_340 & io_enable; // @[Controllers.scala 105:30:@14835.4]
  assign active_0_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 106:32:@14838.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@14554.4]
  assign active_1_clock = clock; // @[:@14508.4]
  assign active_1_reset = reset; // @[:@14509.4]
  assign active_1_io_input_set = _T_374 & io_enable; // @[Controllers.scala 114:32:@14873.4]
  assign active_1_io_input_reset = _T_377 | io_parentAck; // @[Controllers.scala 115:34:@14877.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@14555.4]
  assign active_2_clock = clock; // @[:@14511.4]
  assign active_2_reset = reset; // @[:@14512.4]
  assign active_2_io_input_set = _T_393 & io_enable; // @[Controllers.scala 114:32:@14897.4]
  assign active_2_io_input_reset = _T_396 | io_parentAck; // @[Controllers.scala 115:34:@14901.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@14556.4]
  assign active_3_clock = clock; // @[:@14514.4]
  assign active_3_reset = reset; // @[:@14515.4]
  assign active_3_io_input_set = _T_412 & io_enable; // @[Controllers.scala 114:32:@14921.4]
  assign active_3_io_input_reset = _T_415 | io_parentAck; // @[Controllers.scala 115:34:@14925.4]
  assign active_3_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@14557.4]
  assign active_4_clock = clock; // @[:@14517.4]
  assign active_4_reset = reset; // @[:@14518.4]
  assign active_4_io_input_set = _T_431 & io_enable; // @[Controllers.scala 114:32:@14945.4]
  assign active_4_io_input_reset = _T_434 | io_parentAck; // @[Controllers.scala 115:34:@14949.4]
  assign active_4_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@14558.4]
  assign active_5_clock = clock; // @[:@14520.4]
  assign active_5_reset = reset; // @[:@14521.4]
  assign active_5_io_input_set = _T_450 & io_enable; // @[Controllers.scala 114:32:@14969.4]
  assign active_5_io_input_reset = _T_453 | io_parentAck; // @[Controllers.scala 115:34:@14973.4]
  assign active_5_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@14559.4]
  assign active_6_clock = clock; // @[:@14523.4]
  assign active_6_reset = reset; // @[:@14524.4]
  assign active_6_io_input_set = _T_469 & io_enable; // @[Controllers.scala 114:32:@14993.4]
  assign active_6_io_input_reset = _T_472 | io_parentAck; // @[Controllers.scala 115:34:@14997.4]
  assign active_6_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@14560.4]
  assign done_0_clock = clock; // @[:@14526.4]
  assign done_0_reset = reset; // @[:@14527.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 108:28:@14860.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@14576.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@14561.4]
  assign done_1_clock = clock; // @[:@14529.4]
  assign done_1_reset = reset; // @[:@14530.4]
  assign done_1_io_input_set = done_0_io_output & synchronize; // @[Controllers.scala 117:30:@14884.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@14585.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@14562.4]
  assign done_2_clock = clock; // @[:@14532.4]
  assign done_2_reset = reset; // @[:@14533.4]
  assign done_2_io_input_set = done_1_io_output & synchronize; // @[Controllers.scala 117:30:@14908.4]
  assign done_2_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@14594.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@14563.4]
  assign done_3_clock = clock; // @[:@14535.4]
  assign done_3_reset = reset; // @[:@14536.4]
  assign done_3_io_input_set = done_2_io_output & synchronize; // @[Controllers.scala 117:30:@14932.4]
  assign done_3_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@14603.4]
  assign done_3_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@14564.4]
  assign done_4_clock = clock; // @[:@14538.4]
  assign done_4_reset = reset; // @[:@14539.4]
  assign done_4_io_input_set = done_3_io_output & synchronize; // @[Controllers.scala 117:30:@14956.4]
  assign done_4_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@14612.4]
  assign done_4_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@14565.4]
  assign done_5_clock = clock; // @[:@14541.4]
  assign done_5_reset = reset; // @[:@14542.4]
  assign done_5_io_input_set = done_4_io_output & synchronize; // @[Controllers.scala 117:30:@14980.4]
  assign done_5_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@14621.4]
  assign done_5_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@14566.4]
  assign done_6_clock = clock; // @[:@14544.4]
  assign done_6_reset = reset; // @[:@14545.4]
  assign done_6_io_input_set = done_5_io_output & synchronize; // @[Controllers.scala 117:30:@15004.4]
  assign done_6_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@14630.4]
  assign done_6_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@14567.4]
  assign iterDone_0_clock = clock; // @[:@14633.4]
  assign iterDone_0_reset = reset; // @[:@14634.4]
  assign iterDone_0_io_input_set = io_doneIn_0 | _T_359; // @[Controllers.scala 107:32:@14856.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@14668.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@14653.4]
  assign iterDone_1_clock = clock; // @[:@14636.4]
  assign iterDone_1_reset = reset; // @[:@14637.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 116:34:@14879.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@14677.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@14654.4]
  assign iterDone_2_clock = clock; // @[:@14639.4]
  assign iterDone_2_reset = reset; // @[:@14640.4]
  assign iterDone_2_io_input_set = io_doneIn_2; // @[Controllers.scala 116:34:@14903.4]
  assign iterDone_2_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@14686.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@14655.4]
  assign iterDone_3_clock = clock; // @[:@14642.4]
  assign iterDone_3_reset = reset; // @[:@14643.4]
  assign iterDone_3_io_input_set = io_doneIn_3; // @[Controllers.scala 116:34:@14927.4]
  assign iterDone_3_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@14695.4]
  assign iterDone_3_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@14656.4]
  assign iterDone_4_clock = clock; // @[:@14645.4]
  assign iterDone_4_reset = reset; // @[:@14646.4]
  assign iterDone_4_io_input_set = io_doneIn_4; // @[Controllers.scala 116:34:@14951.4]
  assign iterDone_4_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@14704.4]
  assign iterDone_4_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@14657.4]
  assign iterDone_5_clock = clock; // @[:@14648.4]
  assign iterDone_5_reset = reset; // @[:@14649.4]
  assign iterDone_5_io_input_set = io_doneIn_5; // @[Controllers.scala 116:34:@14975.4]
  assign iterDone_5_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@14713.4]
  assign iterDone_5_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@14658.4]
  assign iterDone_6_clock = clock; // @[:@14651.4]
  assign iterDone_6_reset = reset; // @[:@14652.4]
  assign iterDone_6_io_input_set = io_doneIn_6; // @[Controllers.scala 116:34:@14999.4]
  assign iterDone_6_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@14722.4]
  assign iterDone_6_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@14659.4]
  assign RetimeWrapper_clock = clock; // @[:@14734.4]
  assign RetimeWrapper_reset = reset; // @[:@14735.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@14737.4]
  assign RetimeWrapper_io_in = io_maskIn_0; // @[package.scala 94:16:@14736.4]
  assign RetimeWrapper_1_clock = clock; // @[:@14747.4]
  assign RetimeWrapper_1_reset = reset; // @[:@14748.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@14750.4]
  assign RetimeWrapper_1_io_in = io_maskIn_1; // @[package.scala 94:16:@14749.4]
  assign RetimeWrapper_2_clock = clock; // @[:@14760.4]
  assign RetimeWrapper_2_reset = reset; // @[:@14761.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@14763.4]
  assign RetimeWrapper_2_io_in = io_maskIn_2; // @[package.scala 94:16:@14762.4]
  assign RetimeWrapper_3_clock = clock; // @[:@14773.4]
  assign RetimeWrapper_3_reset = reset; // @[:@14774.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@14776.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@14775.4]
  assign RetimeWrapper_4_clock = clock; // @[:@14786.4]
  assign RetimeWrapper_4_reset = reset; // @[:@14787.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@14789.4]
  assign RetimeWrapper_4_io_in = io_maskIn_4; // @[package.scala 94:16:@14788.4]
  assign RetimeWrapper_5_clock = clock; // @[:@14799.4]
  assign RetimeWrapper_5_reset = reset; // @[:@14800.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@14802.4]
  assign RetimeWrapper_5_io_in = io_maskIn_5; // @[package.scala 94:16:@14801.4]
  assign RetimeWrapper_6_clock = clock; // @[:@14812.4]
  assign RetimeWrapper_6_reset = reset; // @[:@14813.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@14815.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@14814.4]
  assign RetimeWrapper_7_clock = clock; // @[:@14843.4]
  assign RetimeWrapper_7_reset = reset; // @[:@14844.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@14846.4]
  assign RetimeWrapper_7_io_in = io_maskIn_0; // @[package.scala 94:16:@14845.4]
  assign RetimeWrapper_8_clock = clock; // @[:@14863.4]
  assign RetimeWrapper_8_reset = reset; // @[:@14864.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@14866.4]
  assign RetimeWrapper_8_io_in = synchronize & iterDone_0_io_output; // @[package.scala 94:16:@14865.4]
  assign RetimeWrapper_9_clock = clock; // @[:@14887.4]
  assign RetimeWrapper_9_reset = reset; // @[:@14888.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@14890.4]
  assign RetimeWrapper_9_io_in = synchronize & iterDone_1_io_output; // @[package.scala 94:16:@14889.4]
  assign RetimeWrapper_10_clock = clock; // @[:@14911.4]
  assign RetimeWrapper_10_reset = reset; // @[:@14912.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@14914.4]
  assign RetimeWrapper_10_io_in = synchronize & iterDone_2_io_output; // @[package.scala 94:16:@14913.4]
  assign RetimeWrapper_11_clock = clock; // @[:@14935.4]
  assign RetimeWrapper_11_reset = reset; // @[:@14936.4]
  assign RetimeWrapper_11_io_flow = 1'h1; // @[package.scala 95:18:@14938.4]
  assign RetimeWrapper_11_io_in = synchronize & iterDone_3_io_output; // @[package.scala 94:16:@14937.4]
  assign RetimeWrapper_12_clock = clock; // @[:@14959.4]
  assign RetimeWrapper_12_reset = reset; // @[:@14960.4]
  assign RetimeWrapper_12_io_flow = 1'h1; // @[package.scala 95:18:@14962.4]
  assign RetimeWrapper_12_io_in = synchronize & iterDone_4_io_output; // @[package.scala 94:16:@14961.4]
  assign RetimeWrapper_13_clock = clock; // @[:@14983.4]
  assign RetimeWrapper_13_reset = reset; // @[:@14984.4]
  assign RetimeWrapper_13_io_flow = 1'h1; // @[package.scala 95:18:@14986.4]
  assign RetimeWrapper_13_io_in = synchronize & iterDone_5_io_output; // @[package.scala 94:16:@14985.4]
  assign RetimeWrapper_14_clock = clock; // @[:@15082.4]
  assign RetimeWrapper_14_reset = reset; // @[:@15083.4]
  assign RetimeWrapper_14_io_flow = 1'h1; // @[package.scala 95:18:@15085.4]
  assign RetimeWrapper_14_io_in = _T_549 | io_parentAck; // @[package.scala 94:16:@15084.4]
  assign RetimeWrapper_15_clock = clock; // @[:@15099.4]
  assign RetimeWrapper_15_reset = reset; // @[:@15100.4]
  assign RetimeWrapper_15_io_flow = io_enable; // @[package.scala 95:18:@15102.4]
  assign RetimeWrapper_15_io_in = allDone & _T_562; // @[package.scala 94:16:@15101.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_548 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_562 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_548 <= 1'h0;
    end else begin
      _T_548 <= _T_545;
    end
    if (reset) begin
      _T_562 <= 1'h0;
    end else begin
      _T_562 <= _T_545;
    end
  end
endmodule
module RetimeWrapper_178( // @[:@16410.2]
  input         clock, // @[:@16411.4]
  input         reset, // @[:@16412.4]
  input         io_flow, // @[:@16413.4]
  input  [31:0] io_in, // @[:@16413.4]
  output [31:0] io_out // @[:@16413.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16415.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16415.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16415.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16415.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16415.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16415.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@16415.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16428.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16427.4]
  assign sr_init = 32'h6; // @[RetimeShiftRegister.scala 19:16:@16426.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16425.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16424.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16422.4]
endmodule
module NBufCtr_9( // @[:@16430.2]
  input         clock, // @[:@16431.4]
  input         reset, // @[:@16432.4]
  input         io_input_countUp, // @[:@16433.4]
  input         io_input_enable, // @[:@16433.4]
  output [31:0] io_output_count // @[:@16433.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@16470.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@16470.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@16470.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@16470.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@16470.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@16475.4 package.scala 96:25:@16476.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@16436.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@16437.4]
  wire  _T_21; // @[Counter.scala 49:55:@16438.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@16439.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@16440.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@16441.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@16442.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@16443.4]
  wire  _T_33; // @[Counter.scala 51:52:@16447.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@16448.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@16449.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@16450.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@16451.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@16452.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@16453.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@16454.4]
  wire  _T_45; // @[Counter.scala 52:70:@16455.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@16457.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@16458.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@16459.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@16460.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@16461.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@16462.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@16465.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@16466.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@16468.4]
  RetimeWrapper_178 RetimeWrapper ( // @[package.scala 93:22:@16470.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@16475.4 package.scala 96:25:@16476.4]
  assign _T_18 = {{1'd0}, _T_66}; // @[Counter.scala 49:32:@16436.4]
  assign _T_19 = _T_18[31:0]; // @[Counter.scala 49:32:@16437.4]
  assign _T_21 = _T_19 >= 32'h7; // @[Counter.scala 49:55:@16438.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@16439.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh7); // @[Counter.scala 49:91:@16440.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh7); // @[Counter.scala 49:91:@16441.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@16442.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@16443.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@16447.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@16448.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@16449.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@16450.4]
  assign _T_39 = _T_33 ? 32'h6 : _T_38; // @[Counter.scala 51:47:@16451.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@16452.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@16453.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@16454.4]
  assign _T_45 = _T_43 >= 32'h7; // @[Counter.scala 52:70:@16455.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@16457.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@16458.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@16459.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@16460.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@16461.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@16462.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@16465.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@16466.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@16468.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@16478.4]
  assign RetimeWrapper_clock = clock; // @[:@16471.4]
  assign RetimeWrapper_reset = reset; // @[:@16472.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@16474.4]
  assign RetimeWrapper_io_in = reset ? 32'h6 : _T_62; // @[package.scala 94:16:@16473.4]
endmodule
module NBufCtr_11( // @[:@16594.2]
  input         clock, // @[:@16595.4]
  input         reset, // @[:@16596.4]
  input         io_input_countUp, // @[:@16597.4]
  input         io_input_enable, // @[:@16597.4]
  output [31:0] io_output_count // @[:@16597.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@16634.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@16634.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@16634.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@16634.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@16634.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@16639.4 package.scala 96:25:@16640.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@16600.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@16601.4]
  wire  _T_21; // @[Counter.scala 49:55:@16602.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@16603.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@16604.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@16605.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@16606.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@16607.4]
  wire  _T_33; // @[Counter.scala 51:52:@16611.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@16612.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@16613.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@16614.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@16615.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@16616.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@16625.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@16626.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@16629.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@16630.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@16632.4]
  RetimeWrapper_178 RetimeWrapper ( // @[package.scala 93:22:@16634.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@16639.4 package.scala 96:25:@16640.4]
  assign _T_18 = _T_66 + 32'h1; // @[Counter.scala 49:32:@16600.4]
  assign _T_19 = _T_66 + 32'h1; // @[Counter.scala 49:32:@16601.4]
  assign _T_21 = _T_19 >= 32'h7; // @[Counter.scala 49:55:@16602.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@16603.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 49:91:@16604.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 49:91:@16605.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@16606.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@16607.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@16611.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@16612.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@16613.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@16614.4]
  assign _T_39 = _T_33 ? 32'h6 : _T_38; // @[Counter.scala 51:47:@16615.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@16616.4]
  assign _T_53 = {{1'd0}, _T_27}; // @[Counter.scala 52:107:@16625.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@16626.4]
  assign _T_58 = _T_21 ? _T_54 : _T_19; // @[Counter.scala 52:45:@16629.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@16630.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@16632.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@16642.4]
  assign RetimeWrapper_clock = clock; // @[:@16635.4]
  assign RetimeWrapper_reset = reset; // @[:@16636.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@16638.4]
  assign RetimeWrapper_io_in = reset ? 32'h6 : _T_62; // @[package.scala 94:16:@16637.4]
endmodule
module NBufCtr_12( // @[:@16676.2]
  input         clock, // @[:@16677.4]
  input         reset, // @[:@16678.4]
  input         io_input_countUp, // @[:@16679.4]
  input         io_input_enable, // @[:@16679.4]
  output [31:0] io_output_count // @[:@16679.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@16716.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@16716.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@16716.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@16716.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@16716.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@16721.4 package.scala 96:25:@16722.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@16682.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@16683.4]
  wire  _T_21; // @[Counter.scala 49:55:@16684.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@16685.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@16686.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@16687.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@16688.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@16689.4]
  wire  _T_33; // @[Counter.scala 51:52:@16693.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@16694.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@16695.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@16696.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@16697.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@16698.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@16699.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@16700.4]
  wire  _T_45; // @[Counter.scala 52:70:@16701.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@16703.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@16704.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@16705.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@16706.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@16707.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@16708.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@16711.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@16712.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@16714.4]
  RetimeWrapper_178 RetimeWrapper ( // @[package.scala 93:22:@16716.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@16721.4 package.scala 96:25:@16722.4]
  assign _T_18 = _T_66 + 32'h2; // @[Counter.scala 49:32:@16682.4]
  assign _T_19 = _T_66 + 32'h2; // @[Counter.scala 49:32:@16683.4]
  assign _T_21 = _T_19 >= 32'h7; // @[Counter.scala 49:55:@16684.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@16685.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 49:91:@16686.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 49:91:@16687.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@16688.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@16689.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@16693.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@16694.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@16695.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@16696.4]
  assign _T_39 = _T_33 ? 32'h6 : _T_38; // @[Counter.scala 51:47:@16697.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@16698.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@16699.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@16700.4]
  assign _T_45 = _T_43 >= 32'h7; // @[Counter.scala 52:70:@16701.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@16703.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@16704.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@16705.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@16706.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@16707.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@16708.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@16711.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@16712.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@16714.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@16724.4]
  assign RetimeWrapper_clock = clock; // @[:@16717.4]
  assign RetimeWrapper_reset = reset; // @[:@16718.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@16720.4]
  assign RetimeWrapper_io_in = reset ? 32'h6 : _T_62; // @[package.scala 94:16:@16719.4]
endmodule
module NBufCtr_13( // @[:@16758.2]
  input         clock, // @[:@16759.4]
  input         reset, // @[:@16760.4]
  input         io_input_countUp, // @[:@16761.4]
  input         io_input_enable, // @[:@16761.4]
  output [31:0] io_output_count // @[:@16761.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@16798.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@16798.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@16798.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@16798.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@16798.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@16803.4 package.scala 96:25:@16804.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@16764.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@16765.4]
  wire  _T_21; // @[Counter.scala 49:55:@16766.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@16767.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@16768.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@16769.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@16770.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@16771.4]
  wire  _T_33; // @[Counter.scala 51:52:@16775.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@16776.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@16777.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@16778.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@16779.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@16780.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@16781.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@16782.4]
  wire  _T_45; // @[Counter.scala 52:70:@16783.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@16785.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@16786.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@16787.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@16788.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@16789.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@16790.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@16793.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@16794.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@16796.4]
  RetimeWrapper_178 RetimeWrapper ( // @[package.scala 93:22:@16798.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@16803.4 package.scala 96:25:@16804.4]
  assign _T_18 = _T_66 + 32'h3; // @[Counter.scala 49:32:@16764.4]
  assign _T_19 = _T_66 + 32'h3; // @[Counter.scala 49:32:@16765.4]
  assign _T_21 = _T_19 >= 32'h7; // @[Counter.scala 49:55:@16766.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@16767.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh4); // @[Counter.scala 49:91:@16768.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh4); // @[Counter.scala 49:91:@16769.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@16770.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@16771.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@16775.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@16776.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@16777.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@16778.4]
  assign _T_39 = _T_33 ? 32'h6 : _T_38; // @[Counter.scala 51:47:@16779.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@16780.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@16781.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@16782.4]
  assign _T_45 = _T_43 >= 32'h7; // @[Counter.scala 52:70:@16783.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@16785.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@16786.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@16787.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@16788.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@16789.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@16790.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@16793.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@16794.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@16796.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@16806.4]
  assign RetimeWrapper_clock = clock; // @[:@16799.4]
  assign RetimeWrapper_reset = reset; // @[:@16800.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@16802.4]
  assign RetimeWrapper_io_in = reset ? 32'h6 : _T_62; // @[package.scala 94:16:@16801.4]
endmodule
module NBufCtr_14( // @[:@16840.2]
  input         clock, // @[:@16841.4]
  input         reset, // @[:@16842.4]
  input         io_input_countUp, // @[:@16843.4]
  input         io_input_enable, // @[:@16843.4]
  output [31:0] io_output_count // @[:@16843.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@16880.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@16880.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@16880.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@16880.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@16880.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@16885.4 package.scala 96:25:@16886.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@16846.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@16847.4]
  wire  _T_21; // @[Counter.scala 49:55:@16848.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@16849.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@16850.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@16851.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@16852.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@16853.4]
  wire  _T_33; // @[Counter.scala 51:52:@16857.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@16858.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@16859.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@16860.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@16861.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@16862.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@16863.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@16864.4]
  wire  _T_45; // @[Counter.scala 52:70:@16865.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@16867.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@16868.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@16869.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@16870.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@16871.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@16872.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@16875.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@16876.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@16878.4]
  RetimeWrapper_178 RetimeWrapper ( // @[package.scala 93:22:@16880.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@16885.4 package.scala 96:25:@16886.4]
  assign _T_18 = _T_66 + 32'h4; // @[Counter.scala 49:32:@16846.4]
  assign _T_19 = _T_66 + 32'h4; // @[Counter.scala 49:32:@16847.4]
  assign _T_21 = _T_19 >= 32'h7; // @[Counter.scala 49:55:@16848.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@16849.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh3); // @[Counter.scala 49:91:@16850.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh3); // @[Counter.scala 49:91:@16851.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@16852.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@16853.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@16857.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@16858.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@16859.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@16860.4]
  assign _T_39 = _T_33 ? 32'h6 : _T_38; // @[Counter.scala 51:47:@16861.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@16862.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@16863.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@16864.4]
  assign _T_45 = _T_43 >= 32'h7; // @[Counter.scala 52:70:@16865.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@16867.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@16868.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@16869.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@16870.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@16871.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@16872.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@16875.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@16876.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@16878.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@16888.4]
  assign RetimeWrapper_clock = clock; // @[:@16881.4]
  assign RetimeWrapper_reset = reset; // @[:@16882.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@16884.4]
  assign RetimeWrapper_io_in = reset ? 32'h6 : _T_62; // @[package.scala 94:16:@16883.4]
endmodule
module NBufCtr_15( // @[:@16922.2]
  input         clock, // @[:@16923.4]
  input         reset, // @[:@16924.4]
  input         io_input_countUp, // @[:@16925.4]
  input         io_input_enable, // @[:@16925.4]
  output [31:0] io_output_count // @[:@16925.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@16962.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@16962.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@16962.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@16962.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@16962.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@16967.4 package.scala 96:25:@16968.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@16928.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@16929.4]
  wire  _T_21; // @[Counter.scala 49:55:@16930.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@16931.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@16932.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@16933.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@16934.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@16935.4]
  wire  _T_33; // @[Counter.scala 51:52:@16939.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@16940.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@16941.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@16942.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@16943.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@16944.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@16945.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@16946.4]
  wire  _T_45; // @[Counter.scala 52:70:@16947.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@16949.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@16950.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@16951.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@16952.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@16953.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@16954.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@16957.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@16958.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@16960.4]
  RetimeWrapper_178 RetimeWrapper ( // @[package.scala 93:22:@16962.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@16967.4 package.scala 96:25:@16968.4]
  assign _T_18 = _T_66 + 32'h5; // @[Counter.scala 49:32:@16928.4]
  assign _T_19 = _T_66 + 32'h5; // @[Counter.scala 49:32:@16929.4]
  assign _T_21 = _T_19 >= 32'h7; // @[Counter.scala 49:55:@16930.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@16931.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh2); // @[Counter.scala 49:91:@16932.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh2); // @[Counter.scala 49:91:@16933.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@16934.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@16935.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@16939.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@16940.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@16941.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@16942.4]
  assign _T_39 = _T_33 ? 32'h6 : _T_38; // @[Counter.scala 51:47:@16943.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@16944.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@16945.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@16946.4]
  assign _T_45 = _T_43 >= 32'h7; // @[Counter.scala 52:70:@16947.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@16949.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@16950.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@16951.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@16952.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@16953.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@16954.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@16957.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@16958.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@16960.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@16970.4]
  assign RetimeWrapper_clock = clock; // @[:@16963.4]
  assign RetimeWrapper_reset = reset; // @[:@16964.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@16966.4]
  assign RetimeWrapper_io_in = reset ? 32'h6 : _T_62; // @[package.scala 94:16:@16965.4]
endmodule
module NBufCtr_16( // @[:@17004.2]
  input         clock, // @[:@17005.4]
  input         reset, // @[:@17006.4]
  input         io_input_countUp, // @[:@17007.4]
  input         io_input_enable, // @[:@17007.4]
  output [31:0] io_output_count // @[:@17007.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@17044.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@17044.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@17044.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@17044.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@17044.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@17049.4 package.scala 96:25:@17050.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@17010.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@17011.4]
  wire  _T_21; // @[Counter.scala 49:55:@17012.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@17013.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@17014.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@17015.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@17016.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@17017.4]
  wire  _T_33; // @[Counter.scala 51:52:@17021.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@17022.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@17023.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@17024.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@17025.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@17026.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@17027.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@17028.4]
  wire  _T_45; // @[Counter.scala 52:70:@17029.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@17031.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@17032.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@17033.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@17034.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@17035.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@17036.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@17039.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@17040.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@17042.4]
  RetimeWrapper_178 RetimeWrapper ( // @[package.scala 93:22:@17044.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@17049.4 package.scala 96:25:@17050.4]
  assign _T_18 = _T_66 + 32'h6; // @[Counter.scala 49:32:@17010.4]
  assign _T_19 = _T_66 + 32'h6; // @[Counter.scala 49:32:@17011.4]
  assign _T_21 = _T_19 >= 32'h7; // @[Counter.scala 49:55:@17012.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@17013.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 49:91:@17014.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 49:91:@17015.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@17016.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@17017.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@17021.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@17022.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@17023.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@17024.4]
  assign _T_39 = _T_33 ? 32'h6 : _T_38; // @[Counter.scala 51:47:@17025.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@17026.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@17027.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@17028.4]
  assign _T_45 = _T_43 >= 32'h7; // @[Counter.scala 52:70:@17029.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@17031.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 52:121:@17032.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@17033.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@17034.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@17035.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@17036.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@17039.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@17040.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@17042.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@17052.4]
  assign RetimeWrapper_clock = clock; // @[:@17045.4]
  assign RetimeWrapper_reset = reset; // @[:@17046.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@17048.4]
  assign RetimeWrapper_io_in = reset ? 32'h6 : _T_62; // @[package.scala 94:16:@17047.4]
endmodule
module NBufController_3( // @[:@17054.2]
  input        clock, // @[:@17055.4]
  input        reset, // @[:@17056.4]
  input        io_sEn_0, // @[:@17057.4]
  input        io_sEn_1, // @[:@17057.4]
  input        io_sEn_2, // @[:@17057.4]
  input        io_sEn_3, // @[:@17057.4]
  input        io_sEn_4, // @[:@17057.4]
  input        io_sEn_5, // @[:@17057.4]
  input        io_sEn_6, // @[:@17057.4]
  input        io_sDone_0, // @[:@17057.4]
  input        io_sDone_1, // @[:@17057.4]
  input        io_sDone_2, // @[:@17057.4]
  input        io_sDone_3, // @[:@17057.4]
  input        io_sDone_4, // @[:@17057.4]
  input        io_sDone_5, // @[:@17057.4]
  input        io_sDone_6, // @[:@17057.4]
  output [3:0] io_statesInW_0, // @[:@17057.4]
  output [3:0] io_statesInR_1, // @[:@17057.4]
  output [3:0] io_statesInR_2, // @[:@17057.4]
  output [3:0] io_statesInR_3, // @[:@17057.4]
  output [3:0] io_statesInR_4, // @[:@17057.4]
  output [3:0] io_statesInR_5, // @[:@17057.4]
  output [3:0] io_statesInR_6 // @[:@17057.4]
);
  wire  sEn_latch_0_clock; // @[NBuffers.scala 21:52:@17059.4]
  wire  sEn_latch_0_reset; // @[NBuffers.scala 21:52:@17059.4]
  wire  sEn_latch_0_io_input_set; // @[NBuffers.scala 21:52:@17059.4]
  wire  sEn_latch_0_io_input_reset; // @[NBuffers.scala 21:52:@17059.4]
  wire  sEn_latch_0_io_input_asyn_reset; // @[NBuffers.scala 21:52:@17059.4]
  wire  sEn_latch_0_io_output; // @[NBuffers.scala 21:52:@17059.4]
  wire  sEn_latch_1_clock; // @[NBuffers.scala 21:52:@17062.4]
  wire  sEn_latch_1_reset; // @[NBuffers.scala 21:52:@17062.4]
  wire  sEn_latch_1_io_input_set; // @[NBuffers.scala 21:52:@17062.4]
  wire  sEn_latch_1_io_input_reset; // @[NBuffers.scala 21:52:@17062.4]
  wire  sEn_latch_1_io_input_asyn_reset; // @[NBuffers.scala 21:52:@17062.4]
  wire  sEn_latch_1_io_output; // @[NBuffers.scala 21:52:@17062.4]
  wire  sEn_latch_2_clock; // @[NBuffers.scala 21:52:@17065.4]
  wire  sEn_latch_2_reset; // @[NBuffers.scala 21:52:@17065.4]
  wire  sEn_latch_2_io_input_set; // @[NBuffers.scala 21:52:@17065.4]
  wire  sEn_latch_2_io_input_reset; // @[NBuffers.scala 21:52:@17065.4]
  wire  sEn_latch_2_io_input_asyn_reset; // @[NBuffers.scala 21:52:@17065.4]
  wire  sEn_latch_2_io_output; // @[NBuffers.scala 21:52:@17065.4]
  wire  sEn_latch_3_clock; // @[NBuffers.scala 21:52:@17068.4]
  wire  sEn_latch_3_reset; // @[NBuffers.scala 21:52:@17068.4]
  wire  sEn_latch_3_io_input_set; // @[NBuffers.scala 21:52:@17068.4]
  wire  sEn_latch_3_io_input_reset; // @[NBuffers.scala 21:52:@17068.4]
  wire  sEn_latch_3_io_input_asyn_reset; // @[NBuffers.scala 21:52:@17068.4]
  wire  sEn_latch_3_io_output; // @[NBuffers.scala 21:52:@17068.4]
  wire  sEn_latch_4_clock; // @[NBuffers.scala 21:52:@17071.4]
  wire  sEn_latch_4_reset; // @[NBuffers.scala 21:52:@17071.4]
  wire  sEn_latch_4_io_input_set; // @[NBuffers.scala 21:52:@17071.4]
  wire  sEn_latch_4_io_input_reset; // @[NBuffers.scala 21:52:@17071.4]
  wire  sEn_latch_4_io_input_asyn_reset; // @[NBuffers.scala 21:52:@17071.4]
  wire  sEn_latch_4_io_output; // @[NBuffers.scala 21:52:@17071.4]
  wire  sEn_latch_5_clock; // @[NBuffers.scala 21:52:@17074.4]
  wire  sEn_latch_5_reset; // @[NBuffers.scala 21:52:@17074.4]
  wire  sEn_latch_5_io_input_set; // @[NBuffers.scala 21:52:@17074.4]
  wire  sEn_latch_5_io_input_reset; // @[NBuffers.scala 21:52:@17074.4]
  wire  sEn_latch_5_io_input_asyn_reset; // @[NBuffers.scala 21:52:@17074.4]
  wire  sEn_latch_5_io_output; // @[NBuffers.scala 21:52:@17074.4]
  wire  sEn_latch_6_clock; // @[NBuffers.scala 21:52:@17077.4]
  wire  sEn_latch_6_reset; // @[NBuffers.scala 21:52:@17077.4]
  wire  sEn_latch_6_io_input_set; // @[NBuffers.scala 21:52:@17077.4]
  wire  sEn_latch_6_io_input_reset; // @[NBuffers.scala 21:52:@17077.4]
  wire  sEn_latch_6_io_input_asyn_reset; // @[NBuffers.scala 21:52:@17077.4]
  wire  sEn_latch_6_io_output; // @[NBuffers.scala 21:52:@17077.4]
  wire  sDone_latch_0_clock; // @[NBuffers.scala 22:54:@17080.4]
  wire  sDone_latch_0_reset; // @[NBuffers.scala 22:54:@17080.4]
  wire  sDone_latch_0_io_input_set; // @[NBuffers.scala 22:54:@17080.4]
  wire  sDone_latch_0_io_input_reset; // @[NBuffers.scala 22:54:@17080.4]
  wire  sDone_latch_0_io_input_asyn_reset; // @[NBuffers.scala 22:54:@17080.4]
  wire  sDone_latch_0_io_output; // @[NBuffers.scala 22:54:@17080.4]
  wire  sDone_latch_1_clock; // @[NBuffers.scala 22:54:@17083.4]
  wire  sDone_latch_1_reset; // @[NBuffers.scala 22:54:@17083.4]
  wire  sDone_latch_1_io_input_set; // @[NBuffers.scala 22:54:@17083.4]
  wire  sDone_latch_1_io_input_reset; // @[NBuffers.scala 22:54:@17083.4]
  wire  sDone_latch_1_io_input_asyn_reset; // @[NBuffers.scala 22:54:@17083.4]
  wire  sDone_latch_1_io_output; // @[NBuffers.scala 22:54:@17083.4]
  wire  sDone_latch_2_clock; // @[NBuffers.scala 22:54:@17086.4]
  wire  sDone_latch_2_reset; // @[NBuffers.scala 22:54:@17086.4]
  wire  sDone_latch_2_io_input_set; // @[NBuffers.scala 22:54:@17086.4]
  wire  sDone_latch_2_io_input_reset; // @[NBuffers.scala 22:54:@17086.4]
  wire  sDone_latch_2_io_input_asyn_reset; // @[NBuffers.scala 22:54:@17086.4]
  wire  sDone_latch_2_io_output; // @[NBuffers.scala 22:54:@17086.4]
  wire  sDone_latch_3_clock; // @[NBuffers.scala 22:54:@17089.4]
  wire  sDone_latch_3_reset; // @[NBuffers.scala 22:54:@17089.4]
  wire  sDone_latch_3_io_input_set; // @[NBuffers.scala 22:54:@17089.4]
  wire  sDone_latch_3_io_input_reset; // @[NBuffers.scala 22:54:@17089.4]
  wire  sDone_latch_3_io_input_asyn_reset; // @[NBuffers.scala 22:54:@17089.4]
  wire  sDone_latch_3_io_output; // @[NBuffers.scala 22:54:@17089.4]
  wire  sDone_latch_4_clock; // @[NBuffers.scala 22:54:@17092.4]
  wire  sDone_latch_4_reset; // @[NBuffers.scala 22:54:@17092.4]
  wire  sDone_latch_4_io_input_set; // @[NBuffers.scala 22:54:@17092.4]
  wire  sDone_latch_4_io_input_reset; // @[NBuffers.scala 22:54:@17092.4]
  wire  sDone_latch_4_io_input_asyn_reset; // @[NBuffers.scala 22:54:@17092.4]
  wire  sDone_latch_4_io_output; // @[NBuffers.scala 22:54:@17092.4]
  wire  sDone_latch_5_clock; // @[NBuffers.scala 22:54:@17095.4]
  wire  sDone_latch_5_reset; // @[NBuffers.scala 22:54:@17095.4]
  wire  sDone_latch_5_io_input_set; // @[NBuffers.scala 22:54:@17095.4]
  wire  sDone_latch_5_io_input_reset; // @[NBuffers.scala 22:54:@17095.4]
  wire  sDone_latch_5_io_input_asyn_reset; // @[NBuffers.scala 22:54:@17095.4]
  wire  sDone_latch_5_io_output; // @[NBuffers.scala 22:54:@17095.4]
  wire  sDone_latch_6_clock; // @[NBuffers.scala 22:54:@17098.4]
  wire  sDone_latch_6_reset; // @[NBuffers.scala 22:54:@17098.4]
  wire  sDone_latch_6_io_input_set; // @[NBuffers.scala 22:54:@17098.4]
  wire  sDone_latch_6_io_input_reset; // @[NBuffers.scala 22:54:@17098.4]
  wire  sDone_latch_6_io_input_asyn_reset; // @[NBuffers.scala 22:54:@17098.4]
  wire  sDone_latch_6_io_output; // @[NBuffers.scala 22:54:@17098.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@17105.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@17105.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@17105.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@17105.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@17105.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@17113.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@17113.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@17113.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@17113.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@17113.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@17122.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@17122.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@17122.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@17122.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@17122.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@17130.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@17130.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@17130.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@17130.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@17130.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@17141.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@17141.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@17141.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@17141.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@17141.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@17149.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@17149.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@17149.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@17149.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@17149.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@17158.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@17158.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@17158.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@17158.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@17158.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@17166.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@17166.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@17166.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@17166.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@17166.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@17177.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@17177.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@17177.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@17177.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@17177.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@17185.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@17185.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@17185.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@17185.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@17185.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@17194.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@17194.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@17194.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@17194.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@17194.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@17202.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@17202.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@17202.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@17202.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@17202.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@17213.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@17213.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@17213.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@17213.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@17213.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@17221.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@17221.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@17221.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@17221.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@17221.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@17230.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@17230.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@17230.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@17230.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@17230.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@17238.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@17238.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@17238.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@17238.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@17238.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@17249.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@17249.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@17249.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@17249.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@17249.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@17257.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@17257.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@17257.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@17257.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@17257.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@17266.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@17266.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@17266.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@17266.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@17266.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@17274.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@17274.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@17274.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@17274.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@17274.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@17285.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@17285.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@17285.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@17285.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@17285.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@17293.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@17293.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@17293.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@17293.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@17293.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@17302.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@17302.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@17302.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@17302.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@17302.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@17310.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@17310.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@17310.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@17310.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@17310.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@17321.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@17321.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@17321.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@17321.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@17321.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@17329.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@17329.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@17329.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@17329.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@17329.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@17338.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@17338.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@17338.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@17338.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@17338.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@17346.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@17346.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@17346.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@17346.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@17346.4]
  wire  NBufCtr_clock; // @[NBuffers.scala 40:19:@17387.4]
  wire  NBufCtr_reset; // @[NBuffers.scala 40:19:@17387.4]
  wire  NBufCtr_io_input_countUp; // @[NBuffers.scala 40:19:@17387.4]
  wire  NBufCtr_io_input_enable; // @[NBuffers.scala 40:19:@17387.4]
  wire [31:0] NBufCtr_io_output_count; // @[NBuffers.scala 40:19:@17387.4]
  wire  statesInR_0_clock; // @[NBuffers.scala 50:19:@17398.4]
  wire  statesInR_0_reset; // @[NBuffers.scala 50:19:@17398.4]
  wire  statesInR_0_io_input_countUp; // @[NBuffers.scala 50:19:@17398.4]
  wire  statesInR_0_io_input_enable; // @[NBuffers.scala 50:19:@17398.4]
  wire [31:0] statesInR_0_io_output_count; // @[NBuffers.scala 50:19:@17398.4]
  wire  statesInR_1_clock; // @[NBuffers.scala 50:19:@17409.4]
  wire  statesInR_1_reset; // @[NBuffers.scala 50:19:@17409.4]
  wire  statesInR_1_io_input_countUp; // @[NBuffers.scala 50:19:@17409.4]
  wire  statesInR_1_io_input_enable; // @[NBuffers.scala 50:19:@17409.4]
  wire [31:0] statesInR_1_io_output_count; // @[NBuffers.scala 50:19:@17409.4]
  wire  statesInR_2_clock; // @[NBuffers.scala 50:19:@17420.4]
  wire  statesInR_2_reset; // @[NBuffers.scala 50:19:@17420.4]
  wire  statesInR_2_io_input_countUp; // @[NBuffers.scala 50:19:@17420.4]
  wire  statesInR_2_io_input_enable; // @[NBuffers.scala 50:19:@17420.4]
  wire [31:0] statesInR_2_io_output_count; // @[NBuffers.scala 50:19:@17420.4]
  wire  statesInR_3_clock; // @[NBuffers.scala 50:19:@17431.4]
  wire  statesInR_3_reset; // @[NBuffers.scala 50:19:@17431.4]
  wire  statesInR_3_io_input_countUp; // @[NBuffers.scala 50:19:@17431.4]
  wire  statesInR_3_io_input_enable; // @[NBuffers.scala 50:19:@17431.4]
  wire [31:0] statesInR_3_io_output_count; // @[NBuffers.scala 50:19:@17431.4]
  wire  statesInR_4_clock; // @[NBuffers.scala 50:19:@17442.4]
  wire  statesInR_4_reset; // @[NBuffers.scala 50:19:@17442.4]
  wire  statesInR_4_io_input_countUp; // @[NBuffers.scala 50:19:@17442.4]
  wire  statesInR_4_io_input_enable; // @[NBuffers.scala 50:19:@17442.4]
  wire [31:0] statesInR_4_io_output_count; // @[NBuffers.scala 50:19:@17442.4]
  wire  statesInR_5_clock; // @[NBuffers.scala 50:19:@17453.4]
  wire  statesInR_5_reset; // @[NBuffers.scala 50:19:@17453.4]
  wire  statesInR_5_io_input_countUp; // @[NBuffers.scala 50:19:@17453.4]
  wire  statesInR_5_io_input_enable; // @[NBuffers.scala 50:19:@17453.4]
  wire [31:0] statesInR_5_io_output_count; // @[NBuffers.scala 50:19:@17453.4]
  wire  statesInR_6_clock; // @[NBuffers.scala 50:19:@17464.4]
  wire  statesInR_6_reset; // @[NBuffers.scala 50:19:@17464.4]
  wire  statesInR_6_io_input_countUp; // @[NBuffers.scala 50:19:@17464.4]
  wire  statesInR_6_io_input_enable; // @[NBuffers.scala 50:19:@17464.4]
  wire [31:0] statesInR_6_io_output_count; // @[NBuffers.scala 50:19:@17464.4]
  wire  _T_33; // @[NBuffers.scala 26:46:@17102.4]
  wire  _T_48; // @[NBuffers.scala 26:46:@17138.4]
  wire  _T_63; // @[NBuffers.scala 26:46:@17174.4]
  wire  _T_78; // @[NBuffers.scala 26:46:@17210.4]
  wire  _T_93; // @[NBuffers.scala 26:46:@17246.4]
  wire  _T_108; // @[NBuffers.scala 26:46:@17282.4]
  wire  _T_123; // @[NBuffers.scala 26:46:@17318.4]
  wire  _T_137; // @[NBuffers.scala 33:64:@17354.4]
  wire  _T_138; // @[NBuffers.scala 33:64:@17355.4]
  wire  _T_139; // @[NBuffers.scala 33:64:@17356.4]
  wire  _T_140; // @[NBuffers.scala 33:64:@17357.4]
  wire  _T_141; // @[NBuffers.scala 33:64:@17358.4]
  wire  anyEnabled; // @[NBuffers.scala 33:64:@17359.4]
  wire  _T_142; // @[NBuffers.scala 34:124:@17360.4]
  wire  _T_143; // @[NBuffers.scala 34:104:@17361.4]
  wire  _T_144; // @[NBuffers.scala 34:124:@17362.4]
  wire  _T_145; // @[NBuffers.scala 34:104:@17363.4]
  wire  _T_146; // @[NBuffers.scala 34:124:@17364.4]
  wire  _T_147; // @[NBuffers.scala 34:104:@17365.4]
  wire  _T_148; // @[NBuffers.scala 34:124:@17366.4]
  wire  _T_149; // @[NBuffers.scala 34:104:@17367.4]
  wire  _T_150; // @[NBuffers.scala 34:124:@17368.4]
  wire  _T_151; // @[NBuffers.scala 34:104:@17369.4]
  wire  _T_152; // @[NBuffers.scala 34:124:@17370.4]
  wire  _T_153; // @[NBuffers.scala 34:104:@17371.4]
  wire  _T_154; // @[NBuffers.scala 34:124:@17372.4]
  wire  _T_155; // @[NBuffers.scala 34:104:@17373.4]
  wire  _T_156; // @[NBuffers.scala 34:150:@17374.4]
  wire  _T_157; // @[NBuffers.scala 34:150:@17375.4]
  wire  _T_158; // @[NBuffers.scala 34:150:@17376.4]
  wire  _T_159; // @[NBuffers.scala 34:150:@17377.4]
  wire  _T_160; // @[NBuffers.scala 34:150:@17378.4]
  wire  _T_161; // @[NBuffers.scala 34:150:@17379.4]
  wire  _T_162; // @[NBuffers.scala 34:154:@17380.4]
  wire  _T_164; // @[package.scala 100:49:@17381.4]
  reg  _T_167; // @[package.scala 48:56:@17382.4]
  reg [31:0] _RAND_0;
  SRFF sEn_latch_0 ( // @[NBuffers.scala 21:52:@17059.4]
    .clock(sEn_latch_0_clock),
    .reset(sEn_latch_0_reset),
    .io_input_set(sEn_latch_0_io_input_set),
    .io_input_reset(sEn_latch_0_io_input_reset),
    .io_input_asyn_reset(sEn_latch_0_io_input_asyn_reset),
    .io_output(sEn_latch_0_io_output)
  );
  SRFF sEn_latch_1 ( // @[NBuffers.scala 21:52:@17062.4]
    .clock(sEn_latch_1_clock),
    .reset(sEn_latch_1_reset),
    .io_input_set(sEn_latch_1_io_input_set),
    .io_input_reset(sEn_latch_1_io_input_reset),
    .io_input_asyn_reset(sEn_latch_1_io_input_asyn_reset),
    .io_output(sEn_latch_1_io_output)
  );
  SRFF sEn_latch_2 ( // @[NBuffers.scala 21:52:@17065.4]
    .clock(sEn_latch_2_clock),
    .reset(sEn_latch_2_reset),
    .io_input_set(sEn_latch_2_io_input_set),
    .io_input_reset(sEn_latch_2_io_input_reset),
    .io_input_asyn_reset(sEn_latch_2_io_input_asyn_reset),
    .io_output(sEn_latch_2_io_output)
  );
  SRFF sEn_latch_3 ( // @[NBuffers.scala 21:52:@17068.4]
    .clock(sEn_latch_3_clock),
    .reset(sEn_latch_3_reset),
    .io_input_set(sEn_latch_3_io_input_set),
    .io_input_reset(sEn_latch_3_io_input_reset),
    .io_input_asyn_reset(sEn_latch_3_io_input_asyn_reset),
    .io_output(sEn_latch_3_io_output)
  );
  SRFF sEn_latch_4 ( // @[NBuffers.scala 21:52:@17071.4]
    .clock(sEn_latch_4_clock),
    .reset(sEn_latch_4_reset),
    .io_input_set(sEn_latch_4_io_input_set),
    .io_input_reset(sEn_latch_4_io_input_reset),
    .io_input_asyn_reset(sEn_latch_4_io_input_asyn_reset),
    .io_output(sEn_latch_4_io_output)
  );
  SRFF sEn_latch_5 ( // @[NBuffers.scala 21:52:@17074.4]
    .clock(sEn_latch_5_clock),
    .reset(sEn_latch_5_reset),
    .io_input_set(sEn_latch_5_io_input_set),
    .io_input_reset(sEn_latch_5_io_input_reset),
    .io_input_asyn_reset(sEn_latch_5_io_input_asyn_reset),
    .io_output(sEn_latch_5_io_output)
  );
  SRFF sEn_latch_6 ( // @[NBuffers.scala 21:52:@17077.4]
    .clock(sEn_latch_6_clock),
    .reset(sEn_latch_6_reset),
    .io_input_set(sEn_latch_6_io_input_set),
    .io_input_reset(sEn_latch_6_io_input_reset),
    .io_input_asyn_reset(sEn_latch_6_io_input_asyn_reset),
    .io_output(sEn_latch_6_io_output)
  );
  SRFF sDone_latch_0 ( // @[NBuffers.scala 22:54:@17080.4]
    .clock(sDone_latch_0_clock),
    .reset(sDone_latch_0_reset),
    .io_input_set(sDone_latch_0_io_input_set),
    .io_input_reset(sDone_latch_0_io_input_reset),
    .io_input_asyn_reset(sDone_latch_0_io_input_asyn_reset),
    .io_output(sDone_latch_0_io_output)
  );
  SRFF sDone_latch_1 ( // @[NBuffers.scala 22:54:@17083.4]
    .clock(sDone_latch_1_clock),
    .reset(sDone_latch_1_reset),
    .io_input_set(sDone_latch_1_io_input_set),
    .io_input_reset(sDone_latch_1_io_input_reset),
    .io_input_asyn_reset(sDone_latch_1_io_input_asyn_reset),
    .io_output(sDone_latch_1_io_output)
  );
  SRFF sDone_latch_2 ( // @[NBuffers.scala 22:54:@17086.4]
    .clock(sDone_latch_2_clock),
    .reset(sDone_latch_2_reset),
    .io_input_set(sDone_latch_2_io_input_set),
    .io_input_reset(sDone_latch_2_io_input_reset),
    .io_input_asyn_reset(sDone_latch_2_io_input_asyn_reset),
    .io_output(sDone_latch_2_io_output)
  );
  SRFF sDone_latch_3 ( // @[NBuffers.scala 22:54:@17089.4]
    .clock(sDone_latch_3_clock),
    .reset(sDone_latch_3_reset),
    .io_input_set(sDone_latch_3_io_input_set),
    .io_input_reset(sDone_latch_3_io_input_reset),
    .io_input_asyn_reset(sDone_latch_3_io_input_asyn_reset),
    .io_output(sDone_latch_3_io_output)
  );
  SRFF sDone_latch_4 ( // @[NBuffers.scala 22:54:@17092.4]
    .clock(sDone_latch_4_clock),
    .reset(sDone_latch_4_reset),
    .io_input_set(sDone_latch_4_io_input_set),
    .io_input_reset(sDone_latch_4_io_input_reset),
    .io_input_asyn_reset(sDone_latch_4_io_input_asyn_reset),
    .io_output(sDone_latch_4_io_output)
  );
  SRFF sDone_latch_5 ( // @[NBuffers.scala 22:54:@17095.4]
    .clock(sDone_latch_5_clock),
    .reset(sDone_latch_5_reset),
    .io_input_set(sDone_latch_5_io_input_set),
    .io_input_reset(sDone_latch_5_io_input_reset),
    .io_input_asyn_reset(sDone_latch_5_io_input_asyn_reset),
    .io_output(sDone_latch_5_io_output)
  );
  SRFF sDone_latch_6 ( // @[NBuffers.scala 22:54:@17098.4]
    .clock(sDone_latch_6_clock),
    .reset(sDone_latch_6_reset),
    .io_input_set(sDone_latch_6_io_input_set),
    .io_input_reset(sDone_latch_6_io_input_reset),
    .io_input_asyn_reset(sDone_latch_6_io_input_asyn_reset),
    .io_output(sDone_latch_6_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@17105.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@17113.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@17122.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@17130.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@17141.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@17149.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@17158.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@17166.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@17177.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@17185.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@17194.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 ( // @[package.scala 93:22:@17202.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper RetimeWrapper_12 ( // @[package.scala 93:22:@17213.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 ( // @[package.scala 93:22:@17221.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@17230.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@17238.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 ( // @[package.scala 93:22:@17249.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper RetimeWrapper_17 ( // @[package.scala 93:22:@17257.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 ( // @[package.scala 93:22:@17266.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper RetimeWrapper_19 ( // @[package.scala 93:22:@17274.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper RetimeWrapper_20 ( // @[package.scala 93:22:@17285.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper RetimeWrapper_21 ( // @[package.scala 93:22:@17293.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper RetimeWrapper_22 ( // @[package.scala 93:22:@17302.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper RetimeWrapper_23 ( // @[package.scala 93:22:@17310.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper RetimeWrapper_24 ( // @[package.scala 93:22:@17321.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@17329.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper RetimeWrapper_26 ( // @[package.scala 93:22:@17338.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper RetimeWrapper_27 ( // @[package.scala 93:22:@17346.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  NBufCtr_9 NBufCtr ( // @[NBuffers.scala 40:19:@17387.4]
    .clock(NBufCtr_clock),
    .reset(NBufCtr_reset),
    .io_input_countUp(NBufCtr_io_input_countUp),
    .io_input_enable(NBufCtr_io_input_enable),
    .io_output_count(NBufCtr_io_output_count)
  );
  NBufCtr_9 statesInR_0 ( // @[NBuffers.scala 50:19:@17398.4]
    .clock(statesInR_0_clock),
    .reset(statesInR_0_reset),
    .io_input_countUp(statesInR_0_io_input_countUp),
    .io_input_enable(statesInR_0_io_input_enable),
    .io_output_count(statesInR_0_io_output_count)
  );
  NBufCtr_11 statesInR_1 ( // @[NBuffers.scala 50:19:@17409.4]
    .clock(statesInR_1_clock),
    .reset(statesInR_1_reset),
    .io_input_countUp(statesInR_1_io_input_countUp),
    .io_input_enable(statesInR_1_io_input_enable),
    .io_output_count(statesInR_1_io_output_count)
  );
  NBufCtr_12 statesInR_2 ( // @[NBuffers.scala 50:19:@17420.4]
    .clock(statesInR_2_clock),
    .reset(statesInR_2_reset),
    .io_input_countUp(statesInR_2_io_input_countUp),
    .io_input_enable(statesInR_2_io_input_enable),
    .io_output_count(statesInR_2_io_output_count)
  );
  NBufCtr_13 statesInR_3 ( // @[NBuffers.scala 50:19:@17431.4]
    .clock(statesInR_3_clock),
    .reset(statesInR_3_reset),
    .io_input_countUp(statesInR_3_io_input_countUp),
    .io_input_enable(statesInR_3_io_input_enable),
    .io_output_count(statesInR_3_io_output_count)
  );
  NBufCtr_14 statesInR_4 ( // @[NBuffers.scala 50:19:@17442.4]
    .clock(statesInR_4_clock),
    .reset(statesInR_4_reset),
    .io_input_countUp(statesInR_4_io_input_countUp),
    .io_input_enable(statesInR_4_io_input_enable),
    .io_output_count(statesInR_4_io_output_count)
  );
  NBufCtr_15 statesInR_5 ( // @[NBuffers.scala 50:19:@17453.4]
    .clock(statesInR_5_clock),
    .reset(statesInR_5_reset),
    .io_input_countUp(statesInR_5_io_input_countUp),
    .io_input_enable(statesInR_5_io_input_enable),
    .io_output_count(statesInR_5_io_output_count)
  );
  NBufCtr_16 statesInR_6 ( // @[NBuffers.scala 50:19:@17464.4]
    .clock(statesInR_6_clock),
    .reset(statesInR_6_reset),
    .io_input_countUp(statesInR_6_io_input_countUp),
    .io_input_enable(statesInR_6_io_input_enable),
    .io_output_count(statesInR_6_io_output_count)
  );
  assign _T_33 = io_sDone_0 == 1'h0; // @[NBuffers.scala 26:46:@17102.4]
  assign _T_48 = io_sDone_1 == 1'h0; // @[NBuffers.scala 26:46:@17138.4]
  assign _T_63 = io_sDone_2 == 1'h0; // @[NBuffers.scala 26:46:@17174.4]
  assign _T_78 = io_sDone_3 == 1'h0; // @[NBuffers.scala 26:46:@17210.4]
  assign _T_93 = io_sDone_4 == 1'h0; // @[NBuffers.scala 26:46:@17246.4]
  assign _T_108 = io_sDone_5 == 1'h0; // @[NBuffers.scala 26:46:@17282.4]
  assign _T_123 = io_sDone_6 == 1'h0; // @[NBuffers.scala 26:46:@17318.4]
  assign _T_137 = sEn_latch_0_io_output | sEn_latch_1_io_output; // @[NBuffers.scala 33:64:@17354.4]
  assign _T_138 = _T_137 | sEn_latch_2_io_output; // @[NBuffers.scala 33:64:@17355.4]
  assign _T_139 = _T_138 | sEn_latch_3_io_output; // @[NBuffers.scala 33:64:@17356.4]
  assign _T_140 = _T_139 | sEn_latch_4_io_output; // @[NBuffers.scala 33:64:@17357.4]
  assign _T_141 = _T_140 | sEn_latch_5_io_output; // @[NBuffers.scala 33:64:@17358.4]
  assign anyEnabled = _T_141 | sEn_latch_6_io_output; // @[NBuffers.scala 33:64:@17359.4]
  assign _T_142 = sDone_latch_0_io_output | io_sDone_0; // @[NBuffers.scala 34:124:@17360.4]
  assign _T_143 = sEn_latch_0_io_output == _T_142; // @[NBuffers.scala 34:104:@17361.4]
  assign _T_144 = sDone_latch_1_io_output | io_sDone_1; // @[NBuffers.scala 34:124:@17362.4]
  assign _T_145 = sEn_latch_1_io_output == _T_144; // @[NBuffers.scala 34:104:@17363.4]
  assign _T_146 = sDone_latch_2_io_output | io_sDone_2; // @[NBuffers.scala 34:124:@17364.4]
  assign _T_147 = sEn_latch_2_io_output == _T_146; // @[NBuffers.scala 34:104:@17365.4]
  assign _T_148 = sDone_latch_3_io_output | io_sDone_3; // @[NBuffers.scala 34:124:@17366.4]
  assign _T_149 = sEn_latch_3_io_output == _T_148; // @[NBuffers.scala 34:104:@17367.4]
  assign _T_150 = sDone_latch_4_io_output | io_sDone_4; // @[NBuffers.scala 34:124:@17368.4]
  assign _T_151 = sEn_latch_4_io_output == _T_150; // @[NBuffers.scala 34:104:@17369.4]
  assign _T_152 = sDone_latch_5_io_output | io_sDone_5; // @[NBuffers.scala 34:124:@17370.4]
  assign _T_153 = sEn_latch_5_io_output == _T_152; // @[NBuffers.scala 34:104:@17371.4]
  assign _T_154 = sDone_latch_6_io_output | io_sDone_6; // @[NBuffers.scala 34:124:@17372.4]
  assign _T_155 = sEn_latch_6_io_output == _T_154; // @[NBuffers.scala 34:104:@17373.4]
  assign _T_156 = _T_143 & _T_145; // @[NBuffers.scala 34:150:@17374.4]
  assign _T_157 = _T_156 & _T_147; // @[NBuffers.scala 34:150:@17375.4]
  assign _T_158 = _T_157 & _T_149; // @[NBuffers.scala 34:150:@17376.4]
  assign _T_159 = _T_158 & _T_151; // @[NBuffers.scala 34:150:@17377.4]
  assign _T_160 = _T_159 & _T_153; // @[NBuffers.scala 34:150:@17378.4]
  assign _T_161 = _T_160 & _T_155; // @[NBuffers.scala 34:150:@17379.4]
  assign _T_162 = _T_161 & anyEnabled; // @[NBuffers.scala 34:154:@17380.4]
  assign _T_164 = _T_162 == 1'h0; // @[package.scala 100:49:@17381.4]
  assign io_statesInW_0 = NBufCtr_io_output_count[3:0]; // @[NBuffers.scala 44:21:@17397.4]
  assign io_statesInR_1 = statesInR_1_io_output_count[3:0]; // @[NBuffers.scala 54:21:@17419.4]
  assign io_statesInR_2 = statesInR_2_io_output_count[3:0]; // @[NBuffers.scala 54:21:@17430.4]
  assign io_statesInR_3 = statesInR_3_io_output_count[3:0]; // @[NBuffers.scala 54:21:@17441.4]
  assign io_statesInR_4 = statesInR_4_io_output_count[3:0]; // @[NBuffers.scala 54:21:@17452.4]
  assign io_statesInR_5 = statesInR_5_io_output_count[3:0]; // @[NBuffers.scala 54:21:@17463.4]
  assign io_statesInR_6 = statesInR_6_io_output_count[3:0]; // @[NBuffers.scala 54:21:@17474.4]
  assign sEn_latch_0_clock = clock; // @[:@17060.4]
  assign sEn_latch_0_reset = reset; // @[:@17061.4]
  assign sEn_latch_0_io_input_set = io_sEn_0 & _T_33; // @[NBuffers.scala 26:31:@17104.4]
  assign sEn_latch_0_io_input_reset = RetimeWrapper_io_out; // @[NBuffers.scala 27:33:@17112.4]
  assign sEn_latch_0_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[NBuffers.scala 28:38:@17120.4]
  assign sEn_latch_1_clock = clock; // @[:@17063.4]
  assign sEn_latch_1_reset = reset; // @[:@17064.4]
  assign sEn_latch_1_io_input_set = io_sEn_1 & _T_48; // @[NBuffers.scala 26:31:@17140.4]
  assign sEn_latch_1_io_input_reset = RetimeWrapper_4_io_out; // @[NBuffers.scala 27:33:@17148.4]
  assign sEn_latch_1_io_input_asyn_reset = RetimeWrapper_5_io_out; // @[NBuffers.scala 28:38:@17156.4]
  assign sEn_latch_2_clock = clock; // @[:@17066.4]
  assign sEn_latch_2_reset = reset; // @[:@17067.4]
  assign sEn_latch_2_io_input_set = io_sEn_2 & _T_63; // @[NBuffers.scala 26:31:@17176.4]
  assign sEn_latch_2_io_input_reset = RetimeWrapper_8_io_out; // @[NBuffers.scala 27:33:@17184.4]
  assign sEn_latch_2_io_input_asyn_reset = RetimeWrapper_9_io_out; // @[NBuffers.scala 28:38:@17192.4]
  assign sEn_latch_3_clock = clock; // @[:@17069.4]
  assign sEn_latch_3_reset = reset; // @[:@17070.4]
  assign sEn_latch_3_io_input_set = io_sEn_3 & _T_78; // @[NBuffers.scala 26:31:@17212.4]
  assign sEn_latch_3_io_input_reset = RetimeWrapper_12_io_out; // @[NBuffers.scala 27:33:@17220.4]
  assign sEn_latch_3_io_input_asyn_reset = RetimeWrapper_13_io_out; // @[NBuffers.scala 28:38:@17228.4]
  assign sEn_latch_4_clock = clock; // @[:@17072.4]
  assign sEn_latch_4_reset = reset; // @[:@17073.4]
  assign sEn_latch_4_io_input_set = io_sEn_4 & _T_93; // @[NBuffers.scala 26:31:@17248.4]
  assign sEn_latch_4_io_input_reset = RetimeWrapper_16_io_out; // @[NBuffers.scala 27:33:@17256.4]
  assign sEn_latch_4_io_input_asyn_reset = RetimeWrapper_17_io_out; // @[NBuffers.scala 28:38:@17264.4]
  assign sEn_latch_5_clock = clock; // @[:@17075.4]
  assign sEn_latch_5_reset = reset; // @[:@17076.4]
  assign sEn_latch_5_io_input_set = io_sEn_5 & _T_108; // @[NBuffers.scala 26:31:@17284.4]
  assign sEn_latch_5_io_input_reset = RetimeWrapper_20_io_out; // @[NBuffers.scala 27:33:@17292.4]
  assign sEn_latch_5_io_input_asyn_reset = RetimeWrapper_21_io_out; // @[NBuffers.scala 28:38:@17300.4]
  assign sEn_latch_6_clock = clock; // @[:@17078.4]
  assign sEn_latch_6_reset = reset; // @[:@17079.4]
  assign sEn_latch_6_io_input_set = io_sEn_6 & _T_123; // @[NBuffers.scala 26:31:@17320.4]
  assign sEn_latch_6_io_input_reset = RetimeWrapper_24_io_out; // @[NBuffers.scala 27:33:@17328.4]
  assign sEn_latch_6_io_input_asyn_reset = RetimeWrapper_25_io_out; // @[NBuffers.scala 28:38:@17336.4]
  assign sDone_latch_0_clock = clock; // @[:@17081.4]
  assign sDone_latch_0_reset = reset; // @[:@17082.4]
  assign sDone_latch_0_io_input_set = io_sDone_0; // @[NBuffers.scala 29:33:@17121.4]
  assign sDone_latch_0_io_input_reset = RetimeWrapper_2_io_out; // @[NBuffers.scala 30:35:@17129.4]
  assign sDone_latch_0_io_input_asyn_reset = RetimeWrapper_3_io_out; // @[NBuffers.scala 31:40:@17137.4]
  assign sDone_latch_1_clock = clock; // @[:@17084.4]
  assign sDone_latch_1_reset = reset; // @[:@17085.4]
  assign sDone_latch_1_io_input_set = io_sDone_1; // @[NBuffers.scala 29:33:@17157.4]
  assign sDone_latch_1_io_input_reset = RetimeWrapper_6_io_out; // @[NBuffers.scala 30:35:@17165.4]
  assign sDone_latch_1_io_input_asyn_reset = RetimeWrapper_7_io_out; // @[NBuffers.scala 31:40:@17173.4]
  assign sDone_latch_2_clock = clock; // @[:@17087.4]
  assign sDone_latch_2_reset = reset; // @[:@17088.4]
  assign sDone_latch_2_io_input_set = io_sDone_2; // @[NBuffers.scala 29:33:@17193.4]
  assign sDone_latch_2_io_input_reset = RetimeWrapper_10_io_out; // @[NBuffers.scala 30:35:@17201.4]
  assign sDone_latch_2_io_input_asyn_reset = RetimeWrapper_11_io_out; // @[NBuffers.scala 31:40:@17209.4]
  assign sDone_latch_3_clock = clock; // @[:@17090.4]
  assign sDone_latch_3_reset = reset; // @[:@17091.4]
  assign sDone_latch_3_io_input_set = io_sDone_3; // @[NBuffers.scala 29:33:@17229.4]
  assign sDone_latch_3_io_input_reset = RetimeWrapper_14_io_out; // @[NBuffers.scala 30:35:@17237.4]
  assign sDone_latch_3_io_input_asyn_reset = RetimeWrapper_15_io_out; // @[NBuffers.scala 31:40:@17245.4]
  assign sDone_latch_4_clock = clock; // @[:@17093.4]
  assign sDone_latch_4_reset = reset; // @[:@17094.4]
  assign sDone_latch_4_io_input_set = io_sDone_4; // @[NBuffers.scala 29:33:@17265.4]
  assign sDone_latch_4_io_input_reset = RetimeWrapper_18_io_out; // @[NBuffers.scala 30:35:@17273.4]
  assign sDone_latch_4_io_input_asyn_reset = RetimeWrapper_19_io_out; // @[NBuffers.scala 31:40:@17281.4]
  assign sDone_latch_5_clock = clock; // @[:@17096.4]
  assign sDone_latch_5_reset = reset; // @[:@17097.4]
  assign sDone_latch_5_io_input_set = io_sDone_5; // @[NBuffers.scala 29:33:@17301.4]
  assign sDone_latch_5_io_input_reset = RetimeWrapper_22_io_out; // @[NBuffers.scala 30:35:@17309.4]
  assign sDone_latch_5_io_input_asyn_reset = RetimeWrapper_23_io_out; // @[NBuffers.scala 31:40:@17317.4]
  assign sDone_latch_6_clock = clock; // @[:@17099.4]
  assign sDone_latch_6_reset = reset; // @[:@17100.4]
  assign sDone_latch_6_io_input_set = io_sDone_6; // @[NBuffers.scala 29:33:@17337.4]
  assign sDone_latch_6_io_input_reset = RetimeWrapper_26_io_out; // @[NBuffers.scala 30:35:@17345.4]
  assign sDone_latch_6_io_input_asyn_reset = RetimeWrapper_27_io_out; // @[NBuffers.scala 31:40:@17353.4]
  assign RetimeWrapper_clock = clock; // @[:@17106.4]
  assign RetimeWrapper_reset = reset; // @[:@17107.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@17109.4]
  assign RetimeWrapper_io_in = _T_162 & _T_167; // @[package.scala 94:16:@17108.4]
  assign RetimeWrapper_1_clock = clock; // @[:@17114.4]
  assign RetimeWrapper_1_reset = reset; // @[:@17115.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@17117.4]
  assign RetimeWrapper_1_io_in = reset; // @[package.scala 94:16:@17116.4]
  assign RetimeWrapper_2_clock = clock; // @[:@17123.4]
  assign RetimeWrapper_2_reset = reset; // @[:@17124.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@17126.4]
  assign RetimeWrapper_2_io_in = _T_162 & _T_167; // @[package.scala 94:16:@17125.4]
  assign RetimeWrapper_3_clock = clock; // @[:@17131.4]
  assign RetimeWrapper_3_reset = reset; // @[:@17132.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@17134.4]
  assign RetimeWrapper_3_io_in = reset; // @[package.scala 94:16:@17133.4]
  assign RetimeWrapper_4_clock = clock; // @[:@17142.4]
  assign RetimeWrapper_4_reset = reset; // @[:@17143.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@17145.4]
  assign RetimeWrapper_4_io_in = _T_162 & _T_167; // @[package.scala 94:16:@17144.4]
  assign RetimeWrapper_5_clock = clock; // @[:@17150.4]
  assign RetimeWrapper_5_reset = reset; // @[:@17151.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@17153.4]
  assign RetimeWrapper_5_io_in = reset; // @[package.scala 94:16:@17152.4]
  assign RetimeWrapper_6_clock = clock; // @[:@17159.4]
  assign RetimeWrapper_6_reset = reset; // @[:@17160.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@17162.4]
  assign RetimeWrapper_6_io_in = _T_162 & _T_167; // @[package.scala 94:16:@17161.4]
  assign RetimeWrapper_7_clock = clock; // @[:@17167.4]
  assign RetimeWrapper_7_reset = reset; // @[:@17168.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@17170.4]
  assign RetimeWrapper_7_io_in = reset; // @[package.scala 94:16:@17169.4]
  assign RetimeWrapper_8_clock = clock; // @[:@17178.4]
  assign RetimeWrapper_8_reset = reset; // @[:@17179.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@17181.4]
  assign RetimeWrapper_8_io_in = _T_162 & _T_167; // @[package.scala 94:16:@17180.4]
  assign RetimeWrapper_9_clock = clock; // @[:@17186.4]
  assign RetimeWrapper_9_reset = reset; // @[:@17187.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@17189.4]
  assign RetimeWrapper_9_io_in = reset; // @[package.scala 94:16:@17188.4]
  assign RetimeWrapper_10_clock = clock; // @[:@17195.4]
  assign RetimeWrapper_10_reset = reset; // @[:@17196.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@17198.4]
  assign RetimeWrapper_10_io_in = _T_162 & _T_167; // @[package.scala 94:16:@17197.4]
  assign RetimeWrapper_11_clock = clock; // @[:@17203.4]
  assign RetimeWrapper_11_reset = reset; // @[:@17204.4]
  assign RetimeWrapper_11_io_flow = 1'h1; // @[package.scala 95:18:@17206.4]
  assign RetimeWrapper_11_io_in = reset; // @[package.scala 94:16:@17205.4]
  assign RetimeWrapper_12_clock = clock; // @[:@17214.4]
  assign RetimeWrapper_12_reset = reset; // @[:@17215.4]
  assign RetimeWrapper_12_io_flow = 1'h1; // @[package.scala 95:18:@17217.4]
  assign RetimeWrapper_12_io_in = _T_162 & _T_167; // @[package.scala 94:16:@17216.4]
  assign RetimeWrapper_13_clock = clock; // @[:@17222.4]
  assign RetimeWrapper_13_reset = reset; // @[:@17223.4]
  assign RetimeWrapper_13_io_flow = 1'h1; // @[package.scala 95:18:@17225.4]
  assign RetimeWrapper_13_io_in = reset; // @[package.scala 94:16:@17224.4]
  assign RetimeWrapper_14_clock = clock; // @[:@17231.4]
  assign RetimeWrapper_14_reset = reset; // @[:@17232.4]
  assign RetimeWrapper_14_io_flow = 1'h1; // @[package.scala 95:18:@17234.4]
  assign RetimeWrapper_14_io_in = _T_162 & _T_167; // @[package.scala 94:16:@17233.4]
  assign RetimeWrapper_15_clock = clock; // @[:@17239.4]
  assign RetimeWrapper_15_reset = reset; // @[:@17240.4]
  assign RetimeWrapper_15_io_flow = 1'h1; // @[package.scala 95:18:@17242.4]
  assign RetimeWrapper_15_io_in = reset; // @[package.scala 94:16:@17241.4]
  assign RetimeWrapper_16_clock = clock; // @[:@17250.4]
  assign RetimeWrapper_16_reset = reset; // @[:@17251.4]
  assign RetimeWrapper_16_io_flow = 1'h1; // @[package.scala 95:18:@17253.4]
  assign RetimeWrapper_16_io_in = _T_162 & _T_167; // @[package.scala 94:16:@17252.4]
  assign RetimeWrapper_17_clock = clock; // @[:@17258.4]
  assign RetimeWrapper_17_reset = reset; // @[:@17259.4]
  assign RetimeWrapper_17_io_flow = 1'h1; // @[package.scala 95:18:@17261.4]
  assign RetimeWrapper_17_io_in = reset; // @[package.scala 94:16:@17260.4]
  assign RetimeWrapper_18_clock = clock; // @[:@17267.4]
  assign RetimeWrapper_18_reset = reset; // @[:@17268.4]
  assign RetimeWrapper_18_io_flow = 1'h1; // @[package.scala 95:18:@17270.4]
  assign RetimeWrapper_18_io_in = _T_162 & _T_167; // @[package.scala 94:16:@17269.4]
  assign RetimeWrapper_19_clock = clock; // @[:@17275.4]
  assign RetimeWrapper_19_reset = reset; // @[:@17276.4]
  assign RetimeWrapper_19_io_flow = 1'h1; // @[package.scala 95:18:@17278.4]
  assign RetimeWrapper_19_io_in = reset; // @[package.scala 94:16:@17277.4]
  assign RetimeWrapper_20_clock = clock; // @[:@17286.4]
  assign RetimeWrapper_20_reset = reset; // @[:@17287.4]
  assign RetimeWrapper_20_io_flow = 1'h1; // @[package.scala 95:18:@17289.4]
  assign RetimeWrapper_20_io_in = _T_162 & _T_167; // @[package.scala 94:16:@17288.4]
  assign RetimeWrapper_21_clock = clock; // @[:@17294.4]
  assign RetimeWrapper_21_reset = reset; // @[:@17295.4]
  assign RetimeWrapper_21_io_flow = 1'h1; // @[package.scala 95:18:@17297.4]
  assign RetimeWrapper_21_io_in = reset; // @[package.scala 94:16:@17296.4]
  assign RetimeWrapper_22_clock = clock; // @[:@17303.4]
  assign RetimeWrapper_22_reset = reset; // @[:@17304.4]
  assign RetimeWrapper_22_io_flow = 1'h1; // @[package.scala 95:18:@17306.4]
  assign RetimeWrapper_22_io_in = _T_162 & _T_167; // @[package.scala 94:16:@17305.4]
  assign RetimeWrapper_23_clock = clock; // @[:@17311.4]
  assign RetimeWrapper_23_reset = reset; // @[:@17312.4]
  assign RetimeWrapper_23_io_flow = 1'h1; // @[package.scala 95:18:@17314.4]
  assign RetimeWrapper_23_io_in = reset; // @[package.scala 94:16:@17313.4]
  assign RetimeWrapper_24_clock = clock; // @[:@17322.4]
  assign RetimeWrapper_24_reset = reset; // @[:@17323.4]
  assign RetimeWrapper_24_io_flow = 1'h1; // @[package.scala 95:18:@17325.4]
  assign RetimeWrapper_24_io_in = _T_162 & _T_167; // @[package.scala 94:16:@17324.4]
  assign RetimeWrapper_25_clock = clock; // @[:@17330.4]
  assign RetimeWrapper_25_reset = reset; // @[:@17331.4]
  assign RetimeWrapper_25_io_flow = 1'h1; // @[package.scala 95:18:@17333.4]
  assign RetimeWrapper_25_io_in = reset; // @[package.scala 94:16:@17332.4]
  assign RetimeWrapper_26_clock = clock; // @[:@17339.4]
  assign RetimeWrapper_26_reset = reset; // @[:@17340.4]
  assign RetimeWrapper_26_io_flow = 1'h1; // @[package.scala 95:18:@17342.4]
  assign RetimeWrapper_26_io_in = _T_162 & _T_167; // @[package.scala 94:16:@17341.4]
  assign RetimeWrapper_27_clock = clock; // @[:@17347.4]
  assign RetimeWrapper_27_reset = reset; // @[:@17348.4]
  assign RetimeWrapper_27_io_flow = 1'h1; // @[package.scala 95:18:@17350.4]
  assign RetimeWrapper_27_io_in = reset; // @[package.scala 94:16:@17349.4]
  assign NBufCtr_clock = clock; // @[:@17388.4]
  assign NBufCtr_reset = reset; // @[:@17389.4]
  assign NBufCtr_io_input_countUp = 1'h0; // @[NBuffers.scala 43:24:@17396.4]
  assign NBufCtr_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 42:23:@17395.4]
  assign statesInR_0_clock = clock; // @[:@17399.4]
  assign statesInR_0_reset = reset; // @[:@17400.4]
  assign statesInR_0_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@17407.4]
  assign statesInR_0_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@17406.4]
  assign statesInR_1_clock = clock; // @[:@17410.4]
  assign statesInR_1_reset = reset; // @[:@17411.4]
  assign statesInR_1_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@17418.4]
  assign statesInR_1_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@17417.4]
  assign statesInR_2_clock = clock; // @[:@17421.4]
  assign statesInR_2_reset = reset; // @[:@17422.4]
  assign statesInR_2_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@17429.4]
  assign statesInR_2_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@17428.4]
  assign statesInR_3_clock = clock; // @[:@17432.4]
  assign statesInR_3_reset = reset; // @[:@17433.4]
  assign statesInR_3_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@17440.4]
  assign statesInR_3_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@17439.4]
  assign statesInR_4_clock = clock; // @[:@17443.4]
  assign statesInR_4_reset = reset; // @[:@17444.4]
  assign statesInR_4_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@17451.4]
  assign statesInR_4_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@17450.4]
  assign statesInR_5_clock = clock; // @[:@17454.4]
  assign statesInR_5_reset = reset; // @[:@17455.4]
  assign statesInR_5_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@17462.4]
  assign statesInR_5_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@17461.4]
  assign statesInR_6_clock = clock; // @[:@17465.4]
  assign statesInR_6_reset = reset; // @[:@17466.4]
  assign statesInR_6_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@17473.4]
  assign statesInR_6_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@17472.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_167 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_167 <= 1'h0;
    end else begin
      _T_167 <= _T_164;
    end
  end
endmodule
module FF_13( // @[:@17476.2]
  input         clock, // @[:@17477.4]
  input         reset, // @[:@17478.4]
  output [31:0] io_rPort_5_output_0, // @[:@17479.4]
  output [31:0] io_rPort_4_output_0, // @[:@17479.4]
  output [31:0] io_rPort_3_output_0, // @[:@17479.4]
  output [31:0] io_rPort_2_output_0, // @[:@17479.4]
  output [31:0] io_rPort_1_output_0, // @[:@17479.4]
  output [31:0] io_rPort_0_output_0, // @[:@17479.4]
  input  [31:0] io_wPort_0_data_0, // @[:@17479.4]
  input         io_wPort_0_reset, // @[:@17479.4]
  input         io_wPort_0_en_0 // @[:@17479.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@17519.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_198; // @[MemPrimitives.scala 325:32:@17521.4]
  wire [31:0] _T_199; // @[MemPrimitives.scala 325:12:@17522.4]
  assign _T_198 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@17521.4]
  assign _T_199 = io_wPort_0_reset ? 32'h0 : _T_198; // @[MemPrimitives.scala 325:12:@17522.4]
  assign io_rPort_5_output_0 = ff; // @[MemPrimitives.scala 326:34:@17529.4]
  assign io_rPort_4_output_0 = ff; // @[MemPrimitives.scala 326:34:@17528.4]
  assign io_rPort_3_output_0 = ff; // @[MemPrimitives.scala 326:34:@17527.4]
  assign io_rPort_2_output_0 = ff; // @[MemPrimitives.scala 326:34:@17526.4]
  assign io_rPort_1_output_0 = ff; // @[MemPrimitives.scala 326:34:@17525.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@17524.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module NBuf_2( // @[:@17861.2]
  input         clock, // @[:@17862.4]
  input         reset, // @[:@17863.4]
  output [31:0] io_rPort_5_output_0, // @[:@17864.4]
  output [31:0] io_rPort_4_output_0, // @[:@17864.4]
  output [31:0] io_rPort_3_output_0, // @[:@17864.4]
  output [31:0] io_rPort_2_output_0, // @[:@17864.4]
  output [31:0] io_rPort_1_output_0, // @[:@17864.4]
  output [31:0] io_rPort_0_output_0, // @[:@17864.4]
  input  [31:0] io_wPort_0_data_0, // @[:@17864.4]
  input         io_wPort_0_reset, // @[:@17864.4]
  input         io_wPort_0_en_0, // @[:@17864.4]
  input         io_sEn_0, // @[:@17864.4]
  input         io_sEn_1, // @[:@17864.4]
  input         io_sEn_2, // @[:@17864.4]
  input         io_sEn_3, // @[:@17864.4]
  input         io_sEn_4, // @[:@17864.4]
  input         io_sEn_5, // @[:@17864.4]
  input         io_sEn_6, // @[:@17864.4]
  input         io_sDone_0, // @[:@17864.4]
  input         io_sDone_1, // @[:@17864.4]
  input         io_sDone_2, // @[:@17864.4]
  input         io_sDone_3, // @[:@17864.4]
  input         io_sDone_4, // @[:@17864.4]
  input         io_sDone_5, // @[:@17864.4]
  input         io_sDone_6 // @[:@17864.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@17872.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@17872.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@17872.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@17872.4]
  wire  ctrl_io_sEn_2; // @[NBuffers.scala 83:20:@17872.4]
  wire  ctrl_io_sEn_3; // @[NBuffers.scala 83:20:@17872.4]
  wire  ctrl_io_sEn_4; // @[NBuffers.scala 83:20:@17872.4]
  wire  ctrl_io_sEn_5; // @[NBuffers.scala 83:20:@17872.4]
  wire  ctrl_io_sEn_6; // @[NBuffers.scala 83:20:@17872.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@17872.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@17872.4]
  wire  ctrl_io_sDone_2; // @[NBuffers.scala 83:20:@17872.4]
  wire  ctrl_io_sDone_3; // @[NBuffers.scala 83:20:@17872.4]
  wire  ctrl_io_sDone_4; // @[NBuffers.scala 83:20:@17872.4]
  wire  ctrl_io_sDone_5; // @[NBuffers.scala 83:20:@17872.4]
  wire  ctrl_io_sDone_6; // @[NBuffers.scala 83:20:@17872.4]
  wire [3:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@17872.4]
  wire [3:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@17872.4]
  wire [3:0] ctrl_io_statesInR_2; // @[NBuffers.scala 83:20:@17872.4]
  wire [3:0] ctrl_io_statesInR_3; // @[NBuffers.scala 83:20:@17872.4]
  wire [3:0] ctrl_io_statesInR_4; // @[NBuffers.scala 83:20:@17872.4]
  wire [3:0] ctrl_io_statesInR_5; // @[NBuffers.scala 83:20:@17872.4]
  wire [3:0] ctrl_io_statesInR_6; // @[NBuffers.scala 83:20:@17872.4]
  wire  FF_clock; // @[NBuffers.scala 146:23:@17889.4]
  wire  FF_reset; // @[NBuffers.scala 146:23:@17889.4]
  wire [31:0] FF_io_rPort_5_output_0; // @[NBuffers.scala 146:23:@17889.4]
  wire [31:0] FF_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@17889.4]
  wire [31:0] FF_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@17889.4]
  wire [31:0] FF_io_rPort_2_output_0; // @[NBuffers.scala 146:23:@17889.4]
  wire [31:0] FF_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@17889.4]
  wire [31:0] FF_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@17889.4]
  wire [31:0] FF_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@17889.4]
  wire  FF_io_wPort_0_reset; // @[NBuffers.scala 146:23:@17889.4]
  wire  FF_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@17889.4]
  wire  FF_1_clock; // @[NBuffers.scala 146:23:@17930.4]
  wire  FF_1_reset; // @[NBuffers.scala 146:23:@17930.4]
  wire [31:0] FF_1_io_rPort_5_output_0; // @[NBuffers.scala 146:23:@17930.4]
  wire [31:0] FF_1_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@17930.4]
  wire [31:0] FF_1_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@17930.4]
  wire [31:0] FF_1_io_rPort_2_output_0; // @[NBuffers.scala 146:23:@17930.4]
  wire [31:0] FF_1_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@17930.4]
  wire [31:0] FF_1_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@17930.4]
  wire [31:0] FF_1_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@17930.4]
  wire  FF_1_io_wPort_0_reset; // @[NBuffers.scala 146:23:@17930.4]
  wire  FF_1_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@17930.4]
  wire  FF_2_clock; // @[NBuffers.scala 146:23:@17971.4]
  wire  FF_2_reset; // @[NBuffers.scala 146:23:@17971.4]
  wire [31:0] FF_2_io_rPort_5_output_0; // @[NBuffers.scala 146:23:@17971.4]
  wire [31:0] FF_2_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@17971.4]
  wire [31:0] FF_2_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@17971.4]
  wire [31:0] FF_2_io_rPort_2_output_0; // @[NBuffers.scala 146:23:@17971.4]
  wire [31:0] FF_2_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@17971.4]
  wire [31:0] FF_2_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@17971.4]
  wire [31:0] FF_2_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@17971.4]
  wire  FF_2_io_wPort_0_reset; // @[NBuffers.scala 146:23:@17971.4]
  wire  FF_2_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@17971.4]
  wire  FF_3_clock; // @[NBuffers.scala 146:23:@18012.4]
  wire  FF_3_reset; // @[NBuffers.scala 146:23:@18012.4]
  wire [31:0] FF_3_io_rPort_5_output_0; // @[NBuffers.scala 146:23:@18012.4]
  wire [31:0] FF_3_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@18012.4]
  wire [31:0] FF_3_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@18012.4]
  wire [31:0] FF_3_io_rPort_2_output_0; // @[NBuffers.scala 146:23:@18012.4]
  wire [31:0] FF_3_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@18012.4]
  wire [31:0] FF_3_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@18012.4]
  wire [31:0] FF_3_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@18012.4]
  wire  FF_3_io_wPort_0_reset; // @[NBuffers.scala 146:23:@18012.4]
  wire  FF_3_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@18012.4]
  wire  FF_4_clock; // @[NBuffers.scala 146:23:@18053.4]
  wire  FF_4_reset; // @[NBuffers.scala 146:23:@18053.4]
  wire [31:0] FF_4_io_rPort_5_output_0; // @[NBuffers.scala 146:23:@18053.4]
  wire [31:0] FF_4_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@18053.4]
  wire [31:0] FF_4_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@18053.4]
  wire [31:0] FF_4_io_rPort_2_output_0; // @[NBuffers.scala 146:23:@18053.4]
  wire [31:0] FF_4_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@18053.4]
  wire [31:0] FF_4_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@18053.4]
  wire [31:0] FF_4_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@18053.4]
  wire  FF_4_io_wPort_0_reset; // @[NBuffers.scala 146:23:@18053.4]
  wire  FF_4_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@18053.4]
  wire  FF_5_clock; // @[NBuffers.scala 146:23:@18094.4]
  wire  FF_5_reset; // @[NBuffers.scala 146:23:@18094.4]
  wire [31:0] FF_5_io_rPort_5_output_0; // @[NBuffers.scala 146:23:@18094.4]
  wire [31:0] FF_5_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@18094.4]
  wire [31:0] FF_5_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@18094.4]
  wire [31:0] FF_5_io_rPort_2_output_0; // @[NBuffers.scala 146:23:@18094.4]
  wire [31:0] FF_5_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@18094.4]
  wire [31:0] FF_5_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@18094.4]
  wire [31:0] FF_5_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@18094.4]
  wire  FF_5_io_wPort_0_reset; // @[NBuffers.scala 146:23:@18094.4]
  wire  FF_5_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@18094.4]
  wire  FF_6_clock; // @[NBuffers.scala 146:23:@18135.4]
  wire  FF_6_reset; // @[NBuffers.scala 146:23:@18135.4]
  wire [31:0] FF_6_io_rPort_5_output_0; // @[NBuffers.scala 146:23:@18135.4]
  wire [31:0] FF_6_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@18135.4]
  wire [31:0] FF_6_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@18135.4]
  wire [31:0] FF_6_io_rPort_2_output_0; // @[NBuffers.scala 146:23:@18135.4]
  wire [31:0] FF_6_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@18135.4]
  wire [31:0] FF_6_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@18135.4]
  wire [31:0] FF_6_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@18135.4]
  wire  FF_6_io_wPort_0_reset; // @[NBuffers.scala 146:23:@18135.4]
  wire  FF_6_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@18135.4]
  wire  _T_236; // @[NBuffers.scala 153:105:@18183.4]
  wire  _T_240; // @[NBuffers.scala 157:92:@18193.4]
  wire  _T_243; // @[NBuffers.scala 157:92:@18199.4]
  wire  _T_246; // @[NBuffers.scala 157:92:@18205.4]
  wire  _T_249; // @[NBuffers.scala 157:92:@18211.4]
  wire  _T_252; // @[NBuffers.scala 157:92:@18217.4]
  wire  _T_255; // @[NBuffers.scala 157:92:@18223.4]
  wire  _T_258; // @[NBuffers.scala 153:105:@18229.4]
  wire  _T_262; // @[NBuffers.scala 157:92:@18239.4]
  wire  _T_265; // @[NBuffers.scala 157:92:@18245.4]
  wire  _T_268; // @[NBuffers.scala 157:92:@18251.4]
  wire  _T_271; // @[NBuffers.scala 157:92:@18257.4]
  wire  _T_274; // @[NBuffers.scala 157:92:@18263.4]
  wire  _T_277; // @[NBuffers.scala 157:92:@18269.4]
  wire  _T_280; // @[NBuffers.scala 153:105:@18275.4]
  wire  _T_284; // @[NBuffers.scala 157:92:@18285.4]
  wire  _T_287; // @[NBuffers.scala 157:92:@18291.4]
  wire  _T_290; // @[NBuffers.scala 157:92:@18297.4]
  wire  _T_293; // @[NBuffers.scala 157:92:@18303.4]
  wire  _T_296; // @[NBuffers.scala 157:92:@18309.4]
  wire  _T_299; // @[NBuffers.scala 157:92:@18315.4]
  wire  _T_302; // @[NBuffers.scala 153:105:@18321.4]
  wire  _T_306; // @[NBuffers.scala 157:92:@18331.4]
  wire  _T_309; // @[NBuffers.scala 157:92:@18337.4]
  wire  _T_312; // @[NBuffers.scala 157:92:@18343.4]
  wire  _T_315; // @[NBuffers.scala 157:92:@18349.4]
  wire  _T_318; // @[NBuffers.scala 157:92:@18355.4]
  wire  _T_321; // @[NBuffers.scala 157:92:@18361.4]
  wire  _T_324; // @[NBuffers.scala 153:105:@18367.4]
  wire  _T_328; // @[NBuffers.scala 157:92:@18377.4]
  wire  _T_331; // @[NBuffers.scala 157:92:@18383.4]
  wire  _T_334; // @[NBuffers.scala 157:92:@18389.4]
  wire  _T_337; // @[NBuffers.scala 157:92:@18395.4]
  wire  _T_340; // @[NBuffers.scala 157:92:@18401.4]
  wire  _T_343; // @[NBuffers.scala 157:92:@18407.4]
  wire  _T_346; // @[NBuffers.scala 153:105:@18413.4]
  wire  _T_350; // @[NBuffers.scala 157:92:@18423.4]
  wire  _T_353; // @[NBuffers.scala 157:92:@18429.4]
  wire  _T_356; // @[NBuffers.scala 157:92:@18435.4]
  wire  _T_359; // @[NBuffers.scala 157:92:@18441.4]
  wire  _T_362; // @[NBuffers.scala 157:92:@18447.4]
  wire  _T_365; // @[NBuffers.scala 157:92:@18453.4]
  wire  _T_368; // @[NBuffers.scala 153:105:@18459.4]
  wire  _T_372; // @[NBuffers.scala 157:92:@18469.4]
  wire  _T_375; // @[NBuffers.scala 157:92:@18475.4]
  wire  _T_378; // @[NBuffers.scala 157:92:@18481.4]
  wire  _T_381; // @[NBuffers.scala 157:92:@18487.4]
  wire  _T_384; // @[NBuffers.scala 157:92:@18493.4]
  wire  _T_387; // @[NBuffers.scala 157:92:@18499.4]
  wire [31:0] _T_405; // @[Mux.scala 19:72:@18512.4]
  wire [31:0] _T_407; // @[Mux.scala 19:72:@18513.4]
  wire [31:0] _T_409; // @[Mux.scala 19:72:@18514.4]
  wire [31:0] _T_411; // @[Mux.scala 19:72:@18515.4]
  wire [31:0] _T_413; // @[Mux.scala 19:72:@18516.4]
  wire [31:0] _T_415; // @[Mux.scala 19:72:@18517.4]
  wire [31:0] _T_417; // @[Mux.scala 19:72:@18518.4]
  wire [31:0] _T_418; // @[Mux.scala 19:72:@18519.4]
  wire [31:0] _T_419; // @[Mux.scala 19:72:@18520.4]
  wire [31:0] _T_420; // @[Mux.scala 19:72:@18521.4]
  wire [31:0] _T_421; // @[Mux.scala 19:72:@18522.4]
  wire [31:0] _T_422; // @[Mux.scala 19:72:@18523.4]
  wire [31:0] _T_442; // @[Mux.scala 19:72:@18535.4]
  wire [31:0] _T_444; // @[Mux.scala 19:72:@18536.4]
  wire [31:0] _T_446; // @[Mux.scala 19:72:@18537.4]
  wire [31:0] _T_448; // @[Mux.scala 19:72:@18538.4]
  wire [31:0] _T_450; // @[Mux.scala 19:72:@18539.4]
  wire [31:0] _T_452; // @[Mux.scala 19:72:@18540.4]
  wire [31:0] _T_454; // @[Mux.scala 19:72:@18541.4]
  wire [31:0] _T_455; // @[Mux.scala 19:72:@18542.4]
  wire [31:0] _T_456; // @[Mux.scala 19:72:@18543.4]
  wire [31:0] _T_457; // @[Mux.scala 19:72:@18544.4]
  wire [31:0] _T_458; // @[Mux.scala 19:72:@18545.4]
  wire [31:0] _T_459; // @[Mux.scala 19:72:@18546.4]
  wire [31:0] _T_479; // @[Mux.scala 19:72:@18558.4]
  wire [31:0] _T_481; // @[Mux.scala 19:72:@18559.4]
  wire [31:0] _T_483; // @[Mux.scala 19:72:@18560.4]
  wire [31:0] _T_485; // @[Mux.scala 19:72:@18561.4]
  wire [31:0] _T_487; // @[Mux.scala 19:72:@18562.4]
  wire [31:0] _T_489; // @[Mux.scala 19:72:@18563.4]
  wire [31:0] _T_491; // @[Mux.scala 19:72:@18564.4]
  wire [31:0] _T_492; // @[Mux.scala 19:72:@18565.4]
  wire [31:0] _T_493; // @[Mux.scala 19:72:@18566.4]
  wire [31:0] _T_494; // @[Mux.scala 19:72:@18567.4]
  wire [31:0] _T_495; // @[Mux.scala 19:72:@18568.4]
  wire [31:0] _T_496; // @[Mux.scala 19:72:@18569.4]
  wire [31:0] _T_516; // @[Mux.scala 19:72:@18581.4]
  wire [31:0] _T_518; // @[Mux.scala 19:72:@18582.4]
  wire [31:0] _T_520; // @[Mux.scala 19:72:@18583.4]
  wire [31:0] _T_522; // @[Mux.scala 19:72:@18584.4]
  wire [31:0] _T_524; // @[Mux.scala 19:72:@18585.4]
  wire [31:0] _T_526; // @[Mux.scala 19:72:@18586.4]
  wire [31:0] _T_528; // @[Mux.scala 19:72:@18587.4]
  wire [31:0] _T_529; // @[Mux.scala 19:72:@18588.4]
  wire [31:0] _T_530; // @[Mux.scala 19:72:@18589.4]
  wire [31:0] _T_531; // @[Mux.scala 19:72:@18590.4]
  wire [31:0] _T_532; // @[Mux.scala 19:72:@18591.4]
  wire [31:0] _T_533; // @[Mux.scala 19:72:@18592.4]
  wire [31:0] _T_553; // @[Mux.scala 19:72:@18604.4]
  wire [31:0] _T_555; // @[Mux.scala 19:72:@18605.4]
  wire [31:0] _T_557; // @[Mux.scala 19:72:@18606.4]
  wire [31:0] _T_559; // @[Mux.scala 19:72:@18607.4]
  wire [31:0] _T_561; // @[Mux.scala 19:72:@18608.4]
  wire [31:0] _T_563; // @[Mux.scala 19:72:@18609.4]
  wire [31:0] _T_565; // @[Mux.scala 19:72:@18610.4]
  wire [31:0] _T_566; // @[Mux.scala 19:72:@18611.4]
  wire [31:0] _T_567; // @[Mux.scala 19:72:@18612.4]
  wire [31:0] _T_568; // @[Mux.scala 19:72:@18613.4]
  wire [31:0] _T_569; // @[Mux.scala 19:72:@18614.4]
  wire [31:0] _T_570; // @[Mux.scala 19:72:@18615.4]
  wire [31:0] _T_590; // @[Mux.scala 19:72:@18627.4]
  wire [31:0] _T_592; // @[Mux.scala 19:72:@18628.4]
  wire [31:0] _T_594; // @[Mux.scala 19:72:@18629.4]
  wire [31:0] _T_596; // @[Mux.scala 19:72:@18630.4]
  wire [31:0] _T_598; // @[Mux.scala 19:72:@18631.4]
  wire [31:0] _T_600; // @[Mux.scala 19:72:@18632.4]
  wire [31:0] _T_602; // @[Mux.scala 19:72:@18633.4]
  wire [31:0] _T_603; // @[Mux.scala 19:72:@18634.4]
  wire [31:0] _T_604; // @[Mux.scala 19:72:@18635.4]
  wire [31:0] _T_605; // @[Mux.scala 19:72:@18636.4]
  wire [31:0] _T_606; // @[Mux.scala 19:72:@18637.4]
  wire [31:0] _T_607; // @[Mux.scala 19:72:@18638.4]
  NBufController_3 ctrl ( // @[NBuffers.scala 83:20:@17872.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sEn_2(ctrl_io_sEn_2),
    .io_sEn_3(ctrl_io_sEn_3),
    .io_sEn_4(ctrl_io_sEn_4),
    .io_sEn_5(ctrl_io_sEn_5),
    .io_sEn_6(ctrl_io_sEn_6),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_sDone_2(ctrl_io_sDone_2),
    .io_sDone_3(ctrl_io_sDone_3),
    .io_sDone_4(ctrl_io_sDone_4),
    .io_sDone_5(ctrl_io_sDone_5),
    .io_sDone_6(ctrl_io_sDone_6),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1),
    .io_statesInR_2(ctrl_io_statesInR_2),
    .io_statesInR_3(ctrl_io_statesInR_3),
    .io_statesInR_4(ctrl_io_statesInR_4),
    .io_statesInR_5(ctrl_io_statesInR_5),
    .io_statesInR_6(ctrl_io_statesInR_6)
  );
  FF_13 FF ( // @[NBuffers.scala 146:23:@17889.4]
    .clock(FF_clock),
    .reset(FF_reset),
    .io_rPort_5_output_0(FF_io_rPort_5_output_0),
    .io_rPort_4_output_0(FF_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_io_rPort_3_output_0),
    .io_rPort_2_output_0(FF_io_rPort_2_output_0),
    .io_rPort_1_output_0(FF_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_io_wPort_0_en_0)
  );
  FF_13 FF_1 ( // @[NBuffers.scala 146:23:@17930.4]
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_rPort_5_output_0(FF_1_io_rPort_5_output_0),
    .io_rPort_4_output_0(FF_1_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_1_io_rPort_3_output_0),
    .io_rPort_2_output_0(FF_1_io_rPort_2_output_0),
    .io_rPort_1_output_0(FF_1_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_1_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_1_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_1_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_1_io_wPort_0_en_0)
  );
  FF_13 FF_2 ( // @[NBuffers.scala 146:23:@17971.4]
    .clock(FF_2_clock),
    .reset(FF_2_reset),
    .io_rPort_5_output_0(FF_2_io_rPort_5_output_0),
    .io_rPort_4_output_0(FF_2_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_2_io_rPort_3_output_0),
    .io_rPort_2_output_0(FF_2_io_rPort_2_output_0),
    .io_rPort_1_output_0(FF_2_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_2_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_2_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_2_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_2_io_wPort_0_en_0)
  );
  FF_13 FF_3 ( // @[NBuffers.scala 146:23:@18012.4]
    .clock(FF_3_clock),
    .reset(FF_3_reset),
    .io_rPort_5_output_0(FF_3_io_rPort_5_output_0),
    .io_rPort_4_output_0(FF_3_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_3_io_rPort_3_output_0),
    .io_rPort_2_output_0(FF_3_io_rPort_2_output_0),
    .io_rPort_1_output_0(FF_3_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_3_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_3_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_3_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_3_io_wPort_0_en_0)
  );
  FF_13 FF_4 ( // @[NBuffers.scala 146:23:@18053.4]
    .clock(FF_4_clock),
    .reset(FF_4_reset),
    .io_rPort_5_output_0(FF_4_io_rPort_5_output_0),
    .io_rPort_4_output_0(FF_4_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_4_io_rPort_3_output_0),
    .io_rPort_2_output_0(FF_4_io_rPort_2_output_0),
    .io_rPort_1_output_0(FF_4_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_4_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_4_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_4_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_4_io_wPort_0_en_0)
  );
  FF_13 FF_5 ( // @[NBuffers.scala 146:23:@18094.4]
    .clock(FF_5_clock),
    .reset(FF_5_reset),
    .io_rPort_5_output_0(FF_5_io_rPort_5_output_0),
    .io_rPort_4_output_0(FF_5_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_5_io_rPort_3_output_0),
    .io_rPort_2_output_0(FF_5_io_rPort_2_output_0),
    .io_rPort_1_output_0(FF_5_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_5_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_5_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_5_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_5_io_wPort_0_en_0)
  );
  FF_13 FF_6 ( // @[NBuffers.scala 146:23:@18135.4]
    .clock(FF_6_clock),
    .reset(FF_6_reset),
    .io_rPort_5_output_0(FF_6_io_rPort_5_output_0),
    .io_rPort_4_output_0(FF_6_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_6_io_rPort_3_output_0),
    .io_rPort_2_output_0(FF_6_io_rPort_2_output_0),
    .io_rPort_1_output_0(FF_6_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_6_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_6_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_6_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_6_io_wPort_0_en_0)
  );
  assign _T_236 = ctrl_io_statesInW_0 == 4'h0; // @[NBuffers.scala 153:105:@18183.4]
  assign _T_240 = ctrl_io_statesInR_1 == 4'h0; // @[NBuffers.scala 157:92:@18193.4]
  assign _T_243 = ctrl_io_statesInR_2 == 4'h0; // @[NBuffers.scala 157:92:@18199.4]
  assign _T_246 = ctrl_io_statesInR_3 == 4'h0; // @[NBuffers.scala 157:92:@18205.4]
  assign _T_249 = ctrl_io_statesInR_4 == 4'h0; // @[NBuffers.scala 157:92:@18211.4]
  assign _T_252 = ctrl_io_statesInR_5 == 4'h0; // @[NBuffers.scala 157:92:@18217.4]
  assign _T_255 = ctrl_io_statesInR_6 == 4'h0; // @[NBuffers.scala 157:92:@18223.4]
  assign _T_258 = ctrl_io_statesInW_0 == 4'h1; // @[NBuffers.scala 153:105:@18229.4]
  assign _T_262 = ctrl_io_statesInR_1 == 4'h1; // @[NBuffers.scala 157:92:@18239.4]
  assign _T_265 = ctrl_io_statesInR_2 == 4'h1; // @[NBuffers.scala 157:92:@18245.4]
  assign _T_268 = ctrl_io_statesInR_3 == 4'h1; // @[NBuffers.scala 157:92:@18251.4]
  assign _T_271 = ctrl_io_statesInR_4 == 4'h1; // @[NBuffers.scala 157:92:@18257.4]
  assign _T_274 = ctrl_io_statesInR_5 == 4'h1; // @[NBuffers.scala 157:92:@18263.4]
  assign _T_277 = ctrl_io_statesInR_6 == 4'h1; // @[NBuffers.scala 157:92:@18269.4]
  assign _T_280 = ctrl_io_statesInW_0 == 4'h2; // @[NBuffers.scala 153:105:@18275.4]
  assign _T_284 = ctrl_io_statesInR_1 == 4'h2; // @[NBuffers.scala 157:92:@18285.4]
  assign _T_287 = ctrl_io_statesInR_2 == 4'h2; // @[NBuffers.scala 157:92:@18291.4]
  assign _T_290 = ctrl_io_statesInR_3 == 4'h2; // @[NBuffers.scala 157:92:@18297.4]
  assign _T_293 = ctrl_io_statesInR_4 == 4'h2; // @[NBuffers.scala 157:92:@18303.4]
  assign _T_296 = ctrl_io_statesInR_5 == 4'h2; // @[NBuffers.scala 157:92:@18309.4]
  assign _T_299 = ctrl_io_statesInR_6 == 4'h2; // @[NBuffers.scala 157:92:@18315.4]
  assign _T_302 = ctrl_io_statesInW_0 == 4'h3; // @[NBuffers.scala 153:105:@18321.4]
  assign _T_306 = ctrl_io_statesInR_1 == 4'h3; // @[NBuffers.scala 157:92:@18331.4]
  assign _T_309 = ctrl_io_statesInR_2 == 4'h3; // @[NBuffers.scala 157:92:@18337.4]
  assign _T_312 = ctrl_io_statesInR_3 == 4'h3; // @[NBuffers.scala 157:92:@18343.4]
  assign _T_315 = ctrl_io_statesInR_4 == 4'h3; // @[NBuffers.scala 157:92:@18349.4]
  assign _T_318 = ctrl_io_statesInR_5 == 4'h3; // @[NBuffers.scala 157:92:@18355.4]
  assign _T_321 = ctrl_io_statesInR_6 == 4'h3; // @[NBuffers.scala 157:92:@18361.4]
  assign _T_324 = ctrl_io_statesInW_0 == 4'h4; // @[NBuffers.scala 153:105:@18367.4]
  assign _T_328 = ctrl_io_statesInR_1 == 4'h4; // @[NBuffers.scala 157:92:@18377.4]
  assign _T_331 = ctrl_io_statesInR_2 == 4'h4; // @[NBuffers.scala 157:92:@18383.4]
  assign _T_334 = ctrl_io_statesInR_3 == 4'h4; // @[NBuffers.scala 157:92:@18389.4]
  assign _T_337 = ctrl_io_statesInR_4 == 4'h4; // @[NBuffers.scala 157:92:@18395.4]
  assign _T_340 = ctrl_io_statesInR_5 == 4'h4; // @[NBuffers.scala 157:92:@18401.4]
  assign _T_343 = ctrl_io_statesInR_6 == 4'h4; // @[NBuffers.scala 157:92:@18407.4]
  assign _T_346 = ctrl_io_statesInW_0 == 4'h5; // @[NBuffers.scala 153:105:@18413.4]
  assign _T_350 = ctrl_io_statesInR_1 == 4'h5; // @[NBuffers.scala 157:92:@18423.4]
  assign _T_353 = ctrl_io_statesInR_2 == 4'h5; // @[NBuffers.scala 157:92:@18429.4]
  assign _T_356 = ctrl_io_statesInR_3 == 4'h5; // @[NBuffers.scala 157:92:@18435.4]
  assign _T_359 = ctrl_io_statesInR_4 == 4'h5; // @[NBuffers.scala 157:92:@18441.4]
  assign _T_362 = ctrl_io_statesInR_5 == 4'h5; // @[NBuffers.scala 157:92:@18447.4]
  assign _T_365 = ctrl_io_statesInR_6 == 4'h5; // @[NBuffers.scala 157:92:@18453.4]
  assign _T_368 = ctrl_io_statesInW_0 == 4'h6; // @[NBuffers.scala 153:105:@18459.4]
  assign _T_372 = ctrl_io_statesInR_1 == 4'h6; // @[NBuffers.scala 157:92:@18469.4]
  assign _T_375 = ctrl_io_statesInR_2 == 4'h6; // @[NBuffers.scala 157:92:@18475.4]
  assign _T_378 = ctrl_io_statesInR_3 == 4'h6; // @[NBuffers.scala 157:92:@18481.4]
  assign _T_381 = ctrl_io_statesInR_4 == 4'h6; // @[NBuffers.scala 157:92:@18487.4]
  assign _T_384 = ctrl_io_statesInR_5 == 4'h6; // @[NBuffers.scala 157:92:@18493.4]
  assign _T_387 = ctrl_io_statesInR_6 == 4'h6; // @[NBuffers.scala 157:92:@18499.4]
  assign _T_405 = _T_240 ? FF_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@18512.4]
  assign _T_407 = _T_262 ? FF_1_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@18513.4]
  assign _T_409 = _T_284 ? FF_2_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@18514.4]
  assign _T_411 = _T_306 ? FF_3_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@18515.4]
  assign _T_413 = _T_328 ? FF_4_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@18516.4]
  assign _T_415 = _T_350 ? FF_5_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@18517.4]
  assign _T_417 = _T_372 ? FF_6_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@18518.4]
  assign _T_418 = _T_405 | _T_407; // @[Mux.scala 19:72:@18519.4]
  assign _T_419 = _T_418 | _T_409; // @[Mux.scala 19:72:@18520.4]
  assign _T_420 = _T_419 | _T_411; // @[Mux.scala 19:72:@18521.4]
  assign _T_421 = _T_420 | _T_413; // @[Mux.scala 19:72:@18522.4]
  assign _T_422 = _T_421 | _T_415; // @[Mux.scala 19:72:@18523.4]
  assign _T_442 = _T_243 ? FF_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@18535.4]
  assign _T_444 = _T_265 ? FF_1_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@18536.4]
  assign _T_446 = _T_287 ? FF_2_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@18537.4]
  assign _T_448 = _T_309 ? FF_3_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@18538.4]
  assign _T_450 = _T_331 ? FF_4_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@18539.4]
  assign _T_452 = _T_353 ? FF_5_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@18540.4]
  assign _T_454 = _T_375 ? FF_6_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@18541.4]
  assign _T_455 = _T_442 | _T_444; // @[Mux.scala 19:72:@18542.4]
  assign _T_456 = _T_455 | _T_446; // @[Mux.scala 19:72:@18543.4]
  assign _T_457 = _T_456 | _T_448; // @[Mux.scala 19:72:@18544.4]
  assign _T_458 = _T_457 | _T_450; // @[Mux.scala 19:72:@18545.4]
  assign _T_459 = _T_458 | _T_452; // @[Mux.scala 19:72:@18546.4]
  assign _T_479 = _T_246 ? FF_io_rPort_2_output_0 : 32'h0; // @[Mux.scala 19:72:@18558.4]
  assign _T_481 = _T_268 ? FF_1_io_rPort_2_output_0 : 32'h0; // @[Mux.scala 19:72:@18559.4]
  assign _T_483 = _T_290 ? FF_2_io_rPort_2_output_0 : 32'h0; // @[Mux.scala 19:72:@18560.4]
  assign _T_485 = _T_312 ? FF_3_io_rPort_2_output_0 : 32'h0; // @[Mux.scala 19:72:@18561.4]
  assign _T_487 = _T_334 ? FF_4_io_rPort_2_output_0 : 32'h0; // @[Mux.scala 19:72:@18562.4]
  assign _T_489 = _T_356 ? FF_5_io_rPort_2_output_0 : 32'h0; // @[Mux.scala 19:72:@18563.4]
  assign _T_491 = _T_378 ? FF_6_io_rPort_2_output_0 : 32'h0; // @[Mux.scala 19:72:@18564.4]
  assign _T_492 = _T_479 | _T_481; // @[Mux.scala 19:72:@18565.4]
  assign _T_493 = _T_492 | _T_483; // @[Mux.scala 19:72:@18566.4]
  assign _T_494 = _T_493 | _T_485; // @[Mux.scala 19:72:@18567.4]
  assign _T_495 = _T_494 | _T_487; // @[Mux.scala 19:72:@18568.4]
  assign _T_496 = _T_495 | _T_489; // @[Mux.scala 19:72:@18569.4]
  assign _T_516 = _T_249 ? FF_io_rPort_3_output_0 : 32'h0; // @[Mux.scala 19:72:@18581.4]
  assign _T_518 = _T_271 ? FF_1_io_rPort_3_output_0 : 32'h0; // @[Mux.scala 19:72:@18582.4]
  assign _T_520 = _T_293 ? FF_2_io_rPort_3_output_0 : 32'h0; // @[Mux.scala 19:72:@18583.4]
  assign _T_522 = _T_315 ? FF_3_io_rPort_3_output_0 : 32'h0; // @[Mux.scala 19:72:@18584.4]
  assign _T_524 = _T_337 ? FF_4_io_rPort_3_output_0 : 32'h0; // @[Mux.scala 19:72:@18585.4]
  assign _T_526 = _T_359 ? FF_5_io_rPort_3_output_0 : 32'h0; // @[Mux.scala 19:72:@18586.4]
  assign _T_528 = _T_381 ? FF_6_io_rPort_3_output_0 : 32'h0; // @[Mux.scala 19:72:@18587.4]
  assign _T_529 = _T_516 | _T_518; // @[Mux.scala 19:72:@18588.4]
  assign _T_530 = _T_529 | _T_520; // @[Mux.scala 19:72:@18589.4]
  assign _T_531 = _T_530 | _T_522; // @[Mux.scala 19:72:@18590.4]
  assign _T_532 = _T_531 | _T_524; // @[Mux.scala 19:72:@18591.4]
  assign _T_533 = _T_532 | _T_526; // @[Mux.scala 19:72:@18592.4]
  assign _T_553 = _T_252 ? FF_io_rPort_4_output_0 : 32'h0; // @[Mux.scala 19:72:@18604.4]
  assign _T_555 = _T_274 ? FF_1_io_rPort_4_output_0 : 32'h0; // @[Mux.scala 19:72:@18605.4]
  assign _T_557 = _T_296 ? FF_2_io_rPort_4_output_0 : 32'h0; // @[Mux.scala 19:72:@18606.4]
  assign _T_559 = _T_318 ? FF_3_io_rPort_4_output_0 : 32'h0; // @[Mux.scala 19:72:@18607.4]
  assign _T_561 = _T_340 ? FF_4_io_rPort_4_output_0 : 32'h0; // @[Mux.scala 19:72:@18608.4]
  assign _T_563 = _T_362 ? FF_5_io_rPort_4_output_0 : 32'h0; // @[Mux.scala 19:72:@18609.4]
  assign _T_565 = _T_384 ? FF_6_io_rPort_4_output_0 : 32'h0; // @[Mux.scala 19:72:@18610.4]
  assign _T_566 = _T_553 | _T_555; // @[Mux.scala 19:72:@18611.4]
  assign _T_567 = _T_566 | _T_557; // @[Mux.scala 19:72:@18612.4]
  assign _T_568 = _T_567 | _T_559; // @[Mux.scala 19:72:@18613.4]
  assign _T_569 = _T_568 | _T_561; // @[Mux.scala 19:72:@18614.4]
  assign _T_570 = _T_569 | _T_563; // @[Mux.scala 19:72:@18615.4]
  assign _T_590 = _T_255 ? FF_io_rPort_5_output_0 : 32'h0; // @[Mux.scala 19:72:@18627.4]
  assign _T_592 = _T_277 ? FF_1_io_rPort_5_output_0 : 32'h0; // @[Mux.scala 19:72:@18628.4]
  assign _T_594 = _T_299 ? FF_2_io_rPort_5_output_0 : 32'h0; // @[Mux.scala 19:72:@18629.4]
  assign _T_596 = _T_321 ? FF_3_io_rPort_5_output_0 : 32'h0; // @[Mux.scala 19:72:@18630.4]
  assign _T_598 = _T_343 ? FF_4_io_rPort_5_output_0 : 32'h0; // @[Mux.scala 19:72:@18631.4]
  assign _T_600 = _T_365 ? FF_5_io_rPort_5_output_0 : 32'h0; // @[Mux.scala 19:72:@18632.4]
  assign _T_602 = _T_387 ? FF_6_io_rPort_5_output_0 : 32'h0; // @[Mux.scala 19:72:@18633.4]
  assign _T_603 = _T_590 | _T_592; // @[Mux.scala 19:72:@18634.4]
  assign _T_604 = _T_603 | _T_594; // @[Mux.scala 19:72:@18635.4]
  assign _T_605 = _T_604 | _T_596; // @[Mux.scala 19:72:@18636.4]
  assign _T_606 = _T_605 | _T_598; // @[Mux.scala 19:72:@18637.4]
  assign _T_607 = _T_606 | _T_600; // @[Mux.scala 19:72:@18638.4]
  assign io_rPort_5_output_0 = _T_607 | _T_602; // @[NBuffers.scala 163:66:@18642.4]
  assign io_rPort_4_output_0 = _T_570 | _T_565; // @[NBuffers.scala 163:66:@18619.4]
  assign io_rPort_3_output_0 = _T_533 | _T_528; // @[NBuffers.scala 163:66:@18596.4]
  assign io_rPort_2_output_0 = _T_496 | _T_491; // @[NBuffers.scala 163:66:@18573.4]
  assign io_rPort_1_output_0 = _T_459 | _T_454; // @[NBuffers.scala 163:66:@18550.4]
  assign io_rPort_0_output_0 = _T_422 | _T_417; // @[NBuffers.scala 163:66:@18527.4]
  assign ctrl_clock = clock; // @[:@17873.4]
  assign ctrl_reset = reset; // @[:@17874.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@17875.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@17877.4]
  assign ctrl_io_sEn_2 = io_sEn_2; // @[NBuffers.scala 85:20:@17879.4]
  assign ctrl_io_sEn_3 = io_sEn_3; // @[NBuffers.scala 85:20:@17881.4]
  assign ctrl_io_sEn_4 = io_sEn_4; // @[NBuffers.scala 85:20:@17883.4]
  assign ctrl_io_sEn_5 = io_sEn_5; // @[NBuffers.scala 85:20:@17885.4]
  assign ctrl_io_sEn_6 = io_sEn_6; // @[NBuffers.scala 85:20:@17887.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@17876.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@17878.4]
  assign ctrl_io_sDone_2 = io_sDone_2; // @[NBuffers.scala 86:22:@17880.4]
  assign ctrl_io_sDone_3 = io_sDone_3; // @[NBuffers.scala 86:22:@17882.4]
  assign ctrl_io_sDone_4 = io_sDone_4; // @[NBuffers.scala 86:22:@17884.4]
  assign ctrl_io_sDone_5 = io_sDone_5; // @[NBuffers.scala 86:22:@17886.4]
  assign ctrl_io_sDone_6 = io_sDone_6; // @[NBuffers.scala 86:22:@17888.4]
  assign FF_clock = clock; // @[:@17890.4]
  assign FF_reset = reset; // @[:@17891.4]
  assign FF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@18186.4]
  assign FF_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@18187.4]
  assign FF_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_236; // @[MemPrimitives.scala 37:29:@18192.4]
  assign FF_1_clock = clock; // @[:@17931.4]
  assign FF_1_reset = reset; // @[:@17932.4]
  assign FF_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@18232.4]
  assign FF_1_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@18233.4]
  assign FF_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_258; // @[MemPrimitives.scala 37:29:@18238.4]
  assign FF_2_clock = clock; // @[:@17972.4]
  assign FF_2_reset = reset; // @[:@17973.4]
  assign FF_2_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@18278.4]
  assign FF_2_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@18279.4]
  assign FF_2_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_280; // @[MemPrimitives.scala 37:29:@18284.4]
  assign FF_3_clock = clock; // @[:@18013.4]
  assign FF_3_reset = reset; // @[:@18014.4]
  assign FF_3_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@18324.4]
  assign FF_3_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@18325.4]
  assign FF_3_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_302; // @[MemPrimitives.scala 37:29:@18330.4]
  assign FF_4_clock = clock; // @[:@18054.4]
  assign FF_4_reset = reset; // @[:@18055.4]
  assign FF_4_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@18370.4]
  assign FF_4_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@18371.4]
  assign FF_4_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_324; // @[MemPrimitives.scala 37:29:@18376.4]
  assign FF_5_clock = clock; // @[:@18095.4]
  assign FF_5_reset = reset; // @[:@18096.4]
  assign FF_5_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@18416.4]
  assign FF_5_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@18417.4]
  assign FF_5_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_346; // @[MemPrimitives.scala 37:29:@18422.4]
  assign FF_6_clock = clock; // @[:@18136.4]
  assign FF_6_reset = reset; // @[:@18137.4]
  assign FF_6_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@18462.4]
  assign FF_6_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@18463.4]
  assign FF_6_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_368; // @[MemPrimitives.scala 37:29:@18468.4]
endmodule
module b550_chain( // @[:@18644.2]
  input         clock, // @[:@18645.4]
  input         reset, // @[:@18646.4]
  output [31:0] io_rPort_5_output_0, // @[:@18647.4]
  output [31:0] io_rPort_4_output_0, // @[:@18647.4]
  output [31:0] io_rPort_3_output_0, // @[:@18647.4]
  output [31:0] io_rPort_2_output_0, // @[:@18647.4]
  output [31:0] io_rPort_1_output_0, // @[:@18647.4]
  output [31:0] io_rPort_0_output_0, // @[:@18647.4]
  input  [31:0] io_wPort_0_data_0, // @[:@18647.4]
  input         io_wPort_0_reset, // @[:@18647.4]
  input         io_wPort_0_en_0, // @[:@18647.4]
  input         io_sEn_0, // @[:@18647.4]
  input         io_sEn_1, // @[:@18647.4]
  input         io_sEn_2, // @[:@18647.4]
  input         io_sEn_3, // @[:@18647.4]
  input         io_sEn_4, // @[:@18647.4]
  input         io_sEn_5, // @[:@18647.4]
  input         io_sEn_6, // @[:@18647.4]
  input         io_sDone_0, // @[:@18647.4]
  input         io_sDone_1, // @[:@18647.4]
  input         io_sDone_2, // @[:@18647.4]
  input         io_sDone_3, // @[:@18647.4]
  input         io_sDone_4, // @[:@18647.4]
  input         io_sDone_5, // @[:@18647.4]
  input         io_sDone_6 // @[:@18647.4]
);
  wire  nbufFF_clock; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_reset; // @[NBuffers.scala 298:22:@18655.4]
  wire [31:0] nbufFF_io_rPort_5_output_0; // @[NBuffers.scala 298:22:@18655.4]
  wire [31:0] nbufFF_io_rPort_4_output_0; // @[NBuffers.scala 298:22:@18655.4]
  wire [31:0] nbufFF_io_rPort_3_output_0; // @[NBuffers.scala 298:22:@18655.4]
  wire [31:0] nbufFF_io_rPort_2_output_0; // @[NBuffers.scala 298:22:@18655.4]
  wire [31:0] nbufFF_io_rPort_1_output_0; // @[NBuffers.scala 298:22:@18655.4]
  wire [31:0] nbufFF_io_rPort_0_output_0; // @[NBuffers.scala 298:22:@18655.4]
  wire [31:0] nbufFF_io_wPort_0_data_0; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_io_wPort_0_reset; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_io_wPort_0_en_0; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_io_sEn_0; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_io_sEn_1; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_io_sEn_2; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_io_sEn_3; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_io_sEn_4; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_io_sEn_5; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_io_sEn_6; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_io_sDone_0; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_io_sDone_1; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_io_sDone_2; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_io_sDone_3; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_io_sDone_4; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_io_sDone_5; // @[NBuffers.scala 298:22:@18655.4]
  wire  nbufFF_io_sDone_6; // @[NBuffers.scala 298:22:@18655.4]
  NBuf_2 nbufFF ( // @[NBuffers.scala 298:22:@18655.4]
    .clock(nbufFF_clock),
    .reset(nbufFF_reset),
    .io_rPort_5_output_0(nbufFF_io_rPort_5_output_0),
    .io_rPort_4_output_0(nbufFF_io_rPort_4_output_0),
    .io_rPort_3_output_0(nbufFF_io_rPort_3_output_0),
    .io_rPort_2_output_0(nbufFF_io_rPort_2_output_0),
    .io_rPort_1_output_0(nbufFF_io_rPort_1_output_0),
    .io_rPort_0_output_0(nbufFF_io_rPort_0_output_0),
    .io_wPort_0_data_0(nbufFF_io_wPort_0_data_0),
    .io_wPort_0_reset(nbufFF_io_wPort_0_reset),
    .io_wPort_0_en_0(nbufFF_io_wPort_0_en_0),
    .io_sEn_0(nbufFF_io_sEn_0),
    .io_sEn_1(nbufFF_io_sEn_1),
    .io_sEn_2(nbufFF_io_sEn_2),
    .io_sEn_3(nbufFF_io_sEn_3),
    .io_sEn_4(nbufFF_io_sEn_4),
    .io_sEn_5(nbufFF_io_sEn_5),
    .io_sEn_6(nbufFF_io_sEn_6),
    .io_sDone_0(nbufFF_io_sDone_0),
    .io_sDone_1(nbufFF_io_sDone_1),
    .io_sDone_2(nbufFF_io_sDone_2),
    .io_sDone_3(nbufFF_io_sDone_3),
    .io_sDone_4(nbufFF_io_sDone_4),
    .io_sDone_5(nbufFF_io_sDone_5),
    .io_sDone_6(nbufFF_io_sDone_6)
  );
  assign io_rPort_5_output_0 = nbufFF_io_rPort_5_output_0; // @[NBuffers.scala 299:6:@18712.4]
  assign io_rPort_4_output_0 = nbufFF_io_rPort_4_output_0; // @[NBuffers.scala 299:6:@18707.4]
  assign io_rPort_3_output_0 = nbufFF_io_rPort_3_output_0; // @[NBuffers.scala 299:6:@18702.4]
  assign io_rPort_2_output_0 = nbufFF_io_rPort_2_output_0; // @[NBuffers.scala 299:6:@18697.4]
  assign io_rPort_1_output_0 = nbufFF_io_rPort_1_output_0; // @[NBuffers.scala 299:6:@18692.4]
  assign io_rPort_0_output_0 = nbufFF_io_rPort_0_output_0; // @[NBuffers.scala 299:6:@18687.4]
  assign nbufFF_clock = clock; // @[:@18656.4]
  assign nbufFF_reset = reset; // @[:@18657.4]
  assign nbufFF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[NBuffers.scala 299:6:@18684.4]
  assign nbufFF_io_wPort_0_reset = io_wPort_0_reset; // @[NBuffers.scala 299:6:@18683.4]
  assign nbufFF_io_wPort_0_en_0 = io_wPort_0_en_0; // @[NBuffers.scala 299:6:@18680.4]
  assign nbufFF_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 299:6:@18665.4]
  assign nbufFF_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 299:6:@18666.4]
  assign nbufFF_io_sEn_2 = io_sEn_2; // @[NBuffers.scala 299:6:@18667.4]
  assign nbufFF_io_sEn_3 = io_sEn_3; // @[NBuffers.scala 299:6:@18668.4]
  assign nbufFF_io_sEn_4 = io_sEn_4; // @[NBuffers.scala 299:6:@18669.4]
  assign nbufFF_io_sEn_5 = io_sEn_5; // @[NBuffers.scala 299:6:@18670.4]
  assign nbufFF_io_sEn_6 = io_sEn_6; // @[NBuffers.scala 299:6:@18671.4]
  assign nbufFF_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 299:6:@18658.4]
  assign nbufFF_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 299:6:@18659.4]
  assign nbufFF_io_sDone_2 = io_sDone_2; // @[NBuffers.scala 299:6:@18660.4]
  assign nbufFF_io_sDone_3 = io_sDone_3; // @[NBuffers.scala 299:6:@18661.4]
  assign nbufFF_io_sDone_4 = io_sDone_4; // @[NBuffers.scala 299:6:@18662.4]
  assign nbufFF_io_sDone_5 = io_sDone_5; // @[NBuffers.scala 299:6:@18663.4]
  assign nbufFF_io_sDone_6 = io_sDone_6; // @[NBuffers.scala 299:6:@18664.4]
endmodule
module FF_20( // @[:@21122.2]
  input   clock, // @[:@21123.4]
  input   reset, // @[:@21124.4]
  output  io_rPort_4_output_0, // @[:@21125.4]
  output  io_rPort_3_output_0, // @[:@21125.4]
  output  io_rPort_1_output_0, // @[:@21125.4]
  output  io_rPort_0_output_0, // @[:@21125.4]
  input   io_wPort_0_data_0, // @[:@21125.4]
  input   io_wPort_0_reset, // @[:@21125.4]
  input   io_wPort_0_en_0 // @[:@21125.4]
);
  reg  ff; // @[MemPrimitives.scala 321:19:@21165.4]
  reg [31:0] _RAND_0;
  wire  _T_198; // @[MemPrimitives.scala 325:32:@21167.4]
  wire  _T_199; // @[MemPrimitives.scala 325:12:@21168.4]
  assign _T_198 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@21167.4]
  assign _T_199 = io_wPort_0_reset ? 1'h0 : _T_198; // @[MemPrimitives.scala 325:12:@21168.4]
  assign io_rPort_4_output_0 = ff; // @[MemPrimitives.scala 326:34:@21174.4]
  assign io_rPort_3_output_0 = ff; // @[MemPrimitives.scala 326:34:@21173.4]
  assign io_rPort_1_output_0 = ff; // @[MemPrimitives.scala 326:34:@21171.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@21170.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 1'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 1'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module NBuf_3( // @[:@21507.2]
  input   clock, // @[:@21508.4]
  input   reset, // @[:@21509.4]
  output  io_rPort_4_output_0, // @[:@21510.4]
  output  io_rPort_3_output_0, // @[:@21510.4]
  output  io_rPort_1_output_0, // @[:@21510.4]
  output  io_rPort_0_output_0, // @[:@21510.4]
  input   io_wPort_0_data_0, // @[:@21510.4]
  input   io_wPort_0_reset, // @[:@21510.4]
  input   io_wPort_0_en_0, // @[:@21510.4]
  input   io_sEn_0, // @[:@21510.4]
  input   io_sEn_1, // @[:@21510.4]
  input   io_sEn_2, // @[:@21510.4]
  input   io_sEn_3, // @[:@21510.4]
  input   io_sEn_4, // @[:@21510.4]
  input   io_sEn_5, // @[:@21510.4]
  input   io_sEn_6, // @[:@21510.4]
  input   io_sDone_0, // @[:@21510.4]
  input   io_sDone_1, // @[:@21510.4]
  input   io_sDone_2, // @[:@21510.4]
  input   io_sDone_3, // @[:@21510.4]
  input   io_sDone_4, // @[:@21510.4]
  input   io_sDone_5, // @[:@21510.4]
  input   io_sDone_6 // @[:@21510.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@21518.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@21518.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@21518.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@21518.4]
  wire  ctrl_io_sEn_2; // @[NBuffers.scala 83:20:@21518.4]
  wire  ctrl_io_sEn_3; // @[NBuffers.scala 83:20:@21518.4]
  wire  ctrl_io_sEn_4; // @[NBuffers.scala 83:20:@21518.4]
  wire  ctrl_io_sEn_5; // @[NBuffers.scala 83:20:@21518.4]
  wire  ctrl_io_sEn_6; // @[NBuffers.scala 83:20:@21518.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@21518.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@21518.4]
  wire  ctrl_io_sDone_2; // @[NBuffers.scala 83:20:@21518.4]
  wire  ctrl_io_sDone_3; // @[NBuffers.scala 83:20:@21518.4]
  wire  ctrl_io_sDone_4; // @[NBuffers.scala 83:20:@21518.4]
  wire  ctrl_io_sDone_5; // @[NBuffers.scala 83:20:@21518.4]
  wire  ctrl_io_sDone_6; // @[NBuffers.scala 83:20:@21518.4]
  wire [3:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@21518.4]
  wire [3:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@21518.4]
  wire [3:0] ctrl_io_statesInR_2; // @[NBuffers.scala 83:20:@21518.4]
  wire [3:0] ctrl_io_statesInR_3; // @[NBuffers.scala 83:20:@21518.4]
  wire [3:0] ctrl_io_statesInR_4; // @[NBuffers.scala 83:20:@21518.4]
  wire [3:0] ctrl_io_statesInR_5; // @[NBuffers.scala 83:20:@21518.4]
  wire [3:0] ctrl_io_statesInR_6; // @[NBuffers.scala 83:20:@21518.4]
  wire  FF_clock; // @[NBuffers.scala 146:23:@21535.4]
  wire  FF_reset; // @[NBuffers.scala 146:23:@21535.4]
  wire  FF_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@21535.4]
  wire  FF_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@21535.4]
  wire  FF_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@21535.4]
  wire  FF_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@21535.4]
  wire  FF_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@21535.4]
  wire  FF_io_wPort_0_reset; // @[NBuffers.scala 146:23:@21535.4]
  wire  FF_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@21535.4]
  wire  FF_1_clock; // @[NBuffers.scala 146:23:@21576.4]
  wire  FF_1_reset; // @[NBuffers.scala 146:23:@21576.4]
  wire  FF_1_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@21576.4]
  wire  FF_1_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@21576.4]
  wire  FF_1_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@21576.4]
  wire  FF_1_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@21576.4]
  wire  FF_1_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@21576.4]
  wire  FF_1_io_wPort_0_reset; // @[NBuffers.scala 146:23:@21576.4]
  wire  FF_1_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@21576.4]
  wire  FF_2_clock; // @[NBuffers.scala 146:23:@21617.4]
  wire  FF_2_reset; // @[NBuffers.scala 146:23:@21617.4]
  wire  FF_2_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@21617.4]
  wire  FF_2_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@21617.4]
  wire  FF_2_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@21617.4]
  wire  FF_2_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@21617.4]
  wire  FF_2_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@21617.4]
  wire  FF_2_io_wPort_0_reset; // @[NBuffers.scala 146:23:@21617.4]
  wire  FF_2_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@21617.4]
  wire  FF_3_clock; // @[NBuffers.scala 146:23:@21658.4]
  wire  FF_3_reset; // @[NBuffers.scala 146:23:@21658.4]
  wire  FF_3_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@21658.4]
  wire  FF_3_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@21658.4]
  wire  FF_3_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@21658.4]
  wire  FF_3_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@21658.4]
  wire  FF_3_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@21658.4]
  wire  FF_3_io_wPort_0_reset; // @[NBuffers.scala 146:23:@21658.4]
  wire  FF_3_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@21658.4]
  wire  FF_4_clock; // @[NBuffers.scala 146:23:@21699.4]
  wire  FF_4_reset; // @[NBuffers.scala 146:23:@21699.4]
  wire  FF_4_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@21699.4]
  wire  FF_4_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@21699.4]
  wire  FF_4_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@21699.4]
  wire  FF_4_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@21699.4]
  wire  FF_4_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@21699.4]
  wire  FF_4_io_wPort_0_reset; // @[NBuffers.scala 146:23:@21699.4]
  wire  FF_4_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@21699.4]
  wire  FF_5_clock; // @[NBuffers.scala 146:23:@21740.4]
  wire  FF_5_reset; // @[NBuffers.scala 146:23:@21740.4]
  wire  FF_5_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@21740.4]
  wire  FF_5_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@21740.4]
  wire  FF_5_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@21740.4]
  wire  FF_5_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@21740.4]
  wire  FF_5_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@21740.4]
  wire  FF_5_io_wPort_0_reset; // @[NBuffers.scala 146:23:@21740.4]
  wire  FF_5_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@21740.4]
  wire  FF_6_clock; // @[NBuffers.scala 146:23:@21781.4]
  wire  FF_6_reset; // @[NBuffers.scala 146:23:@21781.4]
  wire  FF_6_io_rPort_4_output_0; // @[NBuffers.scala 146:23:@21781.4]
  wire  FF_6_io_rPort_3_output_0; // @[NBuffers.scala 146:23:@21781.4]
  wire  FF_6_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@21781.4]
  wire  FF_6_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@21781.4]
  wire  FF_6_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@21781.4]
  wire  FF_6_io_wPort_0_reset; // @[NBuffers.scala 146:23:@21781.4]
  wire  FF_6_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@21781.4]
  wire  _T_236; // @[NBuffers.scala 153:105:@21829.4]
  wire  _T_240; // @[NBuffers.scala 157:92:@21839.4]
  wire  _T_243; // @[NBuffers.scala 157:92:@21845.4]
  wire  _T_249; // @[NBuffers.scala 157:92:@21857.4]
  wire  _T_252; // @[NBuffers.scala 157:92:@21863.4]
  wire  _T_258; // @[NBuffers.scala 153:105:@21875.4]
  wire  _T_262; // @[NBuffers.scala 157:92:@21885.4]
  wire  _T_265; // @[NBuffers.scala 157:92:@21891.4]
  wire  _T_271; // @[NBuffers.scala 157:92:@21903.4]
  wire  _T_274; // @[NBuffers.scala 157:92:@21909.4]
  wire  _T_280; // @[NBuffers.scala 153:105:@21921.4]
  wire  _T_284; // @[NBuffers.scala 157:92:@21931.4]
  wire  _T_287; // @[NBuffers.scala 157:92:@21937.4]
  wire  _T_293; // @[NBuffers.scala 157:92:@21949.4]
  wire  _T_296; // @[NBuffers.scala 157:92:@21955.4]
  wire  _T_302; // @[NBuffers.scala 153:105:@21967.4]
  wire  _T_306; // @[NBuffers.scala 157:92:@21977.4]
  wire  _T_309; // @[NBuffers.scala 157:92:@21983.4]
  wire  _T_315; // @[NBuffers.scala 157:92:@21995.4]
  wire  _T_318; // @[NBuffers.scala 157:92:@22001.4]
  wire  _T_324; // @[NBuffers.scala 153:105:@22013.4]
  wire  _T_328; // @[NBuffers.scala 157:92:@22023.4]
  wire  _T_331; // @[NBuffers.scala 157:92:@22029.4]
  wire  _T_337; // @[NBuffers.scala 157:92:@22041.4]
  wire  _T_340; // @[NBuffers.scala 157:92:@22047.4]
  wire  _T_346; // @[NBuffers.scala 153:105:@22059.4]
  wire  _T_350; // @[NBuffers.scala 157:92:@22069.4]
  wire  _T_353; // @[NBuffers.scala 157:92:@22075.4]
  wire  _T_359; // @[NBuffers.scala 157:92:@22087.4]
  wire  _T_362; // @[NBuffers.scala 157:92:@22093.4]
  wire  _T_368; // @[NBuffers.scala 153:105:@22105.4]
  wire  _T_372; // @[NBuffers.scala 157:92:@22115.4]
  wire  _T_375; // @[NBuffers.scala 157:92:@22121.4]
  wire  _T_381; // @[NBuffers.scala 157:92:@22133.4]
  wire  _T_384; // @[NBuffers.scala 157:92:@22139.4]
  wire  _T_405; // @[Mux.scala 19:72:@22158.4]
  wire  _T_407; // @[Mux.scala 19:72:@22159.4]
  wire  _T_409; // @[Mux.scala 19:72:@22160.4]
  wire  _T_411; // @[Mux.scala 19:72:@22161.4]
  wire  _T_413; // @[Mux.scala 19:72:@22162.4]
  wire  _T_415; // @[Mux.scala 19:72:@22163.4]
  wire  _T_417; // @[Mux.scala 19:72:@22164.4]
  wire  _T_418; // @[Mux.scala 19:72:@22165.4]
  wire  _T_419; // @[Mux.scala 19:72:@22166.4]
  wire  _T_420; // @[Mux.scala 19:72:@22167.4]
  wire  _T_421; // @[Mux.scala 19:72:@22168.4]
  wire  _T_422; // @[Mux.scala 19:72:@22169.4]
  wire  _T_442; // @[Mux.scala 19:72:@22181.4]
  wire  _T_444; // @[Mux.scala 19:72:@22182.4]
  wire  _T_446; // @[Mux.scala 19:72:@22183.4]
  wire  _T_448; // @[Mux.scala 19:72:@22184.4]
  wire  _T_450; // @[Mux.scala 19:72:@22185.4]
  wire  _T_452; // @[Mux.scala 19:72:@22186.4]
  wire  _T_454; // @[Mux.scala 19:72:@22187.4]
  wire  _T_455; // @[Mux.scala 19:72:@22188.4]
  wire  _T_456; // @[Mux.scala 19:72:@22189.4]
  wire  _T_457; // @[Mux.scala 19:72:@22190.4]
  wire  _T_458; // @[Mux.scala 19:72:@22191.4]
  wire  _T_459; // @[Mux.scala 19:72:@22192.4]
  wire  _T_516; // @[Mux.scala 19:72:@22227.4]
  wire  _T_518; // @[Mux.scala 19:72:@22228.4]
  wire  _T_520; // @[Mux.scala 19:72:@22229.4]
  wire  _T_522; // @[Mux.scala 19:72:@22230.4]
  wire  _T_524; // @[Mux.scala 19:72:@22231.4]
  wire  _T_526; // @[Mux.scala 19:72:@22232.4]
  wire  _T_528; // @[Mux.scala 19:72:@22233.4]
  wire  _T_529; // @[Mux.scala 19:72:@22234.4]
  wire  _T_530; // @[Mux.scala 19:72:@22235.4]
  wire  _T_531; // @[Mux.scala 19:72:@22236.4]
  wire  _T_532; // @[Mux.scala 19:72:@22237.4]
  wire  _T_533; // @[Mux.scala 19:72:@22238.4]
  wire  _T_553; // @[Mux.scala 19:72:@22250.4]
  wire  _T_555; // @[Mux.scala 19:72:@22251.4]
  wire  _T_557; // @[Mux.scala 19:72:@22252.4]
  wire  _T_559; // @[Mux.scala 19:72:@22253.4]
  wire  _T_561; // @[Mux.scala 19:72:@22254.4]
  wire  _T_563; // @[Mux.scala 19:72:@22255.4]
  wire  _T_565; // @[Mux.scala 19:72:@22256.4]
  wire  _T_566; // @[Mux.scala 19:72:@22257.4]
  wire  _T_567; // @[Mux.scala 19:72:@22258.4]
  wire  _T_568; // @[Mux.scala 19:72:@22259.4]
  wire  _T_569; // @[Mux.scala 19:72:@22260.4]
  wire  _T_570; // @[Mux.scala 19:72:@22261.4]
  NBufController_3 ctrl ( // @[NBuffers.scala 83:20:@21518.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sEn_2(ctrl_io_sEn_2),
    .io_sEn_3(ctrl_io_sEn_3),
    .io_sEn_4(ctrl_io_sEn_4),
    .io_sEn_5(ctrl_io_sEn_5),
    .io_sEn_6(ctrl_io_sEn_6),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_sDone_2(ctrl_io_sDone_2),
    .io_sDone_3(ctrl_io_sDone_3),
    .io_sDone_4(ctrl_io_sDone_4),
    .io_sDone_5(ctrl_io_sDone_5),
    .io_sDone_6(ctrl_io_sDone_6),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1),
    .io_statesInR_2(ctrl_io_statesInR_2),
    .io_statesInR_3(ctrl_io_statesInR_3),
    .io_statesInR_4(ctrl_io_statesInR_4),
    .io_statesInR_5(ctrl_io_statesInR_5),
    .io_statesInR_6(ctrl_io_statesInR_6)
  );
  FF_20 FF ( // @[NBuffers.scala 146:23:@21535.4]
    .clock(FF_clock),
    .reset(FF_reset),
    .io_rPort_4_output_0(FF_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_io_rPort_3_output_0),
    .io_rPort_1_output_0(FF_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_io_wPort_0_en_0)
  );
  FF_20 FF_1 ( // @[NBuffers.scala 146:23:@21576.4]
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_rPort_4_output_0(FF_1_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_1_io_rPort_3_output_0),
    .io_rPort_1_output_0(FF_1_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_1_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_1_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_1_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_1_io_wPort_0_en_0)
  );
  FF_20 FF_2 ( // @[NBuffers.scala 146:23:@21617.4]
    .clock(FF_2_clock),
    .reset(FF_2_reset),
    .io_rPort_4_output_0(FF_2_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_2_io_rPort_3_output_0),
    .io_rPort_1_output_0(FF_2_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_2_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_2_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_2_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_2_io_wPort_0_en_0)
  );
  FF_20 FF_3 ( // @[NBuffers.scala 146:23:@21658.4]
    .clock(FF_3_clock),
    .reset(FF_3_reset),
    .io_rPort_4_output_0(FF_3_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_3_io_rPort_3_output_0),
    .io_rPort_1_output_0(FF_3_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_3_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_3_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_3_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_3_io_wPort_0_en_0)
  );
  FF_20 FF_4 ( // @[NBuffers.scala 146:23:@21699.4]
    .clock(FF_4_clock),
    .reset(FF_4_reset),
    .io_rPort_4_output_0(FF_4_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_4_io_rPort_3_output_0),
    .io_rPort_1_output_0(FF_4_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_4_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_4_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_4_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_4_io_wPort_0_en_0)
  );
  FF_20 FF_5 ( // @[NBuffers.scala 146:23:@21740.4]
    .clock(FF_5_clock),
    .reset(FF_5_reset),
    .io_rPort_4_output_0(FF_5_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_5_io_rPort_3_output_0),
    .io_rPort_1_output_0(FF_5_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_5_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_5_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_5_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_5_io_wPort_0_en_0)
  );
  FF_20 FF_6 ( // @[NBuffers.scala 146:23:@21781.4]
    .clock(FF_6_clock),
    .reset(FF_6_reset),
    .io_rPort_4_output_0(FF_6_io_rPort_4_output_0),
    .io_rPort_3_output_0(FF_6_io_rPort_3_output_0),
    .io_rPort_1_output_0(FF_6_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_6_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_6_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_6_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_6_io_wPort_0_en_0)
  );
  assign _T_236 = ctrl_io_statesInW_0 == 4'h0; // @[NBuffers.scala 153:105:@21829.4]
  assign _T_240 = ctrl_io_statesInR_1 == 4'h0; // @[NBuffers.scala 157:92:@21839.4]
  assign _T_243 = ctrl_io_statesInR_2 == 4'h0; // @[NBuffers.scala 157:92:@21845.4]
  assign _T_249 = ctrl_io_statesInR_4 == 4'h0; // @[NBuffers.scala 157:92:@21857.4]
  assign _T_252 = ctrl_io_statesInR_5 == 4'h0; // @[NBuffers.scala 157:92:@21863.4]
  assign _T_258 = ctrl_io_statesInW_0 == 4'h1; // @[NBuffers.scala 153:105:@21875.4]
  assign _T_262 = ctrl_io_statesInR_1 == 4'h1; // @[NBuffers.scala 157:92:@21885.4]
  assign _T_265 = ctrl_io_statesInR_2 == 4'h1; // @[NBuffers.scala 157:92:@21891.4]
  assign _T_271 = ctrl_io_statesInR_4 == 4'h1; // @[NBuffers.scala 157:92:@21903.4]
  assign _T_274 = ctrl_io_statesInR_5 == 4'h1; // @[NBuffers.scala 157:92:@21909.4]
  assign _T_280 = ctrl_io_statesInW_0 == 4'h2; // @[NBuffers.scala 153:105:@21921.4]
  assign _T_284 = ctrl_io_statesInR_1 == 4'h2; // @[NBuffers.scala 157:92:@21931.4]
  assign _T_287 = ctrl_io_statesInR_2 == 4'h2; // @[NBuffers.scala 157:92:@21937.4]
  assign _T_293 = ctrl_io_statesInR_4 == 4'h2; // @[NBuffers.scala 157:92:@21949.4]
  assign _T_296 = ctrl_io_statesInR_5 == 4'h2; // @[NBuffers.scala 157:92:@21955.4]
  assign _T_302 = ctrl_io_statesInW_0 == 4'h3; // @[NBuffers.scala 153:105:@21967.4]
  assign _T_306 = ctrl_io_statesInR_1 == 4'h3; // @[NBuffers.scala 157:92:@21977.4]
  assign _T_309 = ctrl_io_statesInR_2 == 4'h3; // @[NBuffers.scala 157:92:@21983.4]
  assign _T_315 = ctrl_io_statesInR_4 == 4'h3; // @[NBuffers.scala 157:92:@21995.4]
  assign _T_318 = ctrl_io_statesInR_5 == 4'h3; // @[NBuffers.scala 157:92:@22001.4]
  assign _T_324 = ctrl_io_statesInW_0 == 4'h4; // @[NBuffers.scala 153:105:@22013.4]
  assign _T_328 = ctrl_io_statesInR_1 == 4'h4; // @[NBuffers.scala 157:92:@22023.4]
  assign _T_331 = ctrl_io_statesInR_2 == 4'h4; // @[NBuffers.scala 157:92:@22029.4]
  assign _T_337 = ctrl_io_statesInR_4 == 4'h4; // @[NBuffers.scala 157:92:@22041.4]
  assign _T_340 = ctrl_io_statesInR_5 == 4'h4; // @[NBuffers.scala 157:92:@22047.4]
  assign _T_346 = ctrl_io_statesInW_0 == 4'h5; // @[NBuffers.scala 153:105:@22059.4]
  assign _T_350 = ctrl_io_statesInR_1 == 4'h5; // @[NBuffers.scala 157:92:@22069.4]
  assign _T_353 = ctrl_io_statesInR_2 == 4'h5; // @[NBuffers.scala 157:92:@22075.4]
  assign _T_359 = ctrl_io_statesInR_4 == 4'h5; // @[NBuffers.scala 157:92:@22087.4]
  assign _T_362 = ctrl_io_statesInR_5 == 4'h5; // @[NBuffers.scala 157:92:@22093.4]
  assign _T_368 = ctrl_io_statesInW_0 == 4'h6; // @[NBuffers.scala 153:105:@22105.4]
  assign _T_372 = ctrl_io_statesInR_1 == 4'h6; // @[NBuffers.scala 157:92:@22115.4]
  assign _T_375 = ctrl_io_statesInR_2 == 4'h6; // @[NBuffers.scala 157:92:@22121.4]
  assign _T_381 = ctrl_io_statesInR_4 == 4'h6; // @[NBuffers.scala 157:92:@22133.4]
  assign _T_384 = ctrl_io_statesInR_5 == 4'h6; // @[NBuffers.scala 157:92:@22139.4]
  assign _T_405 = _T_240 ? FF_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@22158.4]
  assign _T_407 = _T_262 ? FF_1_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@22159.4]
  assign _T_409 = _T_284 ? FF_2_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@22160.4]
  assign _T_411 = _T_306 ? FF_3_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@22161.4]
  assign _T_413 = _T_328 ? FF_4_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@22162.4]
  assign _T_415 = _T_350 ? FF_5_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@22163.4]
  assign _T_417 = _T_372 ? FF_6_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@22164.4]
  assign _T_418 = _T_405 | _T_407; // @[Mux.scala 19:72:@22165.4]
  assign _T_419 = _T_418 | _T_409; // @[Mux.scala 19:72:@22166.4]
  assign _T_420 = _T_419 | _T_411; // @[Mux.scala 19:72:@22167.4]
  assign _T_421 = _T_420 | _T_413; // @[Mux.scala 19:72:@22168.4]
  assign _T_422 = _T_421 | _T_415; // @[Mux.scala 19:72:@22169.4]
  assign _T_442 = _T_243 ? FF_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@22181.4]
  assign _T_444 = _T_265 ? FF_1_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@22182.4]
  assign _T_446 = _T_287 ? FF_2_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@22183.4]
  assign _T_448 = _T_309 ? FF_3_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@22184.4]
  assign _T_450 = _T_331 ? FF_4_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@22185.4]
  assign _T_452 = _T_353 ? FF_5_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@22186.4]
  assign _T_454 = _T_375 ? FF_6_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@22187.4]
  assign _T_455 = _T_442 | _T_444; // @[Mux.scala 19:72:@22188.4]
  assign _T_456 = _T_455 | _T_446; // @[Mux.scala 19:72:@22189.4]
  assign _T_457 = _T_456 | _T_448; // @[Mux.scala 19:72:@22190.4]
  assign _T_458 = _T_457 | _T_450; // @[Mux.scala 19:72:@22191.4]
  assign _T_459 = _T_458 | _T_452; // @[Mux.scala 19:72:@22192.4]
  assign _T_516 = _T_249 ? FF_io_rPort_3_output_0 : 1'h0; // @[Mux.scala 19:72:@22227.4]
  assign _T_518 = _T_271 ? FF_1_io_rPort_3_output_0 : 1'h0; // @[Mux.scala 19:72:@22228.4]
  assign _T_520 = _T_293 ? FF_2_io_rPort_3_output_0 : 1'h0; // @[Mux.scala 19:72:@22229.4]
  assign _T_522 = _T_315 ? FF_3_io_rPort_3_output_0 : 1'h0; // @[Mux.scala 19:72:@22230.4]
  assign _T_524 = _T_337 ? FF_4_io_rPort_3_output_0 : 1'h0; // @[Mux.scala 19:72:@22231.4]
  assign _T_526 = _T_359 ? FF_5_io_rPort_3_output_0 : 1'h0; // @[Mux.scala 19:72:@22232.4]
  assign _T_528 = _T_381 ? FF_6_io_rPort_3_output_0 : 1'h0; // @[Mux.scala 19:72:@22233.4]
  assign _T_529 = _T_516 | _T_518; // @[Mux.scala 19:72:@22234.4]
  assign _T_530 = _T_529 | _T_520; // @[Mux.scala 19:72:@22235.4]
  assign _T_531 = _T_530 | _T_522; // @[Mux.scala 19:72:@22236.4]
  assign _T_532 = _T_531 | _T_524; // @[Mux.scala 19:72:@22237.4]
  assign _T_533 = _T_532 | _T_526; // @[Mux.scala 19:72:@22238.4]
  assign _T_553 = _T_252 ? FF_io_rPort_4_output_0 : 1'h0; // @[Mux.scala 19:72:@22250.4]
  assign _T_555 = _T_274 ? FF_1_io_rPort_4_output_0 : 1'h0; // @[Mux.scala 19:72:@22251.4]
  assign _T_557 = _T_296 ? FF_2_io_rPort_4_output_0 : 1'h0; // @[Mux.scala 19:72:@22252.4]
  assign _T_559 = _T_318 ? FF_3_io_rPort_4_output_0 : 1'h0; // @[Mux.scala 19:72:@22253.4]
  assign _T_561 = _T_340 ? FF_4_io_rPort_4_output_0 : 1'h0; // @[Mux.scala 19:72:@22254.4]
  assign _T_563 = _T_362 ? FF_5_io_rPort_4_output_0 : 1'h0; // @[Mux.scala 19:72:@22255.4]
  assign _T_565 = _T_384 ? FF_6_io_rPort_4_output_0 : 1'h0; // @[Mux.scala 19:72:@22256.4]
  assign _T_566 = _T_553 | _T_555; // @[Mux.scala 19:72:@22257.4]
  assign _T_567 = _T_566 | _T_557; // @[Mux.scala 19:72:@22258.4]
  assign _T_568 = _T_567 | _T_559; // @[Mux.scala 19:72:@22259.4]
  assign _T_569 = _T_568 | _T_561; // @[Mux.scala 19:72:@22260.4]
  assign _T_570 = _T_569 | _T_563; // @[Mux.scala 19:72:@22261.4]
  assign io_rPort_4_output_0 = _T_570 | _T_565; // @[NBuffers.scala 163:66:@22265.4]
  assign io_rPort_3_output_0 = _T_533 | _T_528; // @[NBuffers.scala 163:66:@22242.4]
  assign io_rPort_1_output_0 = _T_459 | _T_454; // @[NBuffers.scala 163:66:@22196.4]
  assign io_rPort_0_output_0 = _T_422 | _T_417; // @[NBuffers.scala 163:66:@22173.4]
  assign ctrl_clock = clock; // @[:@21519.4]
  assign ctrl_reset = reset; // @[:@21520.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@21521.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@21523.4]
  assign ctrl_io_sEn_2 = io_sEn_2; // @[NBuffers.scala 85:20:@21525.4]
  assign ctrl_io_sEn_3 = io_sEn_3; // @[NBuffers.scala 85:20:@21527.4]
  assign ctrl_io_sEn_4 = io_sEn_4; // @[NBuffers.scala 85:20:@21529.4]
  assign ctrl_io_sEn_5 = io_sEn_5; // @[NBuffers.scala 85:20:@21531.4]
  assign ctrl_io_sEn_6 = io_sEn_6; // @[NBuffers.scala 85:20:@21533.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@21522.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@21524.4]
  assign ctrl_io_sDone_2 = io_sDone_2; // @[NBuffers.scala 86:22:@21526.4]
  assign ctrl_io_sDone_3 = io_sDone_3; // @[NBuffers.scala 86:22:@21528.4]
  assign ctrl_io_sDone_4 = io_sDone_4; // @[NBuffers.scala 86:22:@21530.4]
  assign ctrl_io_sDone_5 = io_sDone_5; // @[NBuffers.scala 86:22:@21532.4]
  assign ctrl_io_sDone_6 = io_sDone_6; // @[NBuffers.scala 86:22:@21534.4]
  assign FF_clock = clock; // @[:@21536.4]
  assign FF_reset = reset; // @[:@21537.4]
  assign FF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@21832.4]
  assign FF_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@21833.4]
  assign FF_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_236; // @[MemPrimitives.scala 37:29:@21838.4]
  assign FF_1_clock = clock; // @[:@21577.4]
  assign FF_1_reset = reset; // @[:@21578.4]
  assign FF_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@21878.4]
  assign FF_1_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@21879.4]
  assign FF_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_258; // @[MemPrimitives.scala 37:29:@21884.4]
  assign FF_2_clock = clock; // @[:@21618.4]
  assign FF_2_reset = reset; // @[:@21619.4]
  assign FF_2_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@21924.4]
  assign FF_2_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@21925.4]
  assign FF_2_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_280; // @[MemPrimitives.scala 37:29:@21930.4]
  assign FF_3_clock = clock; // @[:@21659.4]
  assign FF_3_reset = reset; // @[:@21660.4]
  assign FF_3_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@21970.4]
  assign FF_3_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@21971.4]
  assign FF_3_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_302; // @[MemPrimitives.scala 37:29:@21976.4]
  assign FF_4_clock = clock; // @[:@21700.4]
  assign FF_4_reset = reset; // @[:@21701.4]
  assign FF_4_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@22016.4]
  assign FF_4_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@22017.4]
  assign FF_4_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_324; // @[MemPrimitives.scala 37:29:@22022.4]
  assign FF_5_clock = clock; // @[:@21741.4]
  assign FF_5_reset = reset; // @[:@21742.4]
  assign FF_5_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@22062.4]
  assign FF_5_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@22063.4]
  assign FF_5_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_346; // @[MemPrimitives.scala 37:29:@22068.4]
  assign FF_6_clock = clock; // @[:@21782.4]
  assign FF_6_reset = reset; // @[:@21783.4]
  assign FF_6_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@22108.4]
  assign FF_6_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@22109.4]
  assign FF_6_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_368; // @[MemPrimitives.scala 37:29:@22114.4]
endmodule
module b552_chain( // @[:@22290.2]
  input   clock, // @[:@22291.4]
  input   reset, // @[:@22292.4]
  output  io_rPort_4_output_0, // @[:@22293.4]
  output  io_rPort_3_output_0, // @[:@22293.4]
  output  io_rPort_1_output_0, // @[:@22293.4]
  output  io_rPort_0_output_0, // @[:@22293.4]
  input   io_wPort_0_data_0, // @[:@22293.4]
  input   io_wPort_0_reset, // @[:@22293.4]
  input   io_wPort_0_en_0, // @[:@22293.4]
  input   io_sEn_0, // @[:@22293.4]
  input   io_sEn_1, // @[:@22293.4]
  input   io_sEn_2, // @[:@22293.4]
  input   io_sEn_3, // @[:@22293.4]
  input   io_sEn_4, // @[:@22293.4]
  input   io_sEn_5, // @[:@22293.4]
  input   io_sEn_6, // @[:@22293.4]
  input   io_sDone_0, // @[:@22293.4]
  input   io_sDone_1, // @[:@22293.4]
  input   io_sDone_2, // @[:@22293.4]
  input   io_sDone_3, // @[:@22293.4]
  input   io_sDone_4, // @[:@22293.4]
  input   io_sDone_5, // @[:@22293.4]
  input   io_sDone_6 // @[:@22293.4]
);
  wire  nbufFF_clock; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_reset; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_rPort_4_output_0; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_rPort_3_output_0; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_rPort_1_output_0; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_rPort_0_output_0; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_wPort_0_data_0; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_wPort_0_reset; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_wPort_0_en_0; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_sEn_0; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_sEn_1; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_sEn_2; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_sEn_3; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_sEn_4; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_sEn_5; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_sEn_6; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_sDone_0; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_sDone_1; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_sDone_2; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_sDone_3; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_sDone_4; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_sDone_5; // @[NBuffers.scala 298:22:@22301.4]
  wire  nbufFF_io_sDone_6; // @[NBuffers.scala 298:22:@22301.4]
  NBuf_3 nbufFF ( // @[NBuffers.scala 298:22:@22301.4]
    .clock(nbufFF_clock),
    .reset(nbufFF_reset),
    .io_rPort_4_output_0(nbufFF_io_rPort_4_output_0),
    .io_rPort_3_output_0(nbufFF_io_rPort_3_output_0),
    .io_rPort_1_output_0(nbufFF_io_rPort_1_output_0),
    .io_rPort_0_output_0(nbufFF_io_rPort_0_output_0),
    .io_wPort_0_data_0(nbufFF_io_wPort_0_data_0),
    .io_wPort_0_reset(nbufFF_io_wPort_0_reset),
    .io_wPort_0_en_0(nbufFF_io_wPort_0_en_0),
    .io_sEn_0(nbufFF_io_sEn_0),
    .io_sEn_1(nbufFF_io_sEn_1),
    .io_sEn_2(nbufFF_io_sEn_2),
    .io_sEn_3(nbufFF_io_sEn_3),
    .io_sEn_4(nbufFF_io_sEn_4),
    .io_sEn_5(nbufFF_io_sEn_5),
    .io_sEn_6(nbufFF_io_sEn_6),
    .io_sDone_0(nbufFF_io_sDone_0),
    .io_sDone_1(nbufFF_io_sDone_1),
    .io_sDone_2(nbufFF_io_sDone_2),
    .io_sDone_3(nbufFF_io_sDone_3),
    .io_sDone_4(nbufFF_io_sDone_4),
    .io_sDone_5(nbufFF_io_sDone_5),
    .io_sDone_6(nbufFF_io_sDone_6)
  );
  assign io_rPort_4_output_0 = nbufFF_io_rPort_4_output_0; // @[NBuffers.scala 299:6:@22353.4]
  assign io_rPort_3_output_0 = nbufFF_io_rPort_3_output_0; // @[NBuffers.scala 299:6:@22348.4]
  assign io_rPort_1_output_0 = nbufFF_io_rPort_1_output_0; // @[NBuffers.scala 299:6:@22338.4]
  assign io_rPort_0_output_0 = nbufFF_io_rPort_0_output_0; // @[NBuffers.scala 299:6:@22333.4]
  assign nbufFF_clock = clock; // @[:@22302.4]
  assign nbufFF_reset = reset; // @[:@22303.4]
  assign nbufFF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[NBuffers.scala 299:6:@22330.4]
  assign nbufFF_io_wPort_0_reset = io_wPort_0_reset; // @[NBuffers.scala 299:6:@22329.4]
  assign nbufFF_io_wPort_0_en_0 = io_wPort_0_en_0; // @[NBuffers.scala 299:6:@22326.4]
  assign nbufFF_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 299:6:@22311.4]
  assign nbufFF_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 299:6:@22312.4]
  assign nbufFF_io_sEn_2 = io_sEn_2; // @[NBuffers.scala 299:6:@22313.4]
  assign nbufFF_io_sEn_3 = io_sEn_3; // @[NBuffers.scala 299:6:@22314.4]
  assign nbufFF_io_sEn_4 = io_sEn_4; // @[NBuffers.scala 299:6:@22315.4]
  assign nbufFF_io_sEn_5 = io_sEn_5; // @[NBuffers.scala 299:6:@22316.4]
  assign nbufFF_io_sEn_6 = io_sEn_6; // @[NBuffers.scala 299:6:@22317.4]
  assign nbufFF_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 299:6:@22304.4]
  assign nbufFF_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 299:6:@22305.4]
  assign nbufFF_io_sDone_2 = io_sDone_2; // @[NBuffers.scala 299:6:@22306.4]
  assign nbufFF_io_sDone_3 = io_sDone_3; // @[NBuffers.scala 299:6:@22307.4]
  assign nbufFF_io_sDone_4 = io_sDone_4; // @[NBuffers.scala 299:6:@22308.4]
  assign nbufFF_io_sDone_5 = io_sDone_5; // @[NBuffers.scala 299:6:@22309.4]
  assign nbufFF_io_sDone_6 = io_sDone_6; // @[NBuffers.scala 299:6:@22310.4]
endmodule
module RetimeWrapper_248( // @[:@23332.2]
  input         clock, // @[:@23333.4]
  input         reset, // @[:@23334.4]
  input         io_flow, // @[:@23335.4]
  input  [31:0] io_in, // @[:@23335.4]
  output [31:0] io_out // @[:@23335.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@23337.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@23337.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@23337.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@23337.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@23337.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@23337.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@23337.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@23350.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@23349.4]
  assign sr_init = 32'h5; // @[RetimeShiftRegister.scala 19:16:@23348.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@23347.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@23346.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@23344.4]
endmodule
module NBufCtr_25( // @[:@23352.2]
  input         clock, // @[:@23353.4]
  input         reset, // @[:@23354.4]
  input         io_input_countUp, // @[:@23355.4]
  input         io_input_enable, // @[:@23355.4]
  output [31:0] io_output_count // @[:@23355.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@23392.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@23392.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@23392.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@23392.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@23392.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@23397.4 package.scala 96:25:@23398.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@23358.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@23359.4]
  wire  _T_21; // @[Counter.scala 49:55:@23360.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@23361.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@23362.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@23363.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@23364.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@23365.4]
  wire  _T_33; // @[Counter.scala 51:52:@23369.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@23370.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@23371.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@23372.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@23373.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@23374.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@23375.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@23376.4]
  wire  _T_45; // @[Counter.scala 52:70:@23377.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@23379.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@23380.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@23381.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@23382.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@23383.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@23384.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@23387.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@23388.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@23390.4]
  RetimeWrapper_248 RetimeWrapper ( // @[package.scala 93:22:@23392.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@23397.4 package.scala 96:25:@23398.4]
  assign _T_18 = {{1'd0}, _T_66}; // @[Counter.scala 49:32:@23358.4]
  assign _T_19 = _T_18[31:0]; // @[Counter.scala 49:32:@23359.4]
  assign _T_21 = _T_19 >= 32'h6; // @[Counter.scala 49:55:@23360.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@23361.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 49:91:@23362.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh6); // @[Counter.scala 49:91:@23363.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@23364.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@23365.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@23369.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@23370.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@23371.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@23372.4]
  assign _T_39 = _T_33 ? 32'h5 : _T_38; // @[Counter.scala 51:47:@23373.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@23374.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@23375.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@23376.4]
  assign _T_45 = _T_43 >= 32'h6; // @[Counter.scala 52:70:@23377.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@23379.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@23380.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@23381.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@23382.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@23383.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@23384.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@23387.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@23388.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@23390.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@23400.4]
  assign RetimeWrapper_clock = clock; // @[:@23393.4]
  assign RetimeWrapper_reset = reset; // @[:@23394.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@23396.4]
  assign RetimeWrapper_io_in = reset ? 32'h5 : _T_62; // @[package.scala 94:16:@23395.4]
endmodule
module NBufCtr_26( // @[:@23434.2]
  input         clock, // @[:@23435.4]
  input         reset, // @[:@23436.4]
  input         io_input_countUp, // @[:@23437.4]
  input         io_input_enable, // @[:@23437.4]
  output [31:0] io_output_count // @[:@23437.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@23474.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@23474.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@23474.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@23474.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@23474.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@23479.4 package.scala 96:25:@23480.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@23440.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@23441.4]
  wire  _T_21; // @[Counter.scala 49:55:@23442.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@23443.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@23444.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@23445.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@23446.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@23447.4]
  wire  _T_33; // @[Counter.scala 51:52:@23451.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@23452.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@23453.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@23454.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@23455.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@23456.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@23457.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@23458.4]
  wire  _T_45; // @[Counter.scala 52:70:@23459.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@23461.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@23462.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@23463.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@23464.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@23465.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@23466.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@23469.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@23470.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@23472.4]
  RetimeWrapper_248 RetimeWrapper ( // @[package.scala 93:22:@23474.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@23479.4 package.scala 96:25:@23480.4]
  assign _T_18 = _T_66 + 32'h5; // @[Counter.scala 49:32:@23440.4]
  assign _T_19 = _T_66 + 32'h5; // @[Counter.scala 49:32:@23441.4]
  assign _T_21 = _T_19 >= 32'h6; // @[Counter.scala 49:55:@23442.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@23443.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 49:91:@23444.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 49:91:@23445.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@23446.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@23447.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@23451.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@23452.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@23453.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@23454.4]
  assign _T_39 = _T_33 ? 32'h5 : _T_38; // @[Counter.scala 51:47:@23455.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@23456.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@23457.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@23458.4]
  assign _T_45 = _T_43 >= 32'h6; // @[Counter.scala 52:70:@23459.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@23461.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@23462.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@23463.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@23464.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@23465.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@23466.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@23469.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@23470.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@23472.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@23482.4]
  assign RetimeWrapper_clock = clock; // @[:@23475.4]
  assign RetimeWrapper_reset = reset; // @[:@23476.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@23478.4]
  assign RetimeWrapper_io_in = reset ? 32'h5 : _T_62; // @[package.scala 94:16:@23477.4]
endmodule
module NBufCtr_28( // @[:@23598.2]
  input         clock, // @[:@23599.4]
  input         reset, // @[:@23600.4]
  input         io_input_countUp, // @[:@23601.4]
  input         io_input_enable, // @[:@23601.4]
  output [31:0] io_output_count // @[:@23601.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@23638.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@23638.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@23638.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@23638.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@23638.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@23643.4 package.scala 96:25:@23644.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@23604.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@23605.4]
  wire  _T_21; // @[Counter.scala 49:55:@23606.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@23607.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@23608.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@23609.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@23610.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@23611.4]
  wire  _T_33; // @[Counter.scala 51:52:@23615.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@23616.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@23617.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@23618.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@23619.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@23620.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@23629.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@23630.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@23633.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@23634.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@23636.4]
  RetimeWrapper_248 RetimeWrapper ( // @[package.scala 93:22:@23638.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@23643.4 package.scala 96:25:@23644.4]
  assign _T_18 = _T_66 + 32'h1; // @[Counter.scala 49:32:@23604.4]
  assign _T_19 = _T_66 + 32'h1; // @[Counter.scala 49:32:@23605.4]
  assign _T_21 = _T_19 >= 32'h6; // @[Counter.scala 49:55:@23606.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@23607.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 49:91:@23608.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 49:91:@23609.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@23610.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@23611.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@23615.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@23616.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@23617.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@23618.4]
  assign _T_39 = _T_33 ? 32'h5 : _T_38; // @[Counter.scala 51:47:@23619.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@23620.4]
  assign _T_53 = {{1'd0}, _T_27}; // @[Counter.scala 52:107:@23629.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@23630.4]
  assign _T_58 = _T_21 ? _T_54 : _T_19; // @[Counter.scala 52:45:@23633.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@23634.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@23636.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@23646.4]
  assign RetimeWrapper_clock = clock; // @[:@23639.4]
  assign RetimeWrapper_reset = reset; // @[:@23640.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@23642.4]
  assign RetimeWrapper_io_in = reset ? 32'h5 : _T_62; // @[package.scala 94:16:@23641.4]
endmodule
module NBufCtr_29( // @[:@23680.2]
  input   clock, // @[:@23681.4]
  input   reset, // @[:@23682.4]
  input   io_input_countUp, // @[:@23683.4]
  input   io_input_enable // @[:@23683.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@23720.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@23720.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@23720.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@23720.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@23720.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@23725.4 package.scala 96:25:@23726.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@23689.4]
  wire  _T_33; // @[Counter.scala 51:52:@23697.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@23698.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@23699.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@23700.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@23701.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@23702.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@23703.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@23704.4]
  wire  _T_45; // @[Counter.scala 52:70:@23705.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@23707.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@23708.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@23709.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@23710.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@23711.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@23712.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@23715.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@23716.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@23718.4]
  RetimeWrapper_248 RetimeWrapper ( // @[package.scala 93:22:@23720.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@23725.4 package.scala 96:25:@23726.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@23689.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@23697.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@23698.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@23699.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@23700.4]
  assign _T_39 = _T_33 ? 32'h5 : _T_38; // @[Counter.scala 51:47:@23701.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@23702.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@23703.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@23704.4]
  assign _T_45 = _T_43 >= 32'h6; // @[Counter.scala 52:70:@23705.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@23707.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@23708.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@23709.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@23710.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@23711.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@23712.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@23715.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@23716.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@23718.4]
  assign RetimeWrapper_clock = clock; // @[:@23721.4]
  assign RetimeWrapper_reset = reset; // @[:@23722.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@23724.4]
  assign RetimeWrapper_io_in = reset ? 32'h5 : _T_62; // @[package.scala 94:16:@23723.4]
endmodule
module NBufCtr_30( // @[:@23762.2]
  input   clock, // @[:@23763.4]
  input   reset, // @[:@23764.4]
  input   io_input_countUp, // @[:@23765.4]
  input   io_input_enable // @[:@23765.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@23802.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@23802.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@23802.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@23802.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@23802.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@23807.4 package.scala 96:25:@23808.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@23771.4]
  wire  _T_33; // @[Counter.scala 51:52:@23779.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@23780.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@23781.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@23782.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@23783.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@23784.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@23785.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@23786.4]
  wire  _T_45; // @[Counter.scala 52:70:@23787.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@23789.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@23790.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@23791.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@23792.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@23793.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@23794.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@23797.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@23798.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@23800.4]
  RetimeWrapper_248 RetimeWrapper ( // @[package.scala 93:22:@23802.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@23807.4 package.scala 96:25:@23808.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@23771.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@23779.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@23780.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@23781.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@23782.4]
  assign _T_39 = _T_33 ? 32'h5 : _T_38; // @[Counter.scala 51:47:@23783.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@23784.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@23785.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@23786.4]
  assign _T_45 = _T_43 >= 32'h6; // @[Counter.scala 52:70:@23787.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@23789.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@23790.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@23791.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@23792.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@23793.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@23794.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@23797.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@23798.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@23800.4]
  assign RetimeWrapper_clock = clock; // @[:@23803.4]
  assign RetimeWrapper_reset = reset; // @[:@23804.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@23806.4]
  assign RetimeWrapper_io_in = reset ? 32'h5 : _T_62; // @[package.scala 94:16:@23805.4]
endmodule
module NBufCtr_31( // @[:@23844.2]
  input   clock, // @[:@23845.4]
  input   reset, // @[:@23846.4]
  input   io_input_countUp, // @[:@23847.4]
  input   io_input_enable // @[:@23847.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@23884.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@23884.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@23884.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@23884.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@23884.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@23889.4 package.scala 96:25:@23890.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@23853.4]
  wire  _T_33; // @[Counter.scala 51:52:@23861.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@23862.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@23863.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@23864.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@23865.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@23866.4]
  wire [32:0] _T_42; // @[Counter.scala 52:50:@23867.4]
  wire [31:0] _T_43; // @[Counter.scala 52:50:@23868.4]
  wire  _T_45; // @[Counter.scala 52:70:@23869.4]
  wire [32:0] _T_49; // @[Counter.scala 52:121:@23871.4]
  wire [31:0] _T_50; // @[Counter.scala 52:121:@23872.4]
  wire [31:0] _T_51; // @[Counter.scala 52:121:@23873.4]
  wire [31:0] _T_52; // @[Counter.scala 52:155:@23874.4]
  wire [32:0] _T_53; // @[Counter.scala 52:107:@23875.4]
  wire [31:0] _T_54; // @[Counter.scala 52:107:@23876.4]
  wire [31:0] _T_58; // @[Counter.scala 52:45:@23879.4]
  wire [31:0] _T_59; // @[Counter.scala 52:24:@23880.4]
  wire [31:0] _T_62; // @[Counter.scala 53:52:@23882.4]
  RetimeWrapper_248 RetimeWrapper ( // @[package.scala 93:22:@23884.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@23889.4 package.scala 96:25:@23890.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@23853.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@23861.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@23862.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@23863.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@23864.4]
  assign _T_39 = _T_33 ? 32'h5 : _T_38; // @[Counter.scala 51:47:@23865.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@23866.4]
  assign _T_42 = _T_66 + 32'h1; // @[Counter.scala 52:50:@23867.4]
  assign _T_43 = _T_66 + 32'h1; // @[Counter.scala 52:50:@23868.4]
  assign _T_45 = _T_43 >= 32'h6; // @[Counter.scala 52:70:@23869.4]
  assign _T_49 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@23871.4]
  assign _T_50 = $signed(_T_22) + $signed(-32'sh5); // @[Counter.scala 52:121:@23872.4]
  assign _T_51 = $signed(_T_50); // @[Counter.scala 52:121:@23873.4]
  assign _T_52 = $unsigned(_T_51); // @[Counter.scala 52:155:@23874.4]
  assign _T_53 = {{1'd0}, _T_52}; // @[Counter.scala 52:107:@23875.4]
  assign _T_54 = _T_53[31:0]; // @[Counter.scala 52:107:@23876.4]
  assign _T_58 = _T_45 ? _T_54 : _T_43; // @[Counter.scala 52:45:@23879.4]
  assign _T_59 = io_input_enable ? _T_58 : _T_66; // @[Counter.scala 52:24:@23880.4]
  assign _T_62 = io_input_countUp ? _T_59 : _T_40; // @[Counter.scala 53:52:@23882.4]
  assign RetimeWrapper_clock = clock; // @[:@23885.4]
  assign RetimeWrapper_reset = reset; // @[:@23886.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@23888.4]
  assign RetimeWrapper_io_in = reset ? 32'h5 : _T_62; // @[package.scala 94:16:@23887.4]
endmodule
module NBufController_5( // @[:@23976.2]
  input        clock, // @[:@23977.4]
  input        reset, // @[:@23978.4]
  input        io_sEn_0, // @[:@23979.4]
  input        io_sEn_1, // @[:@23979.4]
  input        io_sEn_2, // @[:@23979.4]
  input        io_sEn_3, // @[:@23979.4]
  input        io_sEn_4, // @[:@23979.4]
  input        io_sEn_5, // @[:@23979.4]
  input        io_sDone_0, // @[:@23979.4]
  input        io_sDone_1, // @[:@23979.4]
  input        io_sDone_2, // @[:@23979.4]
  input        io_sDone_3, // @[:@23979.4]
  input        io_sDone_4, // @[:@23979.4]
  input        io_sDone_5, // @[:@23979.4]
  output [3:0] io_statesInW_0, // @[:@23979.4]
  output [3:0] io_statesInW_1, // @[:@23979.4]
  output [3:0] io_statesInR_1, // @[:@23979.4]
  output [3:0] io_statesInR_5 // @[:@23979.4]
);
  wire  sEn_latch_0_clock; // @[NBuffers.scala 21:52:@23981.4]
  wire  sEn_latch_0_reset; // @[NBuffers.scala 21:52:@23981.4]
  wire  sEn_latch_0_io_input_set; // @[NBuffers.scala 21:52:@23981.4]
  wire  sEn_latch_0_io_input_reset; // @[NBuffers.scala 21:52:@23981.4]
  wire  sEn_latch_0_io_input_asyn_reset; // @[NBuffers.scala 21:52:@23981.4]
  wire  sEn_latch_0_io_output; // @[NBuffers.scala 21:52:@23981.4]
  wire  sEn_latch_1_clock; // @[NBuffers.scala 21:52:@23984.4]
  wire  sEn_latch_1_reset; // @[NBuffers.scala 21:52:@23984.4]
  wire  sEn_latch_1_io_input_set; // @[NBuffers.scala 21:52:@23984.4]
  wire  sEn_latch_1_io_input_reset; // @[NBuffers.scala 21:52:@23984.4]
  wire  sEn_latch_1_io_input_asyn_reset; // @[NBuffers.scala 21:52:@23984.4]
  wire  sEn_latch_1_io_output; // @[NBuffers.scala 21:52:@23984.4]
  wire  sEn_latch_2_clock; // @[NBuffers.scala 21:52:@23987.4]
  wire  sEn_latch_2_reset; // @[NBuffers.scala 21:52:@23987.4]
  wire  sEn_latch_2_io_input_set; // @[NBuffers.scala 21:52:@23987.4]
  wire  sEn_latch_2_io_input_reset; // @[NBuffers.scala 21:52:@23987.4]
  wire  sEn_latch_2_io_input_asyn_reset; // @[NBuffers.scala 21:52:@23987.4]
  wire  sEn_latch_2_io_output; // @[NBuffers.scala 21:52:@23987.4]
  wire  sEn_latch_3_clock; // @[NBuffers.scala 21:52:@23990.4]
  wire  sEn_latch_3_reset; // @[NBuffers.scala 21:52:@23990.4]
  wire  sEn_latch_3_io_input_set; // @[NBuffers.scala 21:52:@23990.4]
  wire  sEn_latch_3_io_input_reset; // @[NBuffers.scala 21:52:@23990.4]
  wire  sEn_latch_3_io_input_asyn_reset; // @[NBuffers.scala 21:52:@23990.4]
  wire  sEn_latch_3_io_output; // @[NBuffers.scala 21:52:@23990.4]
  wire  sEn_latch_4_clock; // @[NBuffers.scala 21:52:@23993.4]
  wire  sEn_latch_4_reset; // @[NBuffers.scala 21:52:@23993.4]
  wire  sEn_latch_4_io_input_set; // @[NBuffers.scala 21:52:@23993.4]
  wire  sEn_latch_4_io_input_reset; // @[NBuffers.scala 21:52:@23993.4]
  wire  sEn_latch_4_io_input_asyn_reset; // @[NBuffers.scala 21:52:@23993.4]
  wire  sEn_latch_4_io_output; // @[NBuffers.scala 21:52:@23993.4]
  wire  sEn_latch_5_clock; // @[NBuffers.scala 21:52:@23996.4]
  wire  sEn_latch_5_reset; // @[NBuffers.scala 21:52:@23996.4]
  wire  sEn_latch_5_io_input_set; // @[NBuffers.scala 21:52:@23996.4]
  wire  sEn_latch_5_io_input_reset; // @[NBuffers.scala 21:52:@23996.4]
  wire  sEn_latch_5_io_input_asyn_reset; // @[NBuffers.scala 21:52:@23996.4]
  wire  sEn_latch_5_io_output; // @[NBuffers.scala 21:52:@23996.4]
  wire  sDone_latch_0_clock; // @[NBuffers.scala 22:54:@23999.4]
  wire  sDone_latch_0_reset; // @[NBuffers.scala 22:54:@23999.4]
  wire  sDone_latch_0_io_input_set; // @[NBuffers.scala 22:54:@23999.4]
  wire  sDone_latch_0_io_input_reset; // @[NBuffers.scala 22:54:@23999.4]
  wire  sDone_latch_0_io_input_asyn_reset; // @[NBuffers.scala 22:54:@23999.4]
  wire  sDone_latch_0_io_output; // @[NBuffers.scala 22:54:@23999.4]
  wire  sDone_latch_1_clock; // @[NBuffers.scala 22:54:@24002.4]
  wire  sDone_latch_1_reset; // @[NBuffers.scala 22:54:@24002.4]
  wire  sDone_latch_1_io_input_set; // @[NBuffers.scala 22:54:@24002.4]
  wire  sDone_latch_1_io_input_reset; // @[NBuffers.scala 22:54:@24002.4]
  wire  sDone_latch_1_io_input_asyn_reset; // @[NBuffers.scala 22:54:@24002.4]
  wire  sDone_latch_1_io_output; // @[NBuffers.scala 22:54:@24002.4]
  wire  sDone_latch_2_clock; // @[NBuffers.scala 22:54:@24005.4]
  wire  sDone_latch_2_reset; // @[NBuffers.scala 22:54:@24005.4]
  wire  sDone_latch_2_io_input_set; // @[NBuffers.scala 22:54:@24005.4]
  wire  sDone_latch_2_io_input_reset; // @[NBuffers.scala 22:54:@24005.4]
  wire  sDone_latch_2_io_input_asyn_reset; // @[NBuffers.scala 22:54:@24005.4]
  wire  sDone_latch_2_io_output; // @[NBuffers.scala 22:54:@24005.4]
  wire  sDone_latch_3_clock; // @[NBuffers.scala 22:54:@24008.4]
  wire  sDone_latch_3_reset; // @[NBuffers.scala 22:54:@24008.4]
  wire  sDone_latch_3_io_input_set; // @[NBuffers.scala 22:54:@24008.4]
  wire  sDone_latch_3_io_input_reset; // @[NBuffers.scala 22:54:@24008.4]
  wire  sDone_latch_3_io_input_asyn_reset; // @[NBuffers.scala 22:54:@24008.4]
  wire  sDone_latch_3_io_output; // @[NBuffers.scala 22:54:@24008.4]
  wire  sDone_latch_4_clock; // @[NBuffers.scala 22:54:@24011.4]
  wire  sDone_latch_4_reset; // @[NBuffers.scala 22:54:@24011.4]
  wire  sDone_latch_4_io_input_set; // @[NBuffers.scala 22:54:@24011.4]
  wire  sDone_latch_4_io_input_reset; // @[NBuffers.scala 22:54:@24011.4]
  wire  sDone_latch_4_io_input_asyn_reset; // @[NBuffers.scala 22:54:@24011.4]
  wire  sDone_latch_4_io_output; // @[NBuffers.scala 22:54:@24011.4]
  wire  sDone_latch_5_clock; // @[NBuffers.scala 22:54:@24014.4]
  wire  sDone_latch_5_reset; // @[NBuffers.scala 22:54:@24014.4]
  wire  sDone_latch_5_io_input_set; // @[NBuffers.scala 22:54:@24014.4]
  wire  sDone_latch_5_io_input_reset; // @[NBuffers.scala 22:54:@24014.4]
  wire  sDone_latch_5_io_input_asyn_reset; // @[NBuffers.scala 22:54:@24014.4]
  wire  sDone_latch_5_io_output; // @[NBuffers.scala 22:54:@24014.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@24021.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@24021.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@24021.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@24021.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@24021.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@24029.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@24029.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@24029.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@24029.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@24029.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@24038.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@24038.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@24038.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@24038.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@24038.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@24046.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@24046.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@24046.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@24046.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@24046.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@24057.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@24057.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@24057.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@24057.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@24057.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@24065.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@24065.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@24065.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@24065.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@24065.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@24074.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@24074.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@24074.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@24074.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@24074.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@24082.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@24082.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@24082.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@24082.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@24082.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@24093.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@24093.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@24093.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@24093.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@24093.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@24101.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@24101.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@24101.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@24101.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@24101.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@24110.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@24110.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@24110.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@24110.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@24110.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@24118.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@24118.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@24118.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@24118.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@24118.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@24129.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@24129.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@24129.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@24129.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@24129.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@24137.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@24137.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@24137.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@24137.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@24137.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@24146.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@24146.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@24146.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@24146.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@24146.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@24154.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@24154.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@24154.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@24154.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@24154.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@24165.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@24165.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@24165.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@24165.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@24165.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@24173.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@24173.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@24173.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@24173.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@24173.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@24182.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@24182.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@24182.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@24182.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@24182.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@24190.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@24190.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@24190.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@24190.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@24190.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@24201.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@24201.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@24201.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@24201.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@24201.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@24209.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@24209.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@24209.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@24209.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@24209.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@24218.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@24218.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@24218.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@24218.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@24218.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@24226.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@24226.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@24226.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@24226.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@24226.4]
  wire  NBufCtr_clock; // @[NBuffers.scala 40:19:@24263.4]
  wire  NBufCtr_reset; // @[NBuffers.scala 40:19:@24263.4]
  wire  NBufCtr_io_input_countUp; // @[NBuffers.scala 40:19:@24263.4]
  wire  NBufCtr_io_input_enable; // @[NBuffers.scala 40:19:@24263.4]
  wire [31:0] NBufCtr_io_output_count; // @[NBuffers.scala 40:19:@24263.4]
  wire  NBufCtr_1_clock; // @[NBuffers.scala 40:19:@24274.4]
  wire  NBufCtr_1_reset; // @[NBuffers.scala 40:19:@24274.4]
  wire  NBufCtr_1_io_input_countUp; // @[NBuffers.scala 40:19:@24274.4]
  wire  NBufCtr_1_io_input_enable; // @[NBuffers.scala 40:19:@24274.4]
  wire [31:0] NBufCtr_1_io_output_count; // @[NBuffers.scala 40:19:@24274.4]
  wire  statesInR_0_clock; // @[NBuffers.scala 50:19:@24285.4]
  wire  statesInR_0_reset; // @[NBuffers.scala 50:19:@24285.4]
  wire  statesInR_0_io_input_countUp; // @[NBuffers.scala 50:19:@24285.4]
  wire  statesInR_0_io_input_enable; // @[NBuffers.scala 50:19:@24285.4]
  wire [31:0] statesInR_0_io_output_count; // @[NBuffers.scala 50:19:@24285.4]
  wire  statesInR_1_clock; // @[NBuffers.scala 50:19:@24296.4]
  wire  statesInR_1_reset; // @[NBuffers.scala 50:19:@24296.4]
  wire  statesInR_1_io_input_countUp; // @[NBuffers.scala 50:19:@24296.4]
  wire  statesInR_1_io_input_enable; // @[NBuffers.scala 50:19:@24296.4]
  wire [31:0] statesInR_1_io_output_count; // @[NBuffers.scala 50:19:@24296.4]
  wire  statesInR_2_clock; // @[NBuffers.scala 50:19:@24307.4]
  wire  statesInR_2_reset; // @[NBuffers.scala 50:19:@24307.4]
  wire  statesInR_2_io_input_countUp; // @[NBuffers.scala 50:19:@24307.4]
  wire  statesInR_2_io_input_enable; // @[NBuffers.scala 50:19:@24307.4]
  wire  statesInR_3_clock; // @[NBuffers.scala 50:19:@24318.4]
  wire  statesInR_3_reset; // @[NBuffers.scala 50:19:@24318.4]
  wire  statesInR_3_io_input_countUp; // @[NBuffers.scala 50:19:@24318.4]
  wire  statesInR_3_io_input_enable; // @[NBuffers.scala 50:19:@24318.4]
  wire  statesInR_4_clock; // @[NBuffers.scala 50:19:@24329.4]
  wire  statesInR_4_reset; // @[NBuffers.scala 50:19:@24329.4]
  wire  statesInR_4_io_input_countUp; // @[NBuffers.scala 50:19:@24329.4]
  wire  statesInR_4_io_input_enable; // @[NBuffers.scala 50:19:@24329.4]
  wire  statesInR_5_clock; // @[NBuffers.scala 50:19:@24340.4]
  wire  statesInR_5_reset; // @[NBuffers.scala 50:19:@24340.4]
  wire  statesInR_5_io_input_countUp; // @[NBuffers.scala 50:19:@24340.4]
  wire  statesInR_5_io_input_enable; // @[NBuffers.scala 50:19:@24340.4]
  wire [31:0] statesInR_5_io_output_count; // @[NBuffers.scala 50:19:@24340.4]
  wire  _T_33; // @[NBuffers.scala 26:46:@24018.4]
  wire  _T_48; // @[NBuffers.scala 26:46:@24054.4]
  wire  _T_63; // @[NBuffers.scala 26:46:@24090.4]
  wire  _T_78; // @[NBuffers.scala 26:46:@24126.4]
  wire  _T_93; // @[NBuffers.scala 26:46:@24162.4]
  wire  _T_108; // @[NBuffers.scala 26:46:@24198.4]
  wire  _T_122; // @[NBuffers.scala 33:64:@24234.4]
  wire  _T_123; // @[NBuffers.scala 33:64:@24235.4]
  wire  _T_124; // @[NBuffers.scala 33:64:@24236.4]
  wire  _T_125; // @[NBuffers.scala 33:64:@24237.4]
  wire  anyEnabled; // @[NBuffers.scala 33:64:@24238.4]
  wire  _T_126; // @[NBuffers.scala 34:124:@24239.4]
  wire  _T_127; // @[NBuffers.scala 34:104:@24240.4]
  wire  _T_128; // @[NBuffers.scala 34:124:@24241.4]
  wire  _T_129; // @[NBuffers.scala 34:104:@24242.4]
  wire  _T_130; // @[NBuffers.scala 34:124:@24243.4]
  wire  _T_131; // @[NBuffers.scala 34:104:@24244.4]
  wire  _T_132; // @[NBuffers.scala 34:124:@24245.4]
  wire  _T_133; // @[NBuffers.scala 34:104:@24246.4]
  wire  _T_134; // @[NBuffers.scala 34:124:@24247.4]
  wire  _T_135; // @[NBuffers.scala 34:104:@24248.4]
  wire  _T_136; // @[NBuffers.scala 34:124:@24249.4]
  wire  _T_137; // @[NBuffers.scala 34:104:@24250.4]
  wire  _T_138; // @[NBuffers.scala 34:150:@24251.4]
  wire  _T_139; // @[NBuffers.scala 34:150:@24252.4]
  wire  _T_140; // @[NBuffers.scala 34:150:@24253.4]
  wire  _T_141; // @[NBuffers.scala 34:150:@24254.4]
  wire  _T_142; // @[NBuffers.scala 34:150:@24255.4]
  wire  _T_143; // @[NBuffers.scala 34:154:@24256.4]
  wire  _T_145; // @[package.scala 100:49:@24257.4]
  reg  _T_148; // @[package.scala 48:56:@24258.4]
  reg [31:0] _RAND_0;
  SRFF sEn_latch_0 ( // @[NBuffers.scala 21:52:@23981.4]
    .clock(sEn_latch_0_clock),
    .reset(sEn_latch_0_reset),
    .io_input_set(sEn_latch_0_io_input_set),
    .io_input_reset(sEn_latch_0_io_input_reset),
    .io_input_asyn_reset(sEn_latch_0_io_input_asyn_reset),
    .io_output(sEn_latch_0_io_output)
  );
  SRFF sEn_latch_1 ( // @[NBuffers.scala 21:52:@23984.4]
    .clock(sEn_latch_1_clock),
    .reset(sEn_latch_1_reset),
    .io_input_set(sEn_latch_1_io_input_set),
    .io_input_reset(sEn_latch_1_io_input_reset),
    .io_input_asyn_reset(sEn_latch_1_io_input_asyn_reset),
    .io_output(sEn_latch_1_io_output)
  );
  SRFF sEn_latch_2 ( // @[NBuffers.scala 21:52:@23987.4]
    .clock(sEn_latch_2_clock),
    .reset(sEn_latch_2_reset),
    .io_input_set(sEn_latch_2_io_input_set),
    .io_input_reset(sEn_latch_2_io_input_reset),
    .io_input_asyn_reset(sEn_latch_2_io_input_asyn_reset),
    .io_output(sEn_latch_2_io_output)
  );
  SRFF sEn_latch_3 ( // @[NBuffers.scala 21:52:@23990.4]
    .clock(sEn_latch_3_clock),
    .reset(sEn_latch_3_reset),
    .io_input_set(sEn_latch_3_io_input_set),
    .io_input_reset(sEn_latch_3_io_input_reset),
    .io_input_asyn_reset(sEn_latch_3_io_input_asyn_reset),
    .io_output(sEn_latch_3_io_output)
  );
  SRFF sEn_latch_4 ( // @[NBuffers.scala 21:52:@23993.4]
    .clock(sEn_latch_4_clock),
    .reset(sEn_latch_4_reset),
    .io_input_set(sEn_latch_4_io_input_set),
    .io_input_reset(sEn_latch_4_io_input_reset),
    .io_input_asyn_reset(sEn_latch_4_io_input_asyn_reset),
    .io_output(sEn_latch_4_io_output)
  );
  SRFF sEn_latch_5 ( // @[NBuffers.scala 21:52:@23996.4]
    .clock(sEn_latch_5_clock),
    .reset(sEn_latch_5_reset),
    .io_input_set(sEn_latch_5_io_input_set),
    .io_input_reset(sEn_latch_5_io_input_reset),
    .io_input_asyn_reset(sEn_latch_5_io_input_asyn_reset),
    .io_output(sEn_latch_5_io_output)
  );
  SRFF sDone_latch_0 ( // @[NBuffers.scala 22:54:@23999.4]
    .clock(sDone_latch_0_clock),
    .reset(sDone_latch_0_reset),
    .io_input_set(sDone_latch_0_io_input_set),
    .io_input_reset(sDone_latch_0_io_input_reset),
    .io_input_asyn_reset(sDone_latch_0_io_input_asyn_reset),
    .io_output(sDone_latch_0_io_output)
  );
  SRFF sDone_latch_1 ( // @[NBuffers.scala 22:54:@24002.4]
    .clock(sDone_latch_1_clock),
    .reset(sDone_latch_1_reset),
    .io_input_set(sDone_latch_1_io_input_set),
    .io_input_reset(sDone_latch_1_io_input_reset),
    .io_input_asyn_reset(sDone_latch_1_io_input_asyn_reset),
    .io_output(sDone_latch_1_io_output)
  );
  SRFF sDone_latch_2 ( // @[NBuffers.scala 22:54:@24005.4]
    .clock(sDone_latch_2_clock),
    .reset(sDone_latch_2_reset),
    .io_input_set(sDone_latch_2_io_input_set),
    .io_input_reset(sDone_latch_2_io_input_reset),
    .io_input_asyn_reset(sDone_latch_2_io_input_asyn_reset),
    .io_output(sDone_latch_2_io_output)
  );
  SRFF sDone_latch_3 ( // @[NBuffers.scala 22:54:@24008.4]
    .clock(sDone_latch_3_clock),
    .reset(sDone_latch_3_reset),
    .io_input_set(sDone_latch_3_io_input_set),
    .io_input_reset(sDone_latch_3_io_input_reset),
    .io_input_asyn_reset(sDone_latch_3_io_input_asyn_reset),
    .io_output(sDone_latch_3_io_output)
  );
  SRFF sDone_latch_4 ( // @[NBuffers.scala 22:54:@24011.4]
    .clock(sDone_latch_4_clock),
    .reset(sDone_latch_4_reset),
    .io_input_set(sDone_latch_4_io_input_set),
    .io_input_reset(sDone_latch_4_io_input_reset),
    .io_input_asyn_reset(sDone_latch_4_io_input_asyn_reset),
    .io_output(sDone_latch_4_io_output)
  );
  SRFF sDone_latch_5 ( // @[NBuffers.scala 22:54:@24014.4]
    .clock(sDone_latch_5_clock),
    .reset(sDone_latch_5_reset),
    .io_input_set(sDone_latch_5_io_input_set),
    .io_input_reset(sDone_latch_5_io_input_reset),
    .io_input_asyn_reset(sDone_latch_5_io_input_asyn_reset),
    .io_output(sDone_latch_5_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@24021.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@24029.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@24038.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@24046.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@24057.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@24065.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@24074.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@24082.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@24093.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@24101.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@24110.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 ( // @[package.scala 93:22:@24118.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper RetimeWrapper_12 ( // @[package.scala 93:22:@24129.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 ( // @[package.scala 93:22:@24137.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@24146.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@24154.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 ( // @[package.scala 93:22:@24165.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper RetimeWrapper_17 ( // @[package.scala 93:22:@24173.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 ( // @[package.scala 93:22:@24182.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper RetimeWrapper_19 ( // @[package.scala 93:22:@24190.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper RetimeWrapper_20 ( // @[package.scala 93:22:@24201.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper RetimeWrapper_21 ( // @[package.scala 93:22:@24209.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper RetimeWrapper_22 ( // @[package.scala 93:22:@24218.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper RetimeWrapper_23 ( // @[package.scala 93:22:@24226.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  NBufCtr_25 NBufCtr ( // @[NBuffers.scala 40:19:@24263.4]
    .clock(NBufCtr_clock),
    .reset(NBufCtr_reset),
    .io_input_countUp(NBufCtr_io_input_countUp),
    .io_input_enable(NBufCtr_io_input_enable),
    .io_output_count(NBufCtr_io_output_count)
  );
  NBufCtr_26 NBufCtr_1 ( // @[NBuffers.scala 40:19:@24274.4]
    .clock(NBufCtr_1_clock),
    .reset(NBufCtr_1_reset),
    .io_input_countUp(NBufCtr_1_io_input_countUp),
    .io_input_enable(NBufCtr_1_io_input_enable),
    .io_output_count(NBufCtr_1_io_output_count)
  );
  NBufCtr_25 statesInR_0 ( // @[NBuffers.scala 50:19:@24285.4]
    .clock(statesInR_0_clock),
    .reset(statesInR_0_reset),
    .io_input_countUp(statesInR_0_io_input_countUp),
    .io_input_enable(statesInR_0_io_input_enable),
    .io_output_count(statesInR_0_io_output_count)
  );
  NBufCtr_28 statesInR_1 ( // @[NBuffers.scala 50:19:@24296.4]
    .clock(statesInR_1_clock),
    .reset(statesInR_1_reset),
    .io_input_countUp(statesInR_1_io_input_countUp),
    .io_input_enable(statesInR_1_io_input_enable),
    .io_output_count(statesInR_1_io_output_count)
  );
  NBufCtr_29 statesInR_2 ( // @[NBuffers.scala 50:19:@24307.4]
    .clock(statesInR_2_clock),
    .reset(statesInR_2_reset),
    .io_input_countUp(statesInR_2_io_input_countUp),
    .io_input_enable(statesInR_2_io_input_enable)
  );
  NBufCtr_30 statesInR_3 ( // @[NBuffers.scala 50:19:@24318.4]
    .clock(statesInR_3_clock),
    .reset(statesInR_3_reset),
    .io_input_countUp(statesInR_3_io_input_countUp),
    .io_input_enable(statesInR_3_io_input_enable)
  );
  NBufCtr_31 statesInR_4 ( // @[NBuffers.scala 50:19:@24329.4]
    .clock(statesInR_4_clock),
    .reset(statesInR_4_reset),
    .io_input_countUp(statesInR_4_io_input_countUp),
    .io_input_enable(statesInR_4_io_input_enable)
  );
  NBufCtr_26 statesInR_5 ( // @[NBuffers.scala 50:19:@24340.4]
    .clock(statesInR_5_clock),
    .reset(statesInR_5_reset),
    .io_input_countUp(statesInR_5_io_input_countUp),
    .io_input_enable(statesInR_5_io_input_enable),
    .io_output_count(statesInR_5_io_output_count)
  );
  assign _T_33 = io_sDone_0 == 1'h0; // @[NBuffers.scala 26:46:@24018.4]
  assign _T_48 = io_sDone_1 == 1'h0; // @[NBuffers.scala 26:46:@24054.4]
  assign _T_63 = io_sDone_2 == 1'h0; // @[NBuffers.scala 26:46:@24090.4]
  assign _T_78 = io_sDone_3 == 1'h0; // @[NBuffers.scala 26:46:@24126.4]
  assign _T_93 = io_sDone_4 == 1'h0; // @[NBuffers.scala 26:46:@24162.4]
  assign _T_108 = io_sDone_5 == 1'h0; // @[NBuffers.scala 26:46:@24198.4]
  assign _T_122 = sEn_latch_0_io_output | sEn_latch_1_io_output; // @[NBuffers.scala 33:64:@24234.4]
  assign _T_123 = _T_122 | sEn_latch_2_io_output; // @[NBuffers.scala 33:64:@24235.4]
  assign _T_124 = _T_123 | sEn_latch_3_io_output; // @[NBuffers.scala 33:64:@24236.4]
  assign _T_125 = _T_124 | sEn_latch_4_io_output; // @[NBuffers.scala 33:64:@24237.4]
  assign anyEnabled = _T_125 | sEn_latch_5_io_output; // @[NBuffers.scala 33:64:@24238.4]
  assign _T_126 = sDone_latch_0_io_output | io_sDone_0; // @[NBuffers.scala 34:124:@24239.4]
  assign _T_127 = sEn_latch_0_io_output == _T_126; // @[NBuffers.scala 34:104:@24240.4]
  assign _T_128 = sDone_latch_1_io_output | io_sDone_1; // @[NBuffers.scala 34:124:@24241.4]
  assign _T_129 = sEn_latch_1_io_output == _T_128; // @[NBuffers.scala 34:104:@24242.4]
  assign _T_130 = sDone_latch_2_io_output | io_sDone_2; // @[NBuffers.scala 34:124:@24243.4]
  assign _T_131 = sEn_latch_2_io_output == _T_130; // @[NBuffers.scala 34:104:@24244.4]
  assign _T_132 = sDone_latch_3_io_output | io_sDone_3; // @[NBuffers.scala 34:124:@24245.4]
  assign _T_133 = sEn_latch_3_io_output == _T_132; // @[NBuffers.scala 34:104:@24246.4]
  assign _T_134 = sDone_latch_4_io_output | io_sDone_4; // @[NBuffers.scala 34:124:@24247.4]
  assign _T_135 = sEn_latch_4_io_output == _T_134; // @[NBuffers.scala 34:104:@24248.4]
  assign _T_136 = sDone_latch_5_io_output | io_sDone_5; // @[NBuffers.scala 34:124:@24249.4]
  assign _T_137 = sEn_latch_5_io_output == _T_136; // @[NBuffers.scala 34:104:@24250.4]
  assign _T_138 = _T_127 & _T_129; // @[NBuffers.scala 34:150:@24251.4]
  assign _T_139 = _T_138 & _T_131; // @[NBuffers.scala 34:150:@24252.4]
  assign _T_140 = _T_139 & _T_133; // @[NBuffers.scala 34:150:@24253.4]
  assign _T_141 = _T_140 & _T_135; // @[NBuffers.scala 34:150:@24254.4]
  assign _T_142 = _T_141 & _T_137; // @[NBuffers.scala 34:150:@24255.4]
  assign _T_143 = _T_142 & anyEnabled; // @[NBuffers.scala 34:154:@24256.4]
  assign _T_145 = _T_143 == 1'h0; // @[package.scala 100:49:@24257.4]
  assign io_statesInW_0 = NBufCtr_io_output_count[3:0]; // @[NBuffers.scala 44:21:@24273.4]
  assign io_statesInW_1 = NBufCtr_1_io_output_count[3:0]; // @[NBuffers.scala 44:21:@24284.4]
  assign io_statesInR_1 = statesInR_1_io_output_count[3:0]; // @[NBuffers.scala 54:21:@24306.4]
  assign io_statesInR_5 = statesInR_5_io_output_count[3:0]; // @[NBuffers.scala 54:21:@24350.4]
  assign sEn_latch_0_clock = clock; // @[:@23982.4]
  assign sEn_latch_0_reset = reset; // @[:@23983.4]
  assign sEn_latch_0_io_input_set = io_sEn_0 & _T_33; // @[NBuffers.scala 26:31:@24020.4]
  assign sEn_latch_0_io_input_reset = RetimeWrapper_io_out; // @[NBuffers.scala 27:33:@24028.4]
  assign sEn_latch_0_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[NBuffers.scala 28:38:@24036.4]
  assign sEn_latch_1_clock = clock; // @[:@23985.4]
  assign sEn_latch_1_reset = reset; // @[:@23986.4]
  assign sEn_latch_1_io_input_set = io_sEn_1 & _T_48; // @[NBuffers.scala 26:31:@24056.4]
  assign sEn_latch_1_io_input_reset = RetimeWrapper_4_io_out; // @[NBuffers.scala 27:33:@24064.4]
  assign sEn_latch_1_io_input_asyn_reset = RetimeWrapper_5_io_out; // @[NBuffers.scala 28:38:@24072.4]
  assign sEn_latch_2_clock = clock; // @[:@23988.4]
  assign sEn_latch_2_reset = reset; // @[:@23989.4]
  assign sEn_latch_2_io_input_set = io_sEn_2 & _T_63; // @[NBuffers.scala 26:31:@24092.4]
  assign sEn_latch_2_io_input_reset = RetimeWrapper_8_io_out; // @[NBuffers.scala 27:33:@24100.4]
  assign sEn_latch_2_io_input_asyn_reset = RetimeWrapper_9_io_out; // @[NBuffers.scala 28:38:@24108.4]
  assign sEn_latch_3_clock = clock; // @[:@23991.4]
  assign sEn_latch_3_reset = reset; // @[:@23992.4]
  assign sEn_latch_3_io_input_set = io_sEn_3 & _T_78; // @[NBuffers.scala 26:31:@24128.4]
  assign sEn_latch_3_io_input_reset = RetimeWrapper_12_io_out; // @[NBuffers.scala 27:33:@24136.4]
  assign sEn_latch_3_io_input_asyn_reset = RetimeWrapper_13_io_out; // @[NBuffers.scala 28:38:@24144.4]
  assign sEn_latch_4_clock = clock; // @[:@23994.4]
  assign sEn_latch_4_reset = reset; // @[:@23995.4]
  assign sEn_latch_4_io_input_set = io_sEn_4 & _T_93; // @[NBuffers.scala 26:31:@24164.4]
  assign sEn_latch_4_io_input_reset = RetimeWrapper_16_io_out; // @[NBuffers.scala 27:33:@24172.4]
  assign sEn_latch_4_io_input_asyn_reset = RetimeWrapper_17_io_out; // @[NBuffers.scala 28:38:@24180.4]
  assign sEn_latch_5_clock = clock; // @[:@23997.4]
  assign sEn_latch_5_reset = reset; // @[:@23998.4]
  assign sEn_latch_5_io_input_set = io_sEn_5 & _T_108; // @[NBuffers.scala 26:31:@24200.4]
  assign sEn_latch_5_io_input_reset = RetimeWrapper_20_io_out; // @[NBuffers.scala 27:33:@24208.4]
  assign sEn_latch_5_io_input_asyn_reset = RetimeWrapper_21_io_out; // @[NBuffers.scala 28:38:@24216.4]
  assign sDone_latch_0_clock = clock; // @[:@24000.4]
  assign sDone_latch_0_reset = reset; // @[:@24001.4]
  assign sDone_latch_0_io_input_set = io_sDone_0; // @[NBuffers.scala 29:33:@24037.4]
  assign sDone_latch_0_io_input_reset = RetimeWrapper_2_io_out; // @[NBuffers.scala 30:35:@24045.4]
  assign sDone_latch_0_io_input_asyn_reset = RetimeWrapper_3_io_out; // @[NBuffers.scala 31:40:@24053.4]
  assign sDone_latch_1_clock = clock; // @[:@24003.4]
  assign sDone_latch_1_reset = reset; // @[:@24004.4]
  assign sDone_latch_1_io_input_set = io_sDone_1; // @[NBuffers.scala 29:33:@24073.4]
  assign sDone_latch_1_io_input_reset = RetimeWrapper_6_io_out; // @[NBuffers.scala 30:35:@24081.4]
  assign sDone_latch_1_io_input_asyn_reset = RetimeWrapper_7_io_out; // @[NBuffers.scala 31:40:@24089.4]
  assign sDone_latch_2_clock = clock; // @[:@24006.4]
  assign sDone_latch_2_reset = reset; // @[:@24007.4]
  assign sDone_latch_2_io_input_set = io_sDone_2; // @[NBuffers.scala 29:33:@24109.4]
  assign sDone_latch_2_io_input_reset = RetimeWrapper_10_io_out; // @[NBuffers.scala 30:35:@24117.4]
  assign sDone_latch_2_io_input_asyn_reset = RetimeWrapper_11_io_out; // @[NBuffers.scala 31:40:@24125.4]
  assign sDone_latch_3_clock = clock; // @[:@24009.4]
  assign sDone_latch_3_reset = reset; // @[:@24010.4]
  assign sDone_latch_3_io_input_set = io_sDone_3; // @[NBuffers.scala 29:33:@24145.4]
  assign sDone_latch_3_io_input_reset = RetimeWrapper_14_io_out; // @[NBuffers.scala 30:35:@24153.4]
  assign sDone_latch_3_io_input_asyn_reset = RetimeWrapper_15_io_out; // @[NBuffers.scala 31:40:@24161.4]
  assign sDone_latch_4_clock = clock; // @[:@24012.4]
  assign sDone_latch_4_reset = reset; // @[:@24013.4]
  assign sDone_latch_4_io_input_set = io_sDone_4; // @[NBuffers.scala 29:33:@24181.4]
  assign sDone_latch_4_io_input_reset = RetimeWrapper_18_io_out; // @[NBuffers.scala 30:35:@24189.4]
  assign sDone_latch_4_io_input_asyn_reset = RetimeWrapper_19_io_out; // @[NBuffers.scala 31:40:@24197.4]
  assign sDone_latch_5_clock = clock; // @[:@24015.4]
  assign sDone_latch_5_reset = reset; // @[:@24016.4]
  assign sDone_latch_5_io_input_set = io_sDone_5; // @[NBuffers.scala 29:33:@24217.4]
  assign sDone_latch_5_io_input_reset = RetimeWrapper_22_io_out; // @[NBuffers.scala 30:35:@24225.4]
  assign sDone_latch_5_io_input_asyn_reset = RetimeWrapper_23_io_out; // @[NBuffers.scala 31:40:@24233.4]
  assign RetimeWrapper_clock = clock; // @[:@24022.4]
  assign RetimeWrapper_reset = reset; // @[:@24023.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@24025.4]
  assign RetimeWrapper_io_in = _T_143 & _T_148; // @[package.scala 94:16:@24024.4]
  assign RetimeWrapper_1_clock = clock; // @[:@24030.4]
  assign RetimeWrapper_1_reset = reset; // @[:@24031.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@24033.4]
  assign RetimeWrapper_1_io_in = reset; // @[package.scala 94:16:@24032.4]
  assign RetimeWrapper_2_clock = clock; // @[:@24039.4]
  assign RetimeWrapper_2_reset = reset; // @[:@24040.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@24042.4]
  assign RetimeWrapper_2_io_in = _T_143 & _T_148; // @[package.scala 94:16:@24041.4]
  assign RetimeWrapper_3_clock = clock; // @[:@24047.4]
  assign RetimeWrapper_3_reset = reset; // @[:@24048.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@24050.4]
  assign RetimeWrapper_3_io_in = reset; // @[package.scala 94:16:@24049.4]
  assign RetimeWrapper_4_clock = clock; // @[:@24058.4]
  assign RetimeWrapper_4_reset = reset; // @[:@24059.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@24061.4]
  assign RetimeWrapper_4_io_in = _T_143 & _T_148; // @[package.scala 94:16:@24060.4]
  assign RetimeWrapper_5_clock = clock; // @[:@24066.4]
  assign RetimeWrapper_5_reset = reset; // @[:@24067.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@24069.4]
  assign RetimeWrapper_5_io_in = reset; // @[package.scala 94:16:@24068.4]
  assign RetimeWrapper_6_clock = clock; // @[:@24075.4]
  assign RetimeWrapper_6_reset = reset; // @[:@24076.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@24078.4]
  assign RetimeWrapper_6_io_in = _T_143 & _T_148; // @[package.scala 94:16:@24077.4]
  assign RetimeWrapper_7_clock = clock; // @[:@24083.4]
  assign RetimeWrapper_7_reset = reset; // @[:@24084.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@24086.4]
  assign RetimeWrapper_7_io_in = reset; // @[package.scala 94:16:@24085.4]
  assign RetimeWrapper_8_clock = clock; // @[:@24094.4]
  assign RetimeWrapper_8_reset = reset; // @[:@24095.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@24097.4]
  assign RetimeWrapper_8_io_in = _T_143 & _T_148; // @[package.scala 94:16:@24096.4]
  assign RetimeWrapper_9_clock = clock; // @[:@24102.4]
  assign RetimeWrapper_9_reset = reset; // @[:@24103.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@24105.4]
  assign RetimeWrapper_9_io_in = reset; // @[package.scala 94:16:@24104.4]
  assign RetimeWrapper_10_clock = clock; // @[:@24111.4]
  assign RetimeWrapper_10_reset = reset; // @[:@24112.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@24114.4]
  assign RetimeWrapper_10_io_in = _T_143 & _T_148; // @[package.scala 94:16:@24113.4]
  assign RetimeWrapper_11_clock = clock; // @[:@24119.4]
  assign RetimeWrapper_11_reset = reset; // @[:@24120.4]
  assign RetimeWrapper_11_io_flow = 1'h1; // @[package.scala 95:18:@24122.4]
  assign RetimeWrapper_11_io_in = reset; // @[package.scala 94:16:@24121.4]
  assign RetimeWrapper_12_clock = clock; // @[:@24130.4]
  assign RetimeWrapper_12_reset = reset; // @[:@24131.4]
  assign RetimeWrapper_12_io_flow = 1'h1; // @[package.scala 95:18:@24133.4]
  assign RetimeWrapper_12_io_in = _T_143 & _T_148; // @[package.scala 94:16:@24132.4]
  assign RetimeWrapper_13_clock = clock; // @[:@24138.4]
  assign RetimeWrapper_13_reset = reset; // @[:@24139.4]
  assign RetimeWrapper_13_io_flow = 1'h1; // @[package.scala 95:18:@24141.4]
  assign RetimeWrapper_13_io_in = reset; // @[package.scala 94:16:@24140.4]
  assign RetimeWrapper_14_clock = clock; // @[:@24147.4]
  assign RetimeWrapper_14_reset = reset; // @[:@24148.4]
  assign RetimeWrapper_14_io_flow = 1'h1; // @[package.scala 95:18:@24150.4]
  assign RetimeWrapper_14_io_in = _T_143 & _T_148; // @[package.scala 94:16:@24149.4]
  assign RetimeWrapper_15_clock = clock; // @[:@24155.4]
  assign RetimeWrapper_15_reset = reset; // @[:@24156.4]
  assign RetimeWrapper_15_io_flow = 1'h1; // @[package.scala 95:18:@24158.4]
  assign RetimeWrapper_15_io_in = reset; // @[package.scala 94:16:@24157.4]
  assign RetimeWrapper_16_clock = clock; // @[:@24166.4]
  assign RetimeWrapper_16_reset = reset; // @[:@24167.4]
  assign RetimeWrapper_16_io_flow = 1'h1; // @[package.scala 95:18:@24169.4]
  assign RetimeWrapper_16_io_in = _T_143 & _T_148; // @[package.scala 94:16:@24168.4]
  assign RetimeWrapper_17_clock = clock; // @[:@24174.4]
  assign RetimeWrapper_17_reset = reset; // @[:@24175.4]
  assign RetimeWrapper_17_io_flow = 1'h1; // @[package.scala 95:18:@24177.4]
  assign RetimeWrapper_17_io_in = reset; // @[package.scala 94:16:@24176.4]
  assign RetimeWrapper_18_clock = clock; // @[:@24183.4]
  assign RetimeWrapper_18_reset = reset; // @[:@24184.4]
  assign RetimeWrapper_18_io_flow = 1'h1; // @[package.scala 95:18:@24186.4]
  assign RetimeWrapper_18_io_in = _T_143 & _T_148; // @[package.scala 94:16:@24185.4]
  assign RetimeWrapper_19_clock = clock; // @[:@24191.4]
  assign RetimeWrapper_19_reset = reset; // @[:@24192.4]
  assign RetimeWrapper_19_io_flow = 1'h1; // @[package.scala 95:18:@24194.4]
  assign RetimeWrapper_19_io_in = reset; // @[package.scala 94:16:@24193.4]
  assign RetimeWrapper_20_clock = clock; // @[:@24202.4]
  assign RetimeWrapper_20_reset = reset; // @[:@24203.4]
  assign RetimeWrapper_20_io_flow = 1'h1; // @[package.scala 95:18:@24205.4]
  assign RetimeWrapper_20_io_in = _T_143 & _T_148; // @[package.scala 94:16:@24204.4]
  assign RetimeWrapper_21_clock = clock; // @[:@24210.4]
  assign RetimeWrapper_21_reset = reset; // @[:@24211.4]
  assign RetimeWrapper_21_io_flow = 1'h1; // @[package.scala 95:18:@24213.4]
  assign RetimeWrapper_21_io_in = reset; // @[package.scala 94:16:@24212.4]
  assign RetimeWrapper_22_clock = clock; // @[:@24219.4]
  assign RetimeWrapper_22_reset = reset; // @[:@24220.4]
  assign RetimeWrapper_22_io_flow = 1'h1; // @[package.scala 95:18:@24222.4]
  assign RetimeWrapper_22_io_in = _T_143 & _T_148; // @[package.scala 94:16:@24221.4]
  assign RetimeWrapper_23_clock = clock; // @[:@24227.4]
  assign RetimeWrapper_23_reset = reset; // @[:@24228.4]
  assign RetimeWrapper_23_io_flow = 1'h1; // @[package.scala 95:18:@24230.4]
  assign RetimeWrapper_23_io_in = reset; // @[package.scala 94:16:@24229.4]
  assign NBufCtr_clock = clock; // @[:@24264.4]
  assign NBufCtr_reset = reset; // @[:@24265.4]
  assign NBufCtr_io_input_countUp = 1'h0; // @[NBuffers.scala 43:24:@24272.4]
  assign NBufCtr_io_input_enable = _T_143 & _T_148; // @[NBuffers.scala 42:23:@24271.4]
  assign NBufCtr_1_clock = clock; // @[:@24275.4]
  assign NBufCtr_1_reset = reset; // @[:@24276.4]
  assign NBufCtr_1_io_input_countUp = 1'h0; // @[NBuffers.scala 43:24:@24283.4]
  assign NBufCtr_1_io_input_enable = _T_143 & _T_148; // @[NBuffers.scala 42:23:@24282.4]
  assign statesInR_0_clock = clock; // @[:@24286.4]
  assign statesInR_0_reset = reset; // @[:@24287.4]
  assign statesInR_0_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@24294.4]
  assign statesInR_0_io_input_enable = _T_143 & _T_148; // @[NBuffers.scala 52:23:@24293.4]
  assign statesInR_1_clock = clock; // @[:@24297.4]
  assign statesInR_1_reset = reset; // @[:@24298.4]
  assign statesInR_1_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@24305.4]
  assign statesInR_1_io_input_enable = _T_143 & _T_148; // @[NBuffers.scala 52:23:@24304.4]
  assign statesInR_2_clock = clock; // @[:@24308.4]
  assign statesInR_2_reset = reset; // @[:@24309.4]
  assign statesInR_2_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@24316.4]
  assign statesInR_2_io_input_enable = _T_143 & _T_148; // @[NBuffers.scala 52:23:@24315.4]
  assign statesInR_3_clock = clock; // @[:@24319.4]
  assign statesInR_3_reset = reset; // @[:@24320.4]
  assign statesInR_3_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@24327.4]
  assign statesInR_3_io_input_enable = _T_143 & _T_148; // @[NBuffers.scala 52:23:@24326.4]
  assign statesInR_4_clock = clock; // @[:@24330.4]
  assign statesInR_4_reset = reset; // @[:@24331.4]
  assign statesInR_4_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@24338.4]
  assign statesInR_4_io_input_enable = _T_143 & _T_148; // @[NBuffers.scala 52:23:@24337.4]
  assign statesInR_5_clock = clock; // @[:@24341.4]
  assign statesInR_5_reset = reset; // @[:@24342.4]
  assign statesInR_5_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@24349.4]
  assign statesInR_5_io_input_enable = _T_143 & _T_148; // @[NBuffers.scala 52:23:@24348.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_148 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_148 <= 1'h0;
    end else begin
      _T_148 <= _T_145;
    end
  end
endmodule
module SRAM_10( // @[:@24498.2]
  input         clock, // @[:@24499.4]
  input         reset, // @[:@24500.4]
  input  [1:0]  io_rPort_0_ofs_0, // @[:@24501.4]
  input         io_rPort_0_en_0, // @[:@24501.4]
  input         io_rPort_0_backpressure, // @[:@24501.4]
  output [31:0] io_rPort_0_output_0, // @[:@24501.4]
  input  [1:0]  io_wPort_1_ofs_0, // @[:@24501.4]
  input  [31:0] io_wPort_1_data_0, // @[:@24501.4]
  input         io_wPort_1_en_0, // @[:@24501.4]
  input  [1:0]  io_wPort_0_ofs_0, // @[:@24501.4]
  input  [31:0] io_wPort_0_data_0, // @[:@24501.4]
  input         io_wPort_0_en_0 // @[:@24501.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@24523.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@24523.4]
  wire [1:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@24523.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@24523.4]
  wire [1:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@24523.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@24523.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@24523.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@24523.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@24553.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@24553.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@24567.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@24567.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@24567.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@24567.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@24567.4]
  wire [34:0] _T_106; // @[Cat.scala 30:58:@24542.4]
  wire [34:0] _T_108; // @[Cat.scala 30:58:@24544.4]
  wire [34:0] _T_109; // @[Mux.scala 31:69:@24545.4]
  wire  _T_115; // @[MemPrimitives.scala 126:35:@24557.4]
  wire [3:0] _T_117; // @[Cat.scala 30:58:@24559.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@24523.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@24553.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@24567.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_106 = {io_wPort_0_en_0,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@24542.4]
  assign _T_108 = {io_wPort_1_en_0,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@24544.4]
  assign _T_109 = io_wPort_0_en_0 ? _T_106 : _T_108; // @[Mux.scala 31:69:@24545.4]
  assign _T_115 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@24557.4]
  assign _T_117 = {_T_115,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@24559.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@24574.4]
  assign Mem1D_clock = clock; // @[:@24524.4]
  assign Mem1D_reset = reset; // @[:@24525.4]
  assign Mem1D_io_r_ofs_0 = _T_117[1:0]; // @[MemPrimitives.scala 131:28:@24563.4]
  assign Mem1D_io_r_backpressure = _T_117[2]; // @[MemPrimitives.scala 132:32:@24564.4]
  assign Mem1D_io_w_ofs_0 = _T_109[1:0]; // @[MemPrimitives.scala 94:28:@24549.4]
  assign Mem1D_io_w_data_0 = _T_109[33:2]; // @[MemPrimitives.scala 95:29:@24550.4]
  assign Mem1D_io_w_en_0 = _T_109[34]; // @[MemPrimitives.scala 96:27:@24551.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@24556.4]
  assign RetimeWrapper_clock = clock; // @[:@24568.4]
  assign RetimeWrapper_reset = reset; // @[:@24569.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@24571.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@24570.4]
endmodule
module x554_tmp_0( // @[:@25696.2]
  input         clock, // @[:@25697.4]
  input         reset, // @[:@25698.4]
  input  [1:0]  io_rPort_0_ofs_0, // @[:@25699.4]
  input         io_rPort_0_en_0, // @[:@25699.4]
  output [31:0] io_rPort_0_output_0, // @[:@25699.4]
  input  [1:0]  io_wPort_1_ofs_0, // @[:@25699.4]
  input  [31:0] io_wPort_1_data_0, // @[:@25699.4]
  input         io_wPort_1_en_0, // @[:@25699.4]
  input  [1:0]  io_wPort_0_ofs_0, // @[:@25699.4]
  input  [31:0] io_wPort_0_data_0, // @[:@25699.4]
  input         io_wPort_0_en_0, // @[:@25699.4]
  input         io_sEn_0, // @[:@25699.4]
  input         io_sEn_1, // @[:@25699.4]
  input         io_sEn_2, // @[:@25699.4]
  input         io_sEn_3, // @[:@25699.4]
  input         io_sEn_4, // @[:@25699.4]
  input         io_sEn_5, // @[:@25699.4]
  input         io_sDone_0, // @[:@25699.4]
  input         io_sDone_1, // @[:@25699.4]
  input         io_sDone_2, // @[:@25699.4]
  input         io_sDone_3, // @[:@25699.4]
  input         io_sDone_4, // @[:@25699.4]
  input         io_sDone_5 // @[:@25699.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@25709.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@25709.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@25709.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@25709.4]
  wire  ctrl_io_sEn_2; // @[NBuffers.scala 83:20:@25709.4]
  wire  ctrl_io_sEn_3; // @[NBuffers.scala 83:20:@25709.4]
  wire  ctrl_io_sEn_4; // @[NBuffers.scala 83:20:@25709.4]
  wire  ctrl_io_sEn_5; // @[NBuffers.scala 83:20:@25709.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@25709.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@25709.4]
  wire  ctrl_io_sDone_2; // @[NBuffers.scala 83:20:@25709.4]
  wire  ctrl_io_sDone_3; // @[NBuffers.scala 83:20:@25709.4]
  wire  ctrl_io_sDone_4; // @[NBuffers.scala 83:20:@25709.4]
  wire  ctrl_io_sDone_5; // @[NBuffers.scala 83:20:@25709.4]
  wire [3:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@25709.4]
  wire [3:0] ctrl_io_statesInW_1; // @[NBuffers.scala 83:20:@25709.4]
  wire [3:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@25709.4]
  wire [3:0] ctrl_io_statesInR_5; // @[NBuffers.scala 83:20:@25709.4]
  wire  SRAM_clock; // @[NBuffers.scala 94:23:@25724.4]
  wire  SRAM_reset; // @[NBuffers.scala 94:23:@25724.4]
  wire [1:0] SRAM_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@25724.4]
  wire  SRAM_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@25724.4]
  wire  SRAM_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@25724.4]
  wire [31:0] SRAM_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@25724.4]
  wire [1:0] SRAM_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@25724.4]
  wire [31:0] SRAM_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@25724.4]
  wire  SRAM_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@25724.4]
  wire [1:0] SRAM_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@25724.4]
  wire [31:0] SRAM_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@25724.4]
  wire  SRAM_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@25724.4]
  wire  SRAM_1_clock; // @[NBuffers.scala 94:23:@25747.4]
  wire  SRAM_1_reset; // @[NBuffers.scala 94:23:@25747.4]
  wire [1:0] SRAM_1_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@25747.4]
  wire  SRAM_1_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@25747.4]
  wire  SRAM_1_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@25747.4]
  wire [31:0] SRAM_1_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@25747.4]
  wire [1:0] SRAM_1_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@25747.4]
  wire [31:0] SRAM_1_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@25747.4]
  wire  SRAM_1_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@25747.4]
  wire [1:0] SRAM_1_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@25747.4]
  wire [31:0] SRAM_1_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@25747.4]
  wire  SRAM_1_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@25747.4]
  wire  SRAM_2_clock; // @[NBuffers.scala 94:23:@25770.4]
  wire  SRAM_2_reset; // @[NBuffers.scala 94:23:@25770.4]
  wire [1:0] SRAM_2_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@25770.4]
  wire  SRAM_2_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@25770.4]
  wire  SRAM_2_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@25770.4]
  wire [31:0] SRAM_2_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@25770.4]
  wire [1:0] SRAM_2_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@25770.4]
  wire [31:0] SRAM_2_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@25770.4]
  wire  SRAM_2_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@25770.4]
  wire [1:0] SRAM_2_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@25770.4]
  wire [31:0] SRAM_2_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@25770.4]
  wire  SRAM_2_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@25770.4]
  wire  SRAM_3_clock; // @[NBuffers.scala 94:23:@25793.4]
  wire  SRAM_3_reset; // @[NBuffers.scala 94:23:@25793.4]
  wire [1:0] SRAM_3_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@25793.4]
  wire  SRAM_3_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@25793.4]
  wire  SRAM_3_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@25793.4]
  wire [31:0] SRAM_3_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@25793.4]
  wire [1:0] SRAM_3_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@25793.4]
  wire [31:0] SRAM_3_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@25793.4]
  wire  SRAM_3_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@25793.4]
  wire [1:0] SRAM_3_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@25793.4]
  wire [31:0] SRAM_3_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@25793.4]
  wire  SRAM_3_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@25793.4]
  wire  SRAM_4_clock; // @[NBuffers.scala 94:23:@25816.4]
  wire  SRAM_4_reset; // @[NBuffers.scala 94:23:@25816.4]
  wire [1:0] SRAM_4_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@25816.4]
  wire  SRAM_4_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@25816.4]
  wire  SRAM_4_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@25816.4]
  wire [31:0] SRAM_4_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@25816.4]
  wire [1:0] SRAM_4_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@25816.4]
  wire [31:0] SRAM_4_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@25816.4]
  wire  SRAM_4_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@25816.4]
  wire [1:0] SRAM_4_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@25816.4]
  wire [31:0] SRAM_4_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@25816.4]
  wire  SRAM_4_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@25816.4]
  wire  SRAM_5_clock; // @[NBuffers.scala 94:23:@25839.4]
  wire  SRAM_5_reset; // @[NBuffers.scala 94:23:@25839.4]
  wire [1:0] SRAM_5_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@25839.4]
  wire  SRAM_5_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@25839.4]
  wire  SRAM_5_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@25839.4]
  wire [31:0] SRAM_5_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@25839.4]
  wire [1:0] SRAM_5_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@25839.4]
  wire [31:0] SRAM_5_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@25839.4]
  wire  SRAM_5_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@25839.4]
  wire [1:0] SRAM_5_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@25839.4]
  wire [31:0] SRAM_5_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@25839.4]
  wire  SRAM_5_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@25839.4]
  wire  _T_148; // @[NBuffers.scala 104:105:@25862.4]
  wire  _T_152; // @[NBuffers.scala 104:105:@25872.4]
  wire  _T_156; // @[NBuffers.scala 108:92:@25882.4]
  wire  _T_159; // @[NBuffers.scala 104:105:@25888.4]
  wire  _T_163; // @[NBuffers.scala 104:105:@25898.4]
  wire  _T_167; // @[NBuffers.scala 108:92:@25908.4]
  wire  _T_170; // @[NBuffers.scala 104:105:@25914.4]
  wire  _T_174; // @[NBuffers.scala 104:105:@25924.4]
  wire  _T_178; // @[NBuffers.scala 108:92:@25934.4]
  wire  _T_181; // @[NBuffers.scala 104:105:@25940.4]
  wire  _T_185; // @[NBuffers.scala 104:105:@25950.4]
  wire  _T_189; // @[NBuffers.scala 108:92:@25960.4]
  wire  _T_192; // @[NBuffers.scala 104:105:@25966.4]
  wire  _T_196; // @[NBuffers.scala 104:105:@25976.4]
  wire  _T_200; // @[NBuffers.scala 108:92:@25986.4]
  wire  _T_203; // @[NBuffers.scala 104:105:@25992.4]
  wire  _T_207; // @[NBuffers.scala 104:105:@26002.4]
  wire  _T_211; // @[NBuffers.scala 108:92:@26012.4]
  wire [31:0] _T_227; // @[Mux.scala 19:72:@26024.4]
  wire [31:0] _T_229; // @[Mux.scala 19:72:@26025.4]
  wire [31:0] _T_231; // @[Mux.scala 19:72:@26026.4]
  wire [31:0] _T_233; // @[Mux.scala 19:72:@26027.4]
  wire [31:0] _T_235; // @[Mux.scala 19:72:@26028.4]
  wire [31:0] _T_237; // @[Mux.scala 19:72:@26029.4]
  wire [31:0] _T_238; // @[Mux.scala 19:72:@26030.4]
  wire [31:0] _T_239; // @[Mux.scala 19:72:@26031.4]
  wire [31:0] _T_240; // @[Mux.scala 19:72:@26032.4]
  wire [31:0] _T_241; // @[Mux.scala 19:72:@26033.4]
  NBufController_5 ctrl ( // @[NBuffers.scala 83:20:@25709.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sEn_2(ctrl_io_sEn_2),
    .io_sEn_3(ctrl_io_sEn_3),
    .io_sEn_4(ctrl_io_sEn_4),
    .io_sEn_5(ctrl_io_sEn_5),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_sDone_2(ctrl_io_sDone_2),
    .io_sDone_3(ctrl_io_sDone_3),
    .io_sDone_4(ctrl_io_sDone_4),
    .io_sDone_5(ctrl_io_sDone_5),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInW_1(ctrl_io_statesInW_1),
    .io_statesInR_1(ctrl_io_statesInR_1),
    .io_statesInR_5(ctrl_io_statesInR_5)
  );
  SRAM_10 SRAM ( // @[NBuffers.scala 94:23:@25724.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_rPort_0_ofs_0(SRAM_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_1 ( // @[NBuffers.scala 94:23:@25747.4]
    .clock(SRAM_1_clock),
    .reset(SRAM_1_reset),
    .io_rPort_0_ofs_0(SRAM_1_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_1_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_1_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_1_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_1_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_1_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_1_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_1_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_1_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_2 ( // @[NBuffers.scala 94:23:@25770.4]
    .clock(SRAM_2_clock),
    .reset(SRAM_2_reset),
    .io_rPort_0_ofs_0(SRAM_2_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_2_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_2_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_2_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_2_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_2_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_2_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_2_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_2_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_2_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_3 ( // @[NBuffers.scala 94:23:@25793.4]
    .clock(SRAM_3_clock),
    .reset(SRAM_3_reset),
    .io_rPort_0_ofs_0(SRAM_3_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_3_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_3_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_3_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_3_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_3_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_3_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_3_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_3_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_3_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_4 ( // @[NBuffers.scala 94:23:@25816.4]
    .clock(SRAM_4_clock),
    .reset(SRAM_4_reset),
    .io_rPort_0_ofs_0(SRAM_4_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_4_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_4_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_4_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_4_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_4_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_4_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_4_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_4_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_4_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_5 ( // @[NBuffers.scala 94:23:@25839.4]
    .clock(SRAM_5_clock),
    .reset(SRAM_5_reset),
    .io_rPort_0_ofs_0(SRAM_5_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_5_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_5_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_5_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_5_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_5_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_5_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_5_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_5_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_5_io_wPort_0_en_0)
  );
  assign _T_148 = ctrl_io_statesInW_0 == 4'h0; // @[NBuffers.scala 104:105:@25862.4]
  assign _T_152 = ctrl_io_statesInW_1 == 4'h0; // @[NBuffers.scala 104:105:@25872.4]
  assign _T_156 = ctrl_io_statesInR_1 == 4'h0; // @[NBuffers.scala 108:92:@25882.4]
  assign _T_159 = ctrl_io_statesInW_0 == 4'h1; // @[NBuffers.scala 104:105:@25888.4]
  assign _T_163 = ctrl_io_statesInW_1 == 4'h1; // @[NBuffers.scala 104:105:@25898.4]
  assign _T_167 = ctrl_io_statesInR_1 == 4'h1; // @[NBuffers.scala 108:92:@25908.4]
  assign _T_170 = ctrl_io_statesInW_0 == 4'h2; // @[NBuffers.scala 104:105:@25914.4]
  assign _T_174 = ctrl_io_statesInW_1 == 4'h2; // @[NBuffers.scala 104:105:@25924.4]
  assign _T_178 = ctrl_io_statesInR_1 == 4'h2; // @[NBuffers.scala 108:92:@25934.4]
  assign _T_181 = ctrl_io_statesInW_0 == 4'h3; // @[NBuffers.scala 104:105:@25940.4]
  assign _T_185 = ctrl_io_statesInW_1 == 4'h3; // @[NBuffers.scala 104:105:@25950.4]
  assign _T_189 = ctrl_io_statesInR_1 == 4'h3; // @[NBuffers.scala 108:92:@25960.4]
  assign _T_192 = ctrl_io_statesInW_0 == 4'h4; // @[NBuffers.scala 104:105:@25966.4]
  assign _T_196 = ctrl_io_statesInW_1 == 4'h4; // @[NBuffers.scala 104:105:@25976.4]
  assign _T_200 = ctrl_io_statesInR_1 == 4'h4; // @[NBuffers.scala 108:92:@25986.4]
  assign _T_203 = ctrl_io_statesInW_0 == 4'h5; // @[NBuffers.scala 104:105:@25992.4]
  assign _T_207 = ctrl_io_statesInW_1 == 4'h5; // @[NBuffers.scala 104:105:@26002.4]
  assign _T_211 = ctrl_io_statesInR_1 == 4'h5; // @[NBuffers.scala 108:92:@26012.4]
  assign _T_227 = _T_156 ? SRAM_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@26024.4]
  assign _T_229 = _T_167 ? SRAM_1_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@26025.4]
  assign _T_231 = _T_178 ? SRAM_2_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@26026.4]
  assign _T_233 = _T_189 ? SRAM_3_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@26027.4]
  assign _T_235 = _T_200 ? SRAM_4_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@26028.4]
  assign _T_237 = _T_211 ? SRAM_5_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@26029.4]
  assign _T_238 = _T_227 | _T_229; // @[Mux.scala 19:72:@26030.4]
  assign _T_239 = _T_238 | _T_231; // @[Mux.scala 19:72:@26031.4]
  assign _T_240 = _T_239 | _T_233; // @[Mux.scala 19:72:@26032.4]
  assign _T_241 = _T_240 | _T_235; // @[Mux.scala 19:72:@26033.4]
  assign io_rPort_0_output_0 = _T_241 | _T_237; // @[NBuffers.scala 115:66:@26037.4]
  assign ctrl_clock = clock; // @[:@25710.4]
  assign ctrl_reset = reset; // @[:@25711.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@25712.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@25714.4]
  assign ctrl_io_sEn_2 = io_sEn_2; // @[NBuffers.scala 85:20:@25716.4]
  assign ctrl_io_sEn_3 = io_sEn_3; // @[NBuffers.scala 85:20:@25718.4]
  assign ctrl_io_sEn_4 = io_sEn_4; // @[NBuffers.scala 85:20:@25720.4]
  assign ctrl_io_sEn_5 = io_sEn_5; // @[NBuffers.scala 85:20:@25722.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@25713.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@25715.4]
  assign ctrl_io_sDone_2 = io_sDone_2; // @[NBuffers.scala 86:22:@25717.4]
  assign ctrl_io_sDone_3 = io_sDone_3; // @[NBuffers.scala 86:22:@25719.4]
  assign ctrl_io_sDone_4 = io_sDone_4; // @[NBuffers.scala 86:22:@25721.4]
  assign ctrl_io_sDone_5 = io_sDone_5; // @[NBuffers.scala 86:22:@25723.4]
  assign SRAM_clock = clock; // @[:@25725.4]
  assign SRAM_reset = reset; // @[:@25726.4]
  assign SRAM_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@25884.4]
  assign SRAM_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_156; // @[MemPrimitives.scala 43:33:@25886.4]
  assign SRAM_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@25887.4]
  assign SRAM_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@25874.4]
  assign SRAM_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@25875.4]
  assign SRAM_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_152; // @[MemPrimitives.scala 37:29:@25881.4]
  assign SRAM_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@25864.4]
  assign SRAM_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@25865.4]
  assign SRAM_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_148; // @[MemPrimitives.scala 37:29:@25871.4]
  assign SRAM_1_clock = clock; // @[:@25748.4]
  assign SRAM_1_reset = reset; // @[:@25749.4]
  assign SRAM_1_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@25910.4]
  assign SRAM_1_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_167; // @[MemPrimitives.scala 43:33:@25912.4]
  assign SRAM_1_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@25913.4]
  assign SRAM_1_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@25900.4]
  assign SRAM_1_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@25901.4]
  assign SRAM_1_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_163; // @[MemPrimitives.scala 37:29:@25907.4]
  assign SRAM_1_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@25890.4]
  assign SRAM_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@25891.4]
  assign SRAM_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_159; // @[MemPrimitives.scala 37:29:@25897.4]
  assign SRAM_2_clock = clock; // @[:@25771.4]
  assign SRAM_2_reset = reset; // @[:@25772.4]
  assign SRAM_2_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@25936.4]
  assign SRAM_2_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_178; // @[MemPrimitives.scala 43:33:@25938.4]
  assign SRAM_2_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@25939.4]
  assign SRAM_2_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@25926.4]
  assign SRAM_2_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@25927.4]
  assign SRAM_2_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_174; // @[MemPrimitives.scala 37:29:@25933.4]
  assign SRAM_2_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@25916.4]
  assign SRAM_2_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@25917.4]
  assign SRAM_2_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_170; // @[MemPrimitives.scala 37:29:@25923.4]
  assign SRAM_3_clock = clock; // @[:@25794.4]
  assign SRAM_3_reset = reset; // @[:@25795.4]
  assign SRAM_3_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@25962.4]
  assign SRAM_3_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_189; // @[MemPrimitives.scala 43:33:@25964.4]
  assign SRAM_3_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@25965.4]
  assign SRAM_3_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@25952.4]
  assign SRAM_3_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@25953.4]
  assign SRAM_3_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_185; // @[MemPrimitives.scala 37:29:@25959.4]
  assign SRAM_3_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@25942.4]
  assign SRAM_3_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@25943.4]
  assign SRAM_3_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_181; // @[MemPrimitives.scala 37:29:@25949.4]
  assign SRAM_4_clock = clock; // @[:@25817.4]
  assign SRAM_4_reset = reset; // @[:@25818.4]
  assign SRAM_4_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@25988.4]
  assign SRAM_4_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_200; // @[MemPrimitives.scala 43:33:@25990.4]
  assign SRAM_4_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@25991.4]
  assign SRAM_4_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@25978.4]
  assign SRAM_4_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@25979.4]
  assign SRAM_4_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_196; // @[MemPrimitives.scala 37:29:@25985.4]
  assign SRAM_4_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@25968.4]
  assign SRAM_4_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@25969.4]
  assign SRAM_4_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_192; // @[MemPrimitives.scala 37:29:@25975.4]
  assign SRAM_5_clock = clock; // @[:@25840.4]
  assign SRAM_5_reset = reset; // @[:@25841.4]
  assign SRAM_5_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@26014.4]
  assign SRAM_5_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_211; // @[MemPrimitives.scala 43:33:@26016.4]
  assign SRAM_5_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@26017.4]
  assign SRAM_5_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@26004.4]
  assign SRAM_5_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@26005.4]
  assign SRAM_5_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_207; // @[MemPrimitives.scala 37:29:@26011.4]
  assign SRAM_5_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@25994.4]
  assign SRAM_5_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@25995.4]
  assign SRAM_5_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_203; // @[MemPrimitives.scala 37:29:@26001.4]
endmodule
module x557_tmp_3( // @[:@36625.2]
  input         clock, // @[:@36626.4]
  input         reset, // @[:@36627.4]
  input  [1:0]  io_rPort_0_ofs_0, // @[:@36628.4]
  input         io_rPort_0_en_0, // @[:@36628.4]
  output [31:0] io_rPort_0_output_0, // @[:@36628.4]
  input  [1:0]  io_wPort_1_ofs_0, // @[:@36628.4]
  input  [31:0] io_wPort_1_data_0, // @[:@36628.4]
  input         io_wPort_1_en_0, // @[:@36628.4]
  input  [1:0]  io_wPort_0_ofs_0, // @[:@36628.4]
  input  [31:0] io_wPort_0_data_0, // @[:@36628.4]
  input         io_wPort_0_en_0, // @[:@36628.4]
  input         io_sEn_0, // @[:@36628.4]
  input         io_sEn_1, // @[:@36628.4]
  input         io_sEn_2, // @[:@36628.4]
  input         io_sEn_3, // @[:@36628.4]
  input         io_sEn_4, // @[:@36628.4]
  input         io_sEn_5, // @[:@36628.4]
  input         io_sDone_0, // @[:@36628.4]
  input         io_sDone_1, // @[:@36628.4]
  input         io_sDone_2, // @[:@36628.4]
  input         io_sDone_3, // @[:@36628.4]
  input         io_sDone_4, // @[:@36628.4]
  input         io_sDone_5 // @[:@36628.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@36638.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@36638.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@36638.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@36638.4]
  wire  ctrl_io_sEn_2; // @[NBuffers.scala 83:20:@36638.4]
  wire  ctrl_io_sEn_3; // @[NBuffers.scala 83:20:@36638.4]
  wire  ctrl_io_sEn_4; // @[NBuffers.scala 83:20:@36638.4]
  wire  ctrl_io_sEn_5; // @[NBuffers.scala 83:20:@36638.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@36638.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@36638.4]
  wire  ctrl_io_sDone_2; // @[NBuffers.scala 83:20:@36638.4]
  wire  ctrl_io_sDone_3; // @[NBuffers.scala 83:20:@36638.4]
  wire  ctrl_io_sDone_4; // @[NBuffers.scala 83:20:@36638.4]
  wire  ctrl_io_sDone_5; // @[NBuffers.scala 83:20:@36638.4]
  wire [3:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@36638.4]
  wire [3:0] ctrl_io_statesInW_1; // @[NBuffers.scala 83:20:@36638.4]
  wire [3:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@36638.4]
  wire [3:0] ctrl_io_statesInR_5; // @[NBuffers.scala 83:20:@36638.4]
  wire  SRAM_clock; // @[NBuffers.scala 94:23:@36653.4]
  wire  SRAM_reset; // @[NBuffers.scala 94:23:@36653.4]
  wire [1:0] SRAM_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@36653.4]
  wire  SRAM_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@36653.4]
  wire  SRAM_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@36653.4]
  wire [31:0] SRAM_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@36653.4]
  wire [1:0] SRAM_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@36653.4]
  wire [31:0] SRAM_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@36653.4]
  wire  SRAM_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@36653.4]
  wire [1:0] SRAM_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@36653.4]
  wire [31:0] SRAM_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@36653.4]
  wire  SRAM_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@36653.4]
  wire  SRAM_1_clock; // @[NBuffers.scala 94:23:@36676.4]
  wire  SRAM_1_reset; // @[NBuffers.scala 94:23:@36676.4]
  wire [1:0] SRAM_1_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@36676.4]
  wire  SRAM_1_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@36676.4]
  wire  SRAM_1_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@36676.4]
  wire [31:0] SRAM_1_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@36676.4]
  wire [1:0] SRAM_1_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@36676.4]
  wire [31:0] SRAM_1_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@36676.4]
  wire  SRAM_1_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@36676.4]
  wire [1:0] SRAM_1_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@36676.4]
  wire [31:0] SRAM_1_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@36676.4]
  wire  SRAM_1_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@36676.4]
  wire  SRAM_2_clock; // @[NBuffers.scala 94:23:@36699.4]
  wire  SRAM_2_reset; // @[NBuffers.scala 94:23:@36699.4]
  wire [1:0] SRAM_2_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@36699.4]
  wire  SRAM_2_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@36699.4]
  wire  SRAM_2_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@36699.4]
  wire [31:0] SRAM_2_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@36699.4]
  wire [1:0] SRAM_2_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@36699.4]
  wire [31:0] SRAM_2_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@36699.4]
  wire  SRAM_2_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@36699.4]
  wire [1:0] SRAM_2_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@36699.4]
  wire [31:0] SRAM_2_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@36699.4]
  wire  SRAM_2_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@36699.4]
  wire  SRAM_3_clock; // @[NBuffers.scala 94:23:@36722.4]
  wire  SRAM_3_reset; // @[NBuffers.scala 94:23:@36722.4]
  wire [1:0] SRAM_3_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@36722.4]
  wire  SRAM_3_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@36722.4]
  wire  SRAM_3_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@36722.4]
  wire [31:0] SRAM_3_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@36722.4]
  wire [1:0] SRAM_3_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@36722.4]
  wire [31:0] SRAM_3_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@36722.4]
  wire  SRAM_3_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@36722.4]
  wire [1:0] SRAM_3_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@36722.4]
  wire [31:0] SRAM_3_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@36722.4]
  wire  SRAM_3_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@36722.4]
  wire  SRAM_4_clock; // @[NBuffers.scala 94:23:@36745.4]
  wire  SRAM_4_reset; // @[NBuffers.scala 94:23:@36745.4]
  wire [1:0] SRAM_4_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@36745.4]
  wire  SRAM_4_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@36745.4]
  wire  SRAM_4_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@36745.4]
  wire [31:0] SRAM_4_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@36745.4]
  wire [1:0] SRAM_4_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@36745.4]
  wire [31:0] SRAM_4_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@36745.4]
  wire  SRAM_4_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@36745.4]
  wire [1:0] SRAM_4_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@36745.4]
  wire [31:0] SRAM_4_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@36745.4]
  wire  SRAM_4_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@36745.4]
  wire  SRAM_5_clock; // @[NBuffers.scala 94:23:@36768.4]
  wire  SRAM_5_reset; // @[NBuffers.scala 94:23:@36768.4]
  wire [1:0] SRAM_5_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@36768.4]
  wire  SRAM_5_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@36768.4]
  wire  SRAM_5_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@36768.4]
  wire [31:0] SRAM_5_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@36768.4]
  wire [1:0] SRAM_5_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@36768.4]
  wire [31:0] SRAM_5_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@36768.4]
  wire  SRAM_5_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@36768.4]
  wire [1:0] SRAM_5_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@36768.4]
  wire [31:0] SRAM_5_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@36768.4]
  wire  SRAM_5_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@36768.4]
  wire  _T_148; // @[NBuffers.scala 104:105:@36791.4]
  wire  _T_152; // @[NBuffers.scala 104:105:@36801.4]
  wire  _T_156; // @[NBuffers.scala 108:92:@36811.4]
  wire  _T_159; // @[NBuffers.scala 104:105:@36817.4]
  wire  _T_163; // @[NBuffers.scala 104:105:@36827.4]
  wire  _T_167; // @[NBuffers.scala 108:92:@36837.4]
  wire  _T_170; // @[NBuffers.scala 104:105:@36843.4]
  wire  _T_174; // @[NBuffers.scala 104:105:@36853.4]
  wire  _T_178; // @[NBuffers.scala 108:92:@36863.4]
  wire  _T_181; // @[NBuffers.scala 104:105:@36869.4]
  wire  _T_185; // @[NBuffers.scala 104:105:@36879.4]
  wire  _T_189; // @[NBuffers.scala 108:92:@36889.4]
  wire  _T_192; // @[NBuffers.scala 104:105:@36895.4]
  wire  _T_196; // @[NBuffers.scala 104:105:@36905.4]
  wire  _T_200; // @[NBuffers.scala 108:92:@36915.4]
  wire  _T_203; // @[NBuffers.scala 104:105:@36921.4]
  wire  _T_207; // @[NBuffers.scala 104:105:@36931.4]
  wire  _T_211; // @[NBuffers.scala 108:92:@36941.4]
  wire [31:0] _T_227; // @[Mux.scala 19:72:@36953.4]
  wire [31:0] _T_229; // @[Mux.scala 19:72:@36954.4]
  wire [31:0] _T_231; // @[Mux.scala 19:72:@36955.4]
  wire [31:0] _T_233; // @[Mux.scala 19:72:@36956.4]
  wire [31:0] _T_235; // @[Mux.scala 19:72:@36957.4]
  wire [31:0] _T_237; // @[Mux.scala 19:72:@36958.4]
  wire [31:0] _T_238; // @[Mux.scala 19:72:@36959.4]
  wire [31:0] _T_239; // @[Mux.scala 19:72:@36960.4]
  wire [31:0] _T_240; // @[Mux.scala 19:72:@36961.4]
  wire [31:0] _T_241; // @[Mux.scala 19:72:@36962.4]
  NBufController_5 ctrl ( // @[NBuffers.scala 83:20:@36638.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sEn_2(ctrl_io_sEn_2),
    .io_sEn_3(ctrl_io_sEn_3),
    .io_sEn_4(ctrl_io_sEn_4),
    .io_sEn_5(ctrl_io_sEn_5),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_sDone_2(ctrl_io_sDone_2),
    .io_sDone_3(ctrl_io_sDone_3),
    .io_sDone_4(ctrl_io_sDone_4),
    .io_sDone_5(ctrl_io_sDone_5),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInW_1(ctrl_io_statesInW_1),
    .io_statesInR_1(ctrl_io_statesInR_1),
    .io_statesInR_5(ctrl_io_statesInR_5)
  );
  SRAM_10 SRAM ( // @[NBuffers.scala 94:23:@36653.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_rPort_0_ofs_0(SRAM_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_1 ( // @[NBuffers.scala 94:23:@36676.4]
    .clock(SRAM_1_clock),
    .reset(SRAM_1_reset),
    .io_rPort_0_ofs_0(SRAM_1_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_1_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_1_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_1_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_1_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_1_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_1_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_1_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_1_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_2 ( // @[NBuffers.scala 94:23:@36699.4]
    .clock(SRAM_2_clock),
    .reset(SRAM_2_reset),
    .io_rPort_0_ofs_0(SRAM_2_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_2_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_2_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_2_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_2_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_2_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_2_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_2_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_2_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_2_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_3 ( // @[NBuffers.scala 94:23:@36722.4]
    .clock(SRAM_3_clock),
    .reset(SRAM_3_reset),
    .io_rPort_0_ofs_0(SRAM_3_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_3_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_3_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_3_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_3_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_3_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_3_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_3_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_3_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_3_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_4 ( // @[NBuffers.scala 94:23:@36745.4]
    .clock(SRAM_4_clock),
    .reset(SRAM_4_reset),
    .io_rPort_0_ofs_0(SRAM_4_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_4_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_4_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_4_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_4_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_4_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_4_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_4_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_4_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_4_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_5 ( // @[NBuffers.scala 94:23:@36768.4]
    .clock(SRAM_5_clock),
    .reset(SRAM_5_reset),
    .io_rPort_0_ofs_0(SRAM_5_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_5_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_5_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_5_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_5_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_5_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_5_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_5_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_5_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_5_io_wPort_0_en_0)
  );
  assign _T_148 = ctrl_io_statesInW_0 == 4'h0; // @[NBuffers.scala 104:105:@36791.4]
  assign _T_152 = ctrl_io_statesInW_1 == 4'h0; // @[NBuffers.scala 104:105:@36801.4]
  assign _T_156 = ctrl_io_statesInR_5 == 4'h0; // @[NBuffers.scala 108:92:@36811.4]
  assign _T_159 = ctrl_io_statesInW_0 == 4'h1; // @[NBuffers.scala 104:105:@36817.4]
  assign _T_163 = ctrl_io_statesInW_1 == 4'h1; // @[NBuffers.scala 104:105:@36827.4]
  assign _T_167 = ctrl_io_statesInR_5 == 4'h1; // @[NBuffers.scala 108:92:@36837.4]
  assign _T_170 = ctrl_io_statesInW_0 == 4'h2; // @[NBuffers.scala 104:105:@36843.4]
  assign _T_174 = ctrl_io_statesInW_1 == 4'h2; // @[NBuffers.scala 104:105:@36853.4]
  assign _T_178 = ctrl_io_statesInR_5 == 4'h2; // @[NBuffers.scala 108:92:@36863.4]
  assign _T_181 = ctrl_io_statesInW_0 == 4'h3; // @[NBuffers.scala 104:105:@36869.4]
  assign _T_185 = ctrl_io_statesInW_1 == 4'h3; // @[NBuffers.scala 104:105:@36879.4]
  assign _T_189 = ctrl_io_statesInR_5 == 4'h3; // @[NBuffers.scala 108:92:@36889.4]
  assign _T_192 = ctrl_io_statesInW_0 == 4'h4; // @[NBuffers.scala 104:105:@36895.4]
  assign _T_196 = ctrl_io_statesInW_1 == 4'h4; // @[NBuffers.scala 104:105:@36905.4]
  assign _T_200 = ctrl_io_statesInR_5 == 4'h4; // @[NBuffers.scala 108:92:@36915.4]
  assign _T_203 = ctrl_io_statesInW_0 == 4'h5; // @[NBuffers.scala 104:105:@36921.4]
  assign _T_207 = ctrl_io_statesInW_1 == 4'h5; // @[NBuffers.scala 104:105:@36931.4]
  assign _T_211 = ctrl_io_statesInR_5 == 4'h5; // @[NBuffers.scala 108:92:@36941.4]
  assign _T_227 = _T_156 ? SRAM_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@36953.4]
  assign _T_229 = _T_167 ? SRAM_1_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@36954.4]
  assign _T_231 = _T_178 ? SRAM_2_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@36955.4]
  assign _T_233 = _T_189 ? SRAM_3_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@36956.4]
  assign _T_235 = _T_200 ? SRAM_4_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@36957.4]
  assign _T_237 = _T_211 ? SRAM_5_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@36958.4]
  assign _T_238 = _T_227 | _T_229; // @[Mux.scala 19:72:@36959.4]
  assign _T_239 = _T_238 | _T_231; // @[Mux.scala 19:72:@36960.4]
  assign _T_240 = _T_239 | _T_233; // @[Mux.scala 19:72:@36961.4]
  assign _T_241 = _T_240 | _T_235; // @[Mux.scala 19:72:@36962.4]
  assign io_rPort_0_output_0 = _T_241 | _T_237; // @[NBuffers.scala 115:66:@36966.4]
  assign ctrl_clock = clock; // @[:@36639.4]
  assign ctrl_reset = reset; // @[:@36640.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@36641.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@36643.4]
  assign ctrl_io_sEn_2 = io_sEn_2; // @[NBuffers.scala 85:20:@36645.4]
  assign ctrl_io_sEn_3 = io_sEn_3; // @[NBuffers.scala 85:20:@36647.4]
  assign ctrl_io_sEn_4 = io_sEn_4; // @[NBuffers.scala 85:20:@36649.4]
  assign ctrl_io_sEn_5 = io_sEn_5; // @[NBuffers.scala 85:20:@36651.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@36642.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@36644.4]
  assign ctrl_io_sDone_2 = io_sDone_2; // @[NBuffers.scala 86:22:@36646.4]
  assign ctrl_io_sDone_3 = io_sDone_3; // @[NBuffers.scala 86:22:@36648.4]
  assign ctrl_io_sDone_4 = io_sDone_4; // @[NBuffers.scala 86:22:@36650.4]
  assign ctrl_io_sDone_5 = io_sDone_5; // @[NBuffers.scala 86:22:@36652.4]
  assign SRAM_clock = clock; // @[:@36654.4]
  assign SRAM_reset = reset; // @[:@36655.4]
  assign SRAM_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@36813.4]
  assign SRAM_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_156; // @[MemPrimitives.scala 43:33:@36815.4]
  assign SRAM_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@36816.4]
  assign SRAM_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@36803.4]
  assign SRAM_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@36804.4]
  assign SRAM_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_152; // @[MemPrimitives.scala 37:29:@36810.4]
  assign SRAM_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@36793.4]
  assign SRAM_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@36794.4]
  assign SRAM_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_148; // @[MemPrimitives.scala 37:29:@36800.4]
  assign SRAM_1_clock = clock; // @[:@36677.4]
  assign SRAM_1_reset = reset; // @[:@36678.4]
  assign SRAM_1_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@36839.4]
  assign SRAM_1_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_167; // @[MemPrimitives.scala 43:33:@36841.4]
  assign SRAM_1_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@36842.4]
  assign SRAM_1_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@36829.4]
  assign SRAM_1_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@36830.4]
  assign SRAM_1_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_163; // @[MemPrimitives.scala 37:29:@36836.4]
  assign SRAM_1_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@36819.4]
  assign SRAM_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@36820.4]
  assign SRAM_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_159; // @[MemPrimitives.scala 37:29:@36826.4]
  assign SRAM_2_clock = clock; // @[:@36700.4]
  assign SRAM_2_reset = reset; // @[:@36701.4]
  assign SRAM_2_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@36865.4]
  assign SRAM_2_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_178; // @[MemPrimitives.scala 43:33:@36867.4]
  assign SRAM_2_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@36868.4]
  assign SRAM_2_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@36855.4]
  assign SRAM_2_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@36856.4]
  assign SRAM_2_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_174; // @[MemPrimitives.scala 37:29:@36862.4]
  assign SRAM_2_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@36845.4]
  assign SRAM_2_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@36846.4]
  assign SRAM_2_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_170; // @[MemPrimitives.scala 37:29:@36852.4]
  assign SRAM_3_clock = clock; // @[:@36723.4]
  assign SRAM_3_reset = reset; // @[:@36724.4]
  assign SRAM_3_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@36891.4]
  assign SRAM_3_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_189; // @[MemPrimitives.scala 43:33:@36893.4]
  assign SRAM_3_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@36894.4]
  assign SRAM_3_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@36881.4]
  assign SRAM_3_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@36882.4]
  assign SRAM_3_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_185; // @[MemPrimitives.scala 37:29:@36888.4]
  assign SRAM_3_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@36871.4]
  assign SRAM_3_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@36872.4]
  assign SRAM_3_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_181; // @[MemPrimitives.scala 37:29:@36878.4]
  assign SRAM_4_clock = clock; // @[:@36746.4]
  assign SRAM_4_reset = reset; // @[:@36747.4]
  assign SRAM_4_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@36917.4]
  assign SRAM_4_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_200; // @[MemPrimitives.scala 43:33:@36919.4]
  assign SRAM_4_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@36920.4]
  assign SRAM_4_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@36907.4]
  assign SRAM_4_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@36908.4]
  assign SRAM_4_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_196; // @[MemPrimitives.scala 37:29:@36914.4]
  assign SRAM_4_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@36897.4]
  assign SRAM_4_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@36898.4]
  assign SRAM_4_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_192; // @[MemPrimitives.scala 37:29:@36904.4]
  assign SRAM_5_clock = clock; // @[:@36769.4]
  assign SRAM_5_reset = reset; // @[:@36770.4]
  assign SRAM_5_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@36943.4]
  assign SRAM_5_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_211; // @[MemPrimitives.scala 43:33:@36945.4]
  assign SRAM_5_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@36946.4]
  assign SRAM_5_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@36933.4]
  assign SRAM_5_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@36934.4]
  assign SRAM_5_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_207; // @[MemPrimitives.scala 37:29:@36940.4]
  assign SRAM_5_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@36923.4]
  assign SRAM_5_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@36924.4]
  assign SRAM_5_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_203; // @[MemPrimitives.scala 37:29:@36930.4]
endmodule
module NBufController_9( // @[:@38784.2]
  input        clock, // @[:@38785.4]
  input        reset, // @[:@38786.4]
  input        io_sEn_0, // @[:@38787.4]
  input        io_sEn_1, // @[:@38787.4]
  input        io_sEn_2, // @[:@38787.4]
  input        io_sEn_3, // @[:@38787.4]
  input        io_sEn_4, // @[:@38787.4]
  input        io_sEn_5, // @[:@38787.4]
  input        io_sEn_6, // @[:@38787.4]
  input        io_sDone_0, // @[:@38787.4]
  input        io_sDone_1, // @[:@38787.4]
  input        io_sDone_2, // @[:@38787.4]
  input        io_sDone_3, // @[:@38787.4]
  input        io_sDone_4, // @[:@38787.4]
  input        io_sDone_5, // @[:@38787.4]
  input        io_sDone_6, // @[:@38787.4]
  output [3:0] io_statesInW_0, // @[:@38787.4]
  output [3:0] io_statesInW_1, // @[:@38787.4]
  output [3:0] io_statesInR_6 // @[:@38787.4]
);
  wire  sEn_latch_0_clock; // @[NBuffers.scala 21:52:@38789.4]
  wire  sEn_latch_0_reset; // @[NBuffers.scala 21:52:@38789.4]
  wire  sEn_latch_0_io_input_set; // @[NBuffers.scala 21:52:@38789.4]
  wire  sEn_latch_0_io_input_reset; // @[NBuffers.scala 21:52:@38789.4]
  wire  sEn_latch_0_io_input_asyn_reset; // @[NBuffers.scala 21:52:@38789.4]
  wire  sEn_latch_0_io_output; // @[NBuffers.scala 21:52:@38789.4]
  wire  sEn_latch_1_clock; // @[NBuffers.scala 21:52:@38792.4]
  wire  sEn_latch_1_reset; // @[NBuffers.scala 21:52:@38792.4]
  wire  sEn_latch_1_io_input_set; // @[NBuffers.scala 21:52:@38792.4]
  wire  sEn_latch_1_io_input_reset; // @[NBuffers.scala 21:52:@38792.4]
  wire  sEn_latch_1_io_input_asyn_reset; // @[NBuffers.scala 21:52:@38792.4]
  wire  sEn_latch_1_io_output; // @[NBuffers.scala 21:52:@38792.4]
  wire  sEn_latch_2_clock; // @[NBuffers.scala 21:52:@38795.4]
  wire  sEn_latch_2_reset; // @[NBuffers.scala 21:52:@38795.4]
  wire  sEn_latch_2_io_input_set; // @[NBuffers.scala 21:52:@38795.4]
  wire  sEn_latch_2_io_input_reset; // @[NBuffers.scala 21:52:@38795.4]
  wire  sEn_latch_2_io_input_asyn_reset; // @[NBuffers.scala 21:52:@38795.4]
  wire  sEn_latch_2_io_output; // @[NBuffers.scala 21:52:@38795.4]
  wire  sEn_latch_3_clock; // @[NBuffers.scala 21:52:@38798.4]
  wire  sEn_latch_3_reset; // @[NBuffers.scala 21:52:@38798.4]
  wire  sEn_latch_3_io_input_set; // @[NBuffers.scala 21:52:@38798.4]
  wire  sEn_latch_3_io_input_reset; // @[NBuffers.scala 21:52:@38798.4]
  wire  sEn_latch_3_io_input_asyn_reset; // @[NBuffers.scala 21:52:@38798.4]
  wire  sEn_latch_3_io_output; // @[NBuffers.scala 21:52:@38798.4]
  wire  sEn_latch_4_clock; // @[NBuffers.scala 21:52:@38801.4]
  wire  sEn_latch_4_reset; // @[NBuffers.scala 21:52:@38801.4]
  wire  sEn_latch_4_io_input_set; // @[NBuffers.scala 21:52:@38801.4]
  wire  sEn_latch_4_io_input_reset; // @[NBuffers.scala 21:52:@38801.4]
  wire  sEn_latch_4_io_input_asyn_reset; // @[NBuffers.scala 21:52:@38801.4]
  wire  sEn_latch_4_io_output; // @[NBuffers.scala 21:52:@38801.4]
  wire  sEn_latch_5_clock; // @[NBuffers.scala 21:52:@38804.4]
  wire  sEn_latch_5_reset; // @[NBuffers.scala 21:52:@38804.4]
  wire  sEn_latch_5_io_input_set; // @[NBuffers.scala 21:52:@38804.4]
  wire  sEn_latch_5_io_input_reset; // @[NBuffers.scala 21:52:@38804.4]
  wire  sEn_latch_5_io_input_asyn_reset; // @[NBuffers.scala 21:52:@38804.4]
  wire  sEn_latch_5_io_output; // @[NBuffers.scala 21:52:@38804.4]
  wire  sEn_latch_6_clock; // @[NBuffers.scala 21:52:@38807.4]
  wire  sEn_latch_6_reset; // @[NBuffers.scala 21:52:@38807.4]
  wire  sEn_latch_6_io_input_set; // @[NBuffers.scala 21:52:@38807.4]
  wire  sEn_latch_6_io_input_reset; // @[NBuffers.scala 21:52:@38807.4]
  wire  sEn_latch_6_io_input_asyn_reset; // @[NBuffers.scala 21:52:@38807.4]
  wire  sEn_latch_6_io_output; // @[NBuffers.scala 21:52:@38807.4]
  wire  sDone_latch_0_clock; // @[NBuffers.scala 22:54:@38810.4]
  wire  sDone_latch_0_reset; // @[NBuffers.scala 22:54:@38810.4]
  wire  sDone_latch_0_io_input_set; // @[NBuffers.scala 22:54:@38810.4]
  wire  sDone_latch_0_io_input_reset; // @[NBuffers.scala 22:54:@38810.4]
  wire  sDone_latch_0_io_input_asyn_reset; // @[NBuffers.scala 22:54:@38810.4]
  wire  sDone_latch_0_io_output; // @[NBuffers.scala 22:54:@38810.4]
  wire  sDone_latch_1_clock; // @[NBuffers.scala 22:54:@38813.4]
  wire  sDone_latch_1_reset; // @[NBuffers.scala 22:54:@38813.4]
  wire  sDone_latch_1_io_input_set; // @[NBuffers.scala 22:54:@38813.4]
  wire  sDone_latch_1_io_input_reset; // @[NBuffers.scala 22:54:@38813.4]
  wire  sDone_latch_1_io_input_asyn_reset; // @[NBuffers.scala 22:54:@38813.4]
  wire  sDone_latch_1_io_output; // @[NBuffers.scala 22:54:@38813.4]
  wire  sDone_latch_2_clock; // @[NBuffers.scala 22:54:@38816.4]
  wire  sDone_latch_2_reset; // @[NBuffers.scala 22:54:@38816.4]
  wire  sDone_latch_2_io_input_set; // @[NBuffers.scala 22:54:@38816.4]
  wire  sDone_latch_2_io_input_reset; // @[NBuffers.scala 22:54:@38816.4]
  wire  sDone_latch_2_io_input_asyn_reset; // @[NBuffers.scala 22:54:@38816.4]
  wire  sDone_latch_2_io_output; // @[NBuffers.scala 22:54:@38816.4]
  wire  sDone_latch_3_clock; // @[NBuffers.scala 22:54:@38819.4]
  wire  sDone_latch_3_reset; // @[NBuffers.scala 22:54:@38819.4]
  wire  sDone_latch_3_io_input_set; // @[NBuffers.scala 22:54:@38819.4]
  wire  sDone_latch_3_io_input_reset; // @[NBuffers.scala 22:54:@38819.4]
  wire  sDone_latch_3_io_input_asyn_reset; // @[NBuffers.scala 22:54:@38819.4]
  wire  sDone_latch_3_io_output; // @[NBuffers.scala 22:54:@38819.4]
  wire  sDone_latch_4_clock; // @[NBuffers.scala 22:54:@38822.4]
  wire  sDone_latch_4_reset; // @[NBuffers.scala 22:54:@38822.4]
  wire  sDone_latch_4_io_input_set; // @[NBuffers.scala 22:54:@38822.4]
  wire  sDone_latch_4_io_input_reset; // @[NBuffers.scala 22:54:@38822.4]
  wire  sDone_latch_4_io_input_asyn_reset; // @[NBuffers.scala 22:54:@38822.4]
  wire  sDone_latch_4_io_output; // @[NBuffers.scala 22:54:@38822.4]
  wire  sDone_latch_5_clock; // @[NBuffers.scala 22:54:@38825.4]
  wire  sDone_latch_5_reset; // @[NBuffers.scala 22:54:@38825.4]
  wire  sDone_latch_5_io_input_set; // @[NBuffers.scala 22:54:@38825.4]
  wire  sDone_latch_5_io_input_reset; // @[NBuffers.scala 22:54:@38825.4]
  wire  sDone_latch_5_io_input_asyn_reset; // @[NBuffers.scala 22:54:@38825.4]
  wire  sDone_latch_5_io_output; // @[NBuffers.scala 22:54:@38825.4]
  wire  sDone_latch_6_clock; // @[NBuffers.scala 22:54:@38828.4]
  wire  sDone_latch_6_reset; // @[NBuffers.scala 22:54:@38828.4]
  wire  sDone_latch_6_io_input_set; // @[NBuffers.scala 22:54:@38828.4]
  wire  sDone_latch_6_io_input_reset; // @[NBuffers.scala 22:54:@38828.4]
  wire  sDone_latch_6_io_input_asyn_reset; // @[NBuffers.scala 22:54:@38828.4]
  wire  sDone_latch_6_io_output; // @[NBuffers.scala 22:54:@38828.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@38835.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@38835.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@38835.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@38835.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@38835.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@38843.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@38843.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@38843.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@38843.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@38843.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@38852.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@38852.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@38852.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@38852.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@38852.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@38860.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@38860.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@38860.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@38860.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@38860.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@38871.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@38871.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@38871.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@38871.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@38871.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@38879.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@38879.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@38879.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@38879.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@38879.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@38888.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@38888.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@38888.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@38888.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@38888.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@38896.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@38896.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@38896.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@38896.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@38896.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@38907.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@38907.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@38907.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@38907.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@38907.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@38915.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@38915.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@38915.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@38915.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@38915.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@38924.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@38924.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@38924.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@38924.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@38924.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@38932.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@38932.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@38932.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@38932.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@38932.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@38943.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@38943.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@38943.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@38943.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@38943.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@38951.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@38951.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@38951.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@38951.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@38951.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@38960.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@38960.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@38960.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@38960.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@38960.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@38968.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@38968.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@38968.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@38968.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@38968.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@38979.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@38979.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@38979.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@38979.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@38979.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@38987.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@38987.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@38987.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@38987.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@38987.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@38996.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@38996.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@38996.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@38996.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@38996.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@39004.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@39004.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@39004.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@39004.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@39004.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@39015.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@39015.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@39015.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@39015.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@39015.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@39023.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@39023.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@39023.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@39023.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@39023.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@39032.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@39032.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@39032.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@39032.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@39032.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@39040.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@39040.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@39040.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@39040.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@39040.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@39051.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@39051.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@39051.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@39051.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@39051.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@39059.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@39059.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@39059.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@39059.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@39059.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@39068.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@39068.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@39068.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@39068.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@39068.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@39076.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@39076.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@39076.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@39076.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@39076.4]
  wire  NBufCtr_clock; // @[NBuffers.scala 40:19:@39117.4]
  wire  NBufCtr_reset; // @[NBuffers.scala 40:19:@39117.4]
  wire  NBufCtr_io_input_countUp; // @[NBuffers.scala 40:19:@39117.4]
  wire  NBufCtr_io_input_enable; // @[NBuffers.scala 40:19:@39117.4]
  wire [31:0] NBufCtr_io_output_count; // @[NBuffers.scala 40:19:@39117.4]
  wire  NBufCtr_1_clock; // @[NBuffers.scala 40:19:@39128.4]
  wire  NBufCtr_1_reset; // @[NBuffers.scala 40:19:@39128.4]
  wire  NBufCtr_1_io_input_countUp; // @[NBuffers.scala 40:19:@39128.4]
  wire  NBufCtr_1_io_input_enable; // @[NBuffers.scala 40:19:@39128.4]
  wire [31:0] NBufCtr_1_io_output_count; // @[NBuffers.scala 40:19:@39128.4]
  wire  statesInR_0_clock; // @[NBuffers.scala 50:19:@39139.4]
  wire  statesInR_0_reset; // @[NBuffers.scala 50:19:@39139.4]
  wire  statesInR_0_io_input_countUp; // @[NBuffers.scala 50:19:@39139.4]
  wire  statesInR_0_io_input_enable; // @[NBuffers.scala 50:19:@39139.4]
  wire [31:0] statesInR_0_io_output_count; // @[NBuffers.scala 50:19:@39139.4]
  wire  statesInR_1_clock; // @[NBuffers.scala 50:19:@39150.4]
  wire  statesInR_1_reset; // @[NBuffers.scala 50:19:@39150.4]
  wire  statesInR_1_io_input_countUp; // @[NBuffers.scala 50:19:@39150.4]
  wire  statesInR_1_io_input_enable; // @[NBuffers.scala 50:19:@39150.4]
  wire [31:0] statesInR_1_io_output_count; // @[NBuffers.scala 50:19:@39150.4]
  wire  statesInR_2_clock; // @[NBuffers.scala 50:19:@39161.4]
  wire  statesInR_2_reset; // @[NBuffers.scala 50:19:@39161.4]
  wire  statesInR_2_io_input_countUp; // @[NBuffers.scala 50:19:@39161.4]
  wire  statesInR_2_io_input_enable; // @[NBuffers.scala 50:19:@39161.4]
  wire [31:0] statesInR_2_io_output_count; // @[NBuffers.scala 50:19:@39161.4]
  wire  statesInR_3_clock; // @[NBuffers.scala 50:19:@39172.4]
  wire  statesInR_3_reset; // @[NBuffers.scala 50:19:@39172.4]
  wire  statesInR_3_io_input_countUp; // @[NBuffers.scala 50:19:@39172.4]
  wire  statesInR_3_io_input_enable; // @[NBuffers.scala 50:19:@39172.4]
  wire [31:0] statesInR_3_io_output_count; // @[NBuffers.scala 50:19:@39172.4]
  wire  statesInR_4_clock; // @[NBuffers.scala 50:19:@39183.4]
  wire  statesInR_4_reset; // @[NBuffers.scala 50:19:@39183.4]
  wire  statesInR_4_io_input_countUp; // @[NBuffers.scala 50:19:@39183.4]
  wire  statesInR_4_io_input_enable; // @[NBuffers.scala 50:19:@39183.4]
  wire [31:0] statesInR_4_io_output_count; // @[NBuffers.scala 50:19:@39183.4]
  wire  statesInR_5_clock; // @[NBuffers.scala 50:19:@39194.4]
  wire  statesInR_5_reset; // @[NBuffers.scala 50:19:@39194.4]
  wire  statesInR_5_io_input_countUp; // @[NBuffers.scala 50:19:@39194.4]
  wire  statesInR_5_io_input_enable; // @[NBuffers.scala 50:19:@39194.4]
  wire [31:0] statesInR_5_io_output_count; // @[NBuffers.scala 50:19:@39194.4]
  wire  statesInR_6_clock; // @[NBuffers.scala 50:19:@39205.4]
  wire  statesInR_6_reset; // @[NBuffers.scala 50:19:@39205.4]
  wire  statesInR_6_io_input_countUp; // @[NBuffers.scala 50:19:@39205.4]
  wire  statesInR_6_io_input_enable; // @[NBuffers.scala 50:19:@39205.4]
  wire [31:0] statesInR_6_io_output_count; // @[NBuffers.scala 50:19:@39205.4]
  wire  _T_33; // @[NBuffers.scala 26:46:@38832.4]
  wire  _T_48; // @[NBuffers.scala 26:46:@38868.4]
  wire  _T_63; // @[NBuffers.scala 26:46:@38904.4]
  wire  _T_78; // @[NBuffers.scala 26:46:@38940.4]
  wire  _T_93; // @[NBuffers.scala 26:46:@38976.4]
  wire  _T_108; // @[NBuffers.scala 26:46:@39012.4]
  wire  _T_123; // @[NBuffers.scala 26:46:@39048.4]
  wire  _T_137; // @[NBuffers.scala 33:64:@39084.4]
  wire  _T_138; // @[NBuffers.scala 33:64:@39085.4]
  wire  _T_139; // @[NBuffers.scala 33:64:@39086.4]
  wire  _T_140; // @[NBuffers.scala 33:64:@39087.4]
  wire  _T_141; // @[NBuffers.scala 33:64:@39088.4]
  wire  anyEnabled; // @[NBuffers.scala 33:64:@39089.4]
  wire  _T_142; // @[NBuffers.scala 34:124:@39090.4]
  wire  _T_143; // @[NBuffers.scala 34:104:@39091.4]
  wire  _T_144; // @[NBuffers.scala 34:124:@39092.4]
  wire  _T_145; // @[NBuffers.scala 34:104:@39093.4]
  wire  _T_146; // @[NBuffers.scala 34:124:@39094.4]
  wire  _T_147; // @[NBuffers.scala 34:104:@39095.4]
  wire  _T_148; // @[NBuffers.scala 34:124:@39096.4]
  wire  _T_149; // @[NBuffers.scala 34:104:@39097.4]
  wire  _T_150; // @[NBuffers.scala 34:124:@39098.4]
  wire  _T_151; // @[NBuffers.scala 34:104:@39099.4]
  wire  _T_152; // @[NBuffers.scala 34:124:@39100.4]
  wire  _T_153; // @[NBuffers.scala 34:104:@39101.4]
  wire  _T_154; // @[NBuffers.scala 34:124:@39102.4]
  wire  _T_155; // @[NBuffers.scala 34:104:@39103.4]
  wire  _T_156; // @[NBuffers.scala 34:150:@39104.4]
  wire  _T_157; // @[NBuffers.scala 34:150:@39105.4]
  wire  _T_158; // @[NBuffers.scala 34:150:@39106.4]
  wire  _T_159; // @[NBuffers.scala 34:150:@39107.4]
  wire  _T_160; // @[NBuffers.scala 34:150:@39108.4]
  wire  _T_161; // @[NBuffers.scala 34:150:@39109.4]
  wire  _T_162; // @[NBuffers.scala 34:154:@39110.4]
  wire  _T_164; // @[package.scala 100:49:@39111.4]
  reg  _T_167; // @[package.scala 48:56:@39112.4]
  reg [31:0] _RAND_0;
  SRFF sEn_latch_0 ( // @[NBuffers.scala 21:52:@38789.4]
    .clock(sEn_latch_0_clock),
    .reset(sEn_latch_0_reset),
    .io_input_set(sEn_latch_0_io_input_set),
    .io_input_reset(sEn_latch_0_io_input_reset),
    .io_input_asyn_reset(sEn_latch_0_io_input_asyn_reset),
    .io_output(sEn_latch_0_io_output)
  );
  SRFF sEn_latch_1 ( // @[NBuffers.scala 21:52:@38792.4]
    .clock(sEn_latch_1_clock),
    .reset(sEn_latch_1_reset),
    .io_input_set(sEn_latch_1_io_input_set),
    .io_input_reset(sEn_latch_1_io_input_reset),
    .io_input_asyn_reset(sEn_latch_1_io_input_asyn_reset),
    .io_output(sEn_latch_1_io_output)
  );
  SRFF sEn_latch_2 ( // @[NBuffers.scala 21:52:@38795.4]
    .clock(sEn_latch_2_clock),
    .reset(sEn_latch_2_reset),
    .io_input_set(sEn_latch_2_io_input_set),
    .io_input_reset(sEn_latch_2_io_input_reset),
    .io_input_asyn_reset(sEn_latch_2_io_input_asyn_reset),
    .io_output(sEn_latch_2_io_output)
  );
  SRFF sEn_latch_3 ( // @[NBuffers.scala 21:52:@38798.4]
    .clock(sEn_latch_3_clock),
    .reset(sEn_latch_3_reset),
    .io_input_set(sEn_latch_3_io_input_set),
    .io_input_reset(sEn_latch_3_io_input_reset),
    .io_input_asyn_reset(sEn_latch_3_io_input_asyn_reset),
    .io_output(sEn_latch_3_io_output)
  );
  SRFF sEn_latch_4 ( // @[NBuffers.scala 21:52:@38801.4]
    .clock(sEn_latch_4_clock),
    .reset(sEn_latch_4_reset),
    .io_input_set(sEn_latch_4_io_input_set),
    .io_input_reset(sEn_latch_4_io_input_reset),
    .io_input_asyn_reset(sEn_latch_4_io_input_asyn_reset),
    .io_output(sEn_latch_4_io_output)
  );
  SRFF sEn_latch_5 ( // @[NBuffers.scala 21:52:@38804.4]
    .clock(sEn_latch_5_clock),
    .reset(sEn_latch_5_reset),
    .io_input_set(sEn_latch_5_io_input_set),
    .io_input_reset(sEn_latch_5_io_input_reset),
    .io_input_asyn_reset(sEn_latch_5_io_input_asyn_reset),
    .io_output(sEn_latch_5_io_output)
  );
  SRFF sEn_latch_6 ( // @[NBuffers.scala 21:52:@38807.4]
    .clock(sEn_latch_6_clock),
    .reset(sEn_latch_6_reset),
    .io_input_set(sEn_latch_6_io_input_set),
    .io_input_reset(sEn_latch_6_io_input_reset),
    .io_input_asyn_reset(sEn_latch_6_io_input_asyn_reset),
    .io_output(sEn_latch_6_io_output)
  );
  SRFF sDone_latch_0 ( // @[NBuffers.scala 22:54:@38810.4]
    .clock(sDone_latch_0_clock),
    .reset(sDone_latch_0_reset),
    .io_input_set(sDone_latch_0_io_input_set),
    .io_input_reset(sDone_latch_0_io_input_reset),
    .io_input_asyn_reset(sDone_latch_0_io_input_asyn_reset),
    .io_output(sDone_latch_0_io_output)
  );
  SRFF sDone_latch_1 ( // @[NBuffers.scala 22:54:@38813.4]
    .clock(sDone_latch_1_clock),
    .reset(sDone_latch_1_reset),
    .io_input_set(sDone_latch_1_io_input_set),
    .io_input_reset(sDone_latch_1_io_input_reset),
    .io_input_asyn_reset(sDone_latch_1_io_input_asyn_reset),
    .io_output(sDone_latch_1_io_output)
  );
  SRFF sDone_latch_2 ( // @[NBuffers.scala 22:54:@38816.4]
    .clock(sDone_latch_2_clock),
    .reset(sDone_latch_2_reset),
    .io_input_set(sDone_latch_2_io_input_set),
    .io_input_reset(sDone_latch_2_io_input_reset),
    .io_input_asyn_reset(sDone_latch_2_io_input_asyn_reset),
    .io_output(sDone_latch_2_io_output)
  );
  SRFF sDone_latch_3 ( // @[NBuffers.scala 22:54:@38819.4]
    .clock(sDone_latch_3_clock),
    .reset(sDone_latch_3_reset),
    .io_input_set(sDone_latch_3_io_input_set),
    .io_input_reset(sDone_latch_3_io_input_reset),
    .io_input_asyn_reset(sDone_latch_3_io_input_asyn_reset),
    .io_output(sDone_latch_3_io_output)
  );
  SRFF sDone_latch_4 ( // @[NBuffers.scala 22:54:@38822.4]
    .clock(sDone_latch_4_clock),
    .reset(sDone_latch_4_reset),
    .io_input_set(sDone_latch_4_io_input_set),
    .io_input_reset(sDone_latch_4_io_input_reset),
    .io_input_asyn_reset(sDone_latch_4_io_input_asyn_reset),
    .io_output(sDone_latch_4_io_output)
  );
  SRFF sDone_latch_5 ( // @[NBuffers.scala 22:54:@38825.4]
    .clock(sDone_latch_5_clock),
    .reset(sDone_latch_5_reset),
    .io_input_set(sDone_latch_5_io_input_set),
    .io_input_reset(sDone_latch_5_io_input_reset),
    .io_input_asyn_reset(sDone_latch_5_io_input_asyn_reset),
    .io_output(sDone_latch_5_io_output)
  );
  SRFF sDone_latch_6 ( // @[NBuffers.scala 22:54:@38828.4]
    .clock(sDone_latch_6_clock),
    .reset(sDone_latch_6_reset),
    .io_input_set(sDone_latch_6_io_input_set),
    .io_input_reset(sDone_latch_6_io_input_reset),
    .io_input_asyn_reset(sDone_latch_6_io_input_asyn_reset),
    .io_output(sDone_latch_6_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@38835.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@38843.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@38852.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@38860.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@38871.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@38879.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@38888.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@38896.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@38907.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@38915.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@38924.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 ( // @[package.scala 93:22:@38932.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper RetimeWrapper_12 ( // @[package.scala 93:22:@38943.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 ( // @[package.scala 93:22:@38951.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@38960.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@38968.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 ( // @[package.scala 93:22:@38979.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper RetimeWrapper_17 ( // @[package.scala 93:22:@38987.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 ( // @[package.scala 93:22:@38996.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper RetimeWrapper_19 ( // @[package.scala 93:22:@39004.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper RetimeWrapper_20 ( // @[package.scala 93:22:@39015.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper RetimeWrapper_21 ( // @[package.scala 93:22:@39023.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper RetimeWrapper_22 ( // @[package.scala 93:22:@39032.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper RetimeWrapper_23 ( // @[package.scala 93:22:@39040.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper RetimeWrapper_24 ( // @[package.scala 93:22:@39051.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@39059.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper RetimeWrapper_26 ( // @[package.scala 93:22:@39068.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper RetimeWrapper_27 ( // @[package.scala 93:22:@39076.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  NBufCtr_9 NBufCtr ( // @[NBuffers.scala 40:19:@39117.4]
    .clock(NBufCtr_clock),
    .reset(NBufCtr_reset),
    .io_input_countUp(NBufCtr_io_input_countUp),
    .io_input_enable(NBufCtr_io_input_enable),
    .io_output_count(NBufCtr_io_output_count)
  );
  NBufCtr_15 NBufCtr_1 ( // @[NBuffers.scala 40:19:@39128.4]
    .clock(NBufCtr_1_clock),
    .reset(NBufCtr_1_reset),
    .io_input_countUp(NBufCtr_1_io_input_countUp),
    .io_input_enable(NBufCtr_1_io_input_enable),
    .io_output_count(NBufCtr_1_io_output_count)
  );
  NBufCtr_9 statesInR_0 ( // @[NBuffers.scala 50:19:@39139.4]
    .clock(statesInR_0_clock),
    .reset(statesInR_0_reset),
    .io_input_countUp(statesInR_0_io_input_countUp),
    .io_input_enable(statesInR_0_io_input_enable),
    .io_output_count(statesInR_0_io_output_count)
  );
  NBufCtr_11 statesInR_1 ( // @[NBuffers.scala 50:19:@39150.4]
    .clock(statesInR_1_clock),
    .reset(statesInR_1_reset),
    .io_input_countUp(statesInR_1_io_input_countUp),
    .io_input_enable(statesInR_1_io_input_enable),
    .io_output_count(statesInR_1_io_output_count)
  );
  NBufCtr_12 statesInR_2 ( // @[NBuffers.scala 50:19:@39161.4]
    .clock(statesInR_2_clock),
    .reset(statesInR_2_reset),
    .io_input_countUp(statesInR_2_io_input_countUp),
    .io_input_enable(statesInR_2_io_input_enable),
    .io_output_count(statesInR_2_io_output_count)
  );
  NBufCtr_13 statesInR_3 ( // @[NBuffers.scala 50:19:@39172.4]
    .clock(statesInR_3_clock),
    .reset(statesInR_3_reset),
    .io_input_countUp(statesInR_3_io_input_countUp),
    .io_input_enable(statesInR_3_io_input_enable),
    .io_output_count(statesInR_3_io_output_count)
  );
  NBufCtr_14 statesInR_4 ( // @[NBuffers.scala 50:19:@39183.4]
    .clock(statesInR_4_clock),
    .reset(statesInR_4_reset),
    .io_input_countUp(statesInR_4_io_input_countUp),
    .io_input_enable(statesInR_4_io_input_enable),
    .io_output_count(statesInR_4_io_output_count)
  );
  NBufCtr_15 statesInR_5 ( // @[NBuffers.scala 50:19:@39194.4]
    .clock(statesInR_5_clock),
    .reset(statesInR_5_reset),
    .io_input_countUp(statesInR_5_io_input_countUp),
    .io_input_enable(statesInR_5_io_input_enable),
    .io_output_count(statesInR_5_io_output_count)
  );
  NBufCtr_16 statesInR_6 ( // @[NBuffers.scala 50:19:@39205.4]
    .clock(statesInR_6_clock),
    .reset(statesInR_6_reset),
    .io_input_countUp(statesInR_6_io_input_countUp),
    .io_input_enable(statesInR_6_io_input_enable),
    .io_output_count(statesInR_6_io_output_count)
  );
  assign _T_33 = io_sDone_0 == 1'h0; // @[NBuffers.scala 26:46:@38832.4]
  assign _T_48 = io_sDone_1 == 1'h0; // @[NBuffers.scala 26:46:@38868.4]
  assign _T_63 = io_sDone_2 == 1'h0; // @[NBuffers.scala 26:46:@38904.4]
  assign _T_78 = io_sDone_3 == 1'h0; // @[NBuffers.scala 26:46:@38940.4]
  assign _T_93 = io_sDone_4 == 1'h0; // @[NBuffers.scala 26:46:@38976.4]
  assign _T_108 = io_sDone_5 == 1'h0; // @[NBuffers.scala 26:46:@39012.4]
  assign _T_123 = io_sDone_6 == 1'h0; // @[NBuffers.scala 26:46:@39048.4]
  assign _T_137 = sEn_latch_0_io_output | sEn_latch_1_io_output; // @[NBuffers.scala 33:64:@39084.4]
  assign _T_138 = _T_137 | sEn_latch_2_io_output; // @[NBuffers.scala 33:64:@39085.4]
  assign _T_139 = _T_138 | sEn_latch_3_io_output; // @[NBuffers.scala 33:64:@39086.4]
  assign _T_140 = _T_139 | sEn_latch_4_io_output; // @[NBuffers.scala 33:64:@39087.4]
  assign _T_141 = _T_140 | sEn_latch_5_io_output; // @[NBuffers.scala 33:64:@39088.4]
  assign anyEnabled = _T_141 | sEn_latch_6_io_output; // @[NBuffers.scala 33:64:@39089.4]
  assign _T_142 = sDone_latch_0_io_output | io_sDone_0; // @[NBuffers.scala 34:124:@39090.4]
  assign _T_143 = sEn_latch_0_io_output == _T_142; // @[NBuffers.scala 34:104:@39091.4]
  assign _T_144 = sDone_latch_1_io_output | io_sDone_1; // @[NBuffers.scala 34:124:@39092.4]
  assign _T_145 = sEn_latch_1_io_output == _T_144; // @[NBuffers.scala 34:104:@39093.4]
  assign _T_146 = sDone_latch_2_io_output | io_sDone_2; // @[NBuffers.scala 34:124:@39094.4]
  assign _T_147 = sEn_latch_2_io_output == _T_146; // @[NBuffers.scala 34:104:@39095.4]
  assign _T_148 = sDone_latch_3_io_output | io_sDone_3; // @[NBuffers.scala 34:124:@39096.4]
  assign _T_149 = sEn_latch_3_io_output == _T_148; // @[NBuffers.scala 34:104:@39097.4]
  assign _T_150 = sDone_latch_4_io_output | io_sDone_4; // @[NBuffers.scala 34:124:@39098.4]
  assign _T_151 = sEn_latch_4_io_output == _T_150; // @[NBuffers.scala 34:104:@39099.4]
  assign _T_152 = sDone_latch_5_io_output | io_sDone_5; // @[NBuffers.scala 34:124:@39100.4]
  assign _T_153 = sEn_latch_5_io_output == _T_152; // @[NBuffers.scala 34:104:@39101.4]
  assign _T_154 = sDone_latch_6_io_output | io_sDone_6; // @[NBuffers.scala 34:124:@39102.4]
  assign _T_155 = sEn_latch_6_io_output == _T_154; // @[NBuffers.scala 34:104:@39103.4]
  assign _T_156 = _T_143 & _T_145; // @[NBuffers.scala 34:150:@39104.4]
  assign _T_157 = _T_156 & _T_147; // @[NBuffers.scala 34:150:@39105.4]
  assign _T_158 = _T_157 & _T_149; // @[NBuffers.scala 34:150:@39106.4]
  assign _T_159 = _T_158 & _T_151; // @[NBuffers.scala 34:150:@39107.4]
  assign _T_160 = _T_159 & _T_153; // @[NBuffers.scala 34:150:@39108.4]
  assign _T_161 = _T_160 & _T_155; // @[NBuffers.scala 34:150:@39109.4]
  assign _T_162 = _T_161 & anyEnabled; // @[NBuffers.scala 34:154:@39110.4]
  assign _T_164 = _T_162 == 1'h0; // @[package.scala 100:49:@39111.4]
  assign io_statesInW_0 = NBufCtr_io_output_count[3:0]; // @[NBuffers.scala 44:21:@39127.4]
  assign io_statesInW_1 = NBufCtr_1_io_output_count[3:0]; // @[NBuffers.scala 44:21:@39138.4]
  assign io_statesInR_6 = statesInR_6_io_output_count[3:0]; // @[NBuffers.scala 54:21:@39215.4]
  assign sEn_latch_0_clock = clock; // @[:@38790.4]
  assign sEn_latch_0_reset = reset; // @[:@38791.4]
  assign sEn_latch_0_io_input_set = io_sEn_0 & _T_33; // @[NBuffers.scala 26:31:@38834.4]
  assign sEn_latch_0_io_input_reset = RetimeWrapper_io_out; // @[NBuffers.scala 27:33:@38842.4]
  assign sEn_latch_0_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[NBuffers.scala 28:38:@38850.4]
  assign sEn_latch_1_clock = clock; // @[:@38793.4]
  assign sEn_latch_1_reset = reset; // @[:@38794.4]
  assign sEn_latch_1_io_input_set = io_sEn_1 & _T_48; // @[NBuffers.scala 26:31:@38870.4]
  assign sEn_latch_1_io_input_reset = RetimeWrapper_4_io_out; // @[NBuffers.scala 27:33:@38878.4]
  assign sEn_latch_1_io_input_asyn_reset = RetimeWrapper_5_io_out; // @[NBuffers.scala 28:38:@38886.4]
  assign sEn_latch_2_clock = clock; // @[:@38796.4]
  assign sEn_latch_2_reset = reset; // @[:@38797.4]
  assign sEn_latch_2_io_input_set = io_sEn_2 & _T_63; // @[NBuffers.scala 26:31:@38906.4]
  assign sEn_latch_2_io_input_reset = RetimeWrapper_8_io_out; // @[NBuffers.scala 27:33:@38914.4]
  assign sEn_latch_2_io_input_asyn_reset = RetimeWrapper_9_io_out; // @[NBuffers.scala 28:38:@38922.4]
  assign sEn_latch_3_clock = clock; // @[:@38799.4]
  assign sEn_latch_3_reset = reset; // @[:@38800.4]
  assign sEn_latch_3_io_input_set = io_sEn_3 & _T_78; // @[NBuffers.scala 26:31:@38942.4]
  assign sEn_latch_3_io_input_reset = RetimeWrapper_12_io_out; // @[NBuffers.scala 27:33:@38950.4]
  assign sEn_latch_3_io_input_asyn_reset = RetimeWrapper_13_io_out; // @[NBuffers.scala 28:38:@38958.4]
  assign sEn_latch_4_clock = clock; // @[:@38802.4]
  assign sEn_latch_4_reset = reset; // @[:@38803.4]
  assign sEn_latch_4_io_input_set = io_sEn_4 & _T_93; // @[NBuffers.scala 26:31:@38978.4]
  assign sEn_latch_4_io_input_reset = RetimeWrapper_16_io_out; // @[NBuffers.scala 27:33:@38986.4]
  assign sEn_latch_4_io_input_asyn_reset = RetimeWrapper_17_io_out; // @[NBuffers.scala 28:38:@38994.4]
  assign sEn_latch_5_clock = clock; // @[:@38805.4]
  assign sEn_latch_5_reset = reset; // @[:@38806.4]
  assign sEn_latch_5_io_input_set = io_sEn_5 & _T_108; // @[NBuffers.scala 26:31:@39014.4]
  assign sEn_latch_5_io_input_reset = RetimeWrapper_20_io_out; // @[NBuffers.scala 27:33:@39022.4]
  assign sEn_latch_5_io_input_asyn_reset = RetimeWrapper_21_io_out; // @[NBuffers.scala 28:38:@39030.4]
  assign sEn_latch_6_clock = clock; // @[:@38808.4]
  assign sEn_latch_6_reset = reset; // @[:@38809.4]
  assign sEn_latch_6_io_input_set = io_sEn_6 & _T_123; // @[NBuffers.scala 26:31:@39050.4]
  assign sEn_latch_6_io_input_reset = RetimeWrapper_24_io_out; // @[NBuffers.scala 27:33:@39058.4]
  assign sEn_latch_6_io_input_asyn_reset = RetimeWrapper_25_io_out; // @[NBuffers.scala 28:38:@39066.4]
  assign sDone_latch_0_clock = clock; // @[:@38811.4]
  assign sDone_latch_0_reset = reset; // @[:@38812.4]
  assign sDone_latch_0_io_input_set = io_sDone_0; // @[NBuffers.scala 29:33:@38851.4]
  assign sDone_latch_0_io_input_reset = RetimeWrapper_2_io_out; // @[NBuffers.scala 30:35:@38859.4]
  assign sDone_latch_0_io_input_asyn_reset = RetimeWrapper_3_io_out; // @[NBuffers.scala 31:40:@38867.4]
  assign sDone_latch_1_clock = clock; // @[:@38814.4]
  assign sDone_latch_1_reset = reset; // @[:@38815.4]
  assign sDone_latch_1_io_input_set = io_sDone_1; // @[NBuffers.scala 29:33:@38887.4]
  assign sDone_latch_1_io_input_reset = RetimeWrapper_6_io_out; // @[NBuffers.scala 30:35:@38895.4]
  assign sDone_latch_1_io_input_asyn_reset = RetimeWrapper_7_io_out; // @[NBuffers.scala 31:40:@38903.4]
  assign sDone_latch_2_clock = clock; // @[:@38817.4]
  assign sDone_latch_2_reset = reset; // @[:@38818.4]
  assign sDone_latch_2_io_input_set = io_sDone_2; // @[NBuffers.scala 29:33:@38923.4]
  assign sDone_latch_2_io_input_reset = RetimeWrapper_10_io_out; // @[NBuffers.scala 30:35:@38931.4]
  assign sDone_latch_2_io_input_asyn_reset = RetimeWrapper_11_io_out; // @[NBuffers.scala 31:40:@38939.4]
  assign sDone_latch_3_clock = clock; // @[:@38820.4]
  assign sDone_latch_3_reset = reset; // @[:@38821.4]
  assign sDone_latch_3_io_input_set = io_sDone_3; // @[NBuffers.scala 29:33:@38959.4]
  assign sDone_latch_3_io_input_reset = RetimeWrapper_14_io_out; // @[NBuffers.scala 30:35:@38967.4]
  assign sDone_latch_3_io_input_asyn_reset = RetimeWrapper_15_io_out; // @[NBuffers.scala 31:40:@38975.4]
  assign sDone_latch_4_clock = clock; // @[:@38823.4]
  assign sDone_latch_4_reset = reset; // @[:@38824.4]
  assign sDone_latch_4_io_input_set = io_sDone_4; // @[NBuffers.scala 29:33:@38995.4]
  assign sDone_latch_4_io_input_reset = RetimeWrapper_18_io_out; // @[NBuffers.scala 30:35:@39003.4]
  assign sDone_latch_4_io_input_asyn_reset = RetimeWrapper_19_io_out; // @[NBuffers.scala 31:40:@39011.4]
  assign sDone_latch_5_clock = clock; // @[:@38826.4]
  assign sDone_latch_5_reset = reset; // @[:@38827.4]
  assign sDone_latch_5_io_input_set = io_sDone_5; // @[NBuffers.scala 29:33:@39031.4]
  assign sDone_latch_5_io_input_reset = RetimeWrapper_22_io_out; // @[NBuffers.scala 30:35:@39039.4]
  assign sDone_latch_5_io_input_asyn_reset = RetimeWrapper_23_io_out; // @[NBuffers.scala 31:40:@39047.4]
  assign sDone_latch_6_clock = clock; // @[:@38829.4]
  assign sDone_latch_6_reset = reset; // @[:@38830.4]
  assign sDone_latch_6_io_input_set = io_sDone_6; // @[NBuffers.scala 29:33:@39067.4]
  assign sDone_latch_6_io_input_reset = RetimeWrapper_26_io_out; // @[NBuffers.scala 30:35:@39075.4]
  assign sDone_latch_6_io_input_asyn_reset = RetimeWrapper_27_io_out; // @[NBuffers.scala 31:40:@39083.4]
  assign RetimeWrapper_clock = clock; // @[:@38836.4]
  assign RetimeWrapper_reset = reset; // @[:@38837.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@38839.4]
  assign RetimeWrapper_io_in = _T_162 & _T_167; // @[package.scala 94:16:@38838.4]
  assign RetimeWrapper_1_clock = clock; // @[:@38844.4]
  assign RetimeWrapper_1_reset = reset; // @[:@38845.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@38847.4]
  assign RetimeWrapper_1_io_in = reset; // @[package.scala 94:16:@38846.4]
  assign RetimeWrapper_2_clock = clock; // @[:@38853.4]
  assign RetimeWrapper_2_reset = reset; // @[:@38854.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@38856.4]
  assign RetimeWrapper_2_io_in = _T_162 & _T_167; // @[package.scala 94:16:@38855.4]
  assign RetimeWrapper_3_clock = clock; // @[:@38861.4]
  assign RetimeWrapper_3_reset = reset; // @[:@38862.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@38864.4]
  assign RetimeWrapper_3_io_in = reset; // @[package.scala 94:16:@38863.4]
  assign RetimeWrapper_4_clock = clock; // @[:@38872.4]
  assign RetimeWrapper_4_reset = reset; // @[:@38873.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@38875.4]
  assign RetimeWrapper_4_io_in = _T_162 & _T_167; // @[package.scala 94:16:@38874.4]
  assign RetimeWrapper_5_clock = clock; // @[:@38880.4]
  assign RetimeWrapper_5_reset = reset; // @[:@38881.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@38883.4]
  assign RetimeWrapper_5_io_in = reset; // @[package.scala 94:16:@38882.4]
  assign RetimeWrapper_6_clock = clock; // @[:@38889.4]
  assign RetimeWrapper_6_reset = reset; // @[:@38890.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@38892.4]
  assign RetimeWrapper_6_io_in = _T_162 & _T_167; // @[package.scala 94:16:@38891.4]
  assign RetimeWrapper_7_clock = clock; // @[:@38897.4]
  assign RetimeWrapper_7_reset = reset; // @[:@38898.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@38900.4]
  assign RetimeWrapper_7_io_in = reset; // @[package.scala 94:16:@38899.4]
  assign RetimeWrapper_8_clock = clock; // @[:@38908.4]
  assign RetimeWrapper_8_reset = reset; // @[:@38909.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@38911.4]
  assign RetimeWrapper_8_io_in = _T_162 & _T_167; // @[package.scala 94:16:@38910.4]
  assign RetimeWrapper_9_clock = clock; // @[:@38916.4]
  assign RetimeWrapper_9_reset = reset; // @[:@38917.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@38919.4]
  assign RetimeWrapper_9_io_in = reset; // @[package.scala 94:16:@38918.4]
  assign RetimeWrapper_10_clock = clock; // @[:@38925.4]
  assign RetimeWrapper_10_reset = reset; // @[:@38926.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@38928.4]
  assign RetimeWrapper_10_io_in = _T_162 & _T_167; // @[package.scala 94:16:@38927.4]
  assign RetimeWrapper_11_clock = clock; // @[:@38933.4]
  assign RetimeWrapper_11_reset = reset; // @[:@38934.4]
  assign RetimeWrapper_11_io_flow = 1'h1; // @[package.scala 95:18:@38936.4]
  assign RetimeWrapper_11_io_in = reset; // @[package.scala 94:16:@38935.4]
  assign RetimeWrapper_12_clock = clock; // @[:@38944.4]
  assign RetimeWrapper_12_reset = reset; // @[:@38945.4]
  assign RetimeWrapper_12_io_flow = 1'h1; // @[package.scala 95:18:@38947.4]
  assign RetimeWrapper_12_io_in = _T_162 & _T_167; // @[package.scala 94:16:@38946.4]
  assign RetimeWrapper_13_clock = clock; // @[:@38952.4]
  assign RetimeWrapper_13_reset = reset; // @[:@38953.4]
  assign RetimeWrapper_13_io_flow = 1'h1; // @[package.scala 95:18:@38955.4]
  assign RetimeWrapper_13_io_in = reset; // @[package.scala 94:16:@38954.4]
  assign RetimeWrapper_14_clock = clock; // @[:@38961.4]
  assign RetimeWrapper_14_reset = reset; // @[:@38962.4]
  assign RetimeWrapper_14_io_flow = 1'h1; // @[package.scala 95:18:@38964.4]
  assign RetimeWrapper_14_io_in = _T_162 & _T_167; // @[package.scala 94:16:@38963.4]
  assign RetimeWrapper_15_clock = clock; // @[:@38969.4]
  assign RetimeWrapper_15_reset = reset; // @[:@38970.4]
  assign RetimeWrapper_15_io_flow = 1'h1; // @[package.scala 95:18:@38972.4]
  assign RetimeWrapper_15_io_in = reset; // @[package.scala 94:16:@38971.4]
  assign RetimeWrapper_16_clock = clock; // @[:@38980.4]
  assign RetimeWrapper_16_reset = reset; // @[:@38981.4]
  assign RetimeWrapper_16_io_flow = 1'h1; // @[package.scala 95:18:@38983.4]
  assign RetimeWrapper_16_io_in = _T_162 & _T_167; // @[package.scala 94:16:@38982.4]
  assign RetimeWrapper_17_clock = clock; // @[:@38988.4]
  assign RetimeWrapper_17_reset = reset; // @[:@38989.4]
  assign RetimeWrapper_17_io_flow = 1'h1; // @[package.scala 95:18:@38991.4]
  assign RetimeWrapper_17_io_in = reset; // @[package.scala 94:16:@38990.4]
  assign RetimeWrapper_18_clock = clock; // @[:@38997.4]
  assign RetimeWrapper_18_reset = reset; // @[:@38998.4]
  assign RetimeWrapper_18_io_flow = 1'h1; // @[package.scala 95:18:@39000.4]
  assign RetimeWrapper_18_io_in = _T_162 & _T_167; // @[package.scala 94:16:@38999.4]
  assign RetimeWrapper_19_clock = clock; // @[:@39005.4]
  assign RetimeWrapper_19_reset = reset; // @[:@39006.4]
  assign RetimeWrapper_19_io_flow = 1'h1; // @[package.scala 95:18:@39008.4]
  assign RetimeWrapper_19_io_in = reset; // @[package.scala 94:16:@39007.4]
  assign RetimeWrapper_20_clock = clock; // @[:@39016.4]
  assign RetimeWrapper_20_reset = reset; // @[:@39017.4]
  assign RetimeWrapper_20_io_flow = 1'h1; // @[package.scala 95:18:@39019.4]
  assign RetimeWrapper_20_io_in = _T_162 & _T_167; // @[package.scala 94:16:@39018.4]
  assign RetimeWrapper_21_clock = clock; // @[:@39024.4]
  assign RetimeWrapper_21_reset = reset; // @[:@39025.4]
  assign RetimeWrapper_21_io_flow = 1'h1; // @[package.scala 95:18:@39027.4]
  assign RetimeWrapper_21_io_in = reset; // @[package.scala 94:16:@39026.4]
  assign RetimeWrapper_22_clock = clock; // @[:@39033.4]
  assign RetimeWrapper_22_reset = reset; // @[:@39034.4]
  assign RetimeWrapper_22_io_flow = 1'h1; // @[package.scala 95:18:@39036.4]
  assign RetimeWrapper_22_io_in = _T_162 & _T_167; // @[package.scala 94:16:@39035.4]
  assign RetimeWrapper_23_clock = clock; // @[:@39041.4]
  assign RetimeWrapper_23_reset = reset; // @[:@39042.4]
  assign RetimeWrapper_23_io_flow = 1'h1; // @[package.scala 95:18:@39044.4]
  assign RetimeWrapper_23_io_in = reset; // @[package.scala 94:16:@39043.4]
  assign RetimeWrapper_24_clock = clock; // @[:@39052.4]
  assign RetimeWrapper_24_reset = reset; // @[:@39053.4]
  assign RetimeWrapper_24_io_flow = 1'h1; // @[package.scala 95:18:@39055.4]
  assign RetimeWrapper_24_io_in = _T_162 & _T_167; // @[package.scala 94:16:@39054.4]
  assign RetimeWrapper_25_clock = clock; // @[:@39060.4]
  assign RetimeWrapper_25_reset = reset; // @[:@39061.4]
  assign RetimeWrapper_25_io_flow = 1'h1; // @[package.scala 95:18:@39063.4]
  assign RetimeWrapper_25_io_in = reset; // @[package.scala 94:16:@39062.4]
  assign RetimeWrapper_26_clock = clock; // @[:@39069.4]
  assign RetimeWrapper_26_reset = reset; // @[:@39070.4]
  assign RetimeWrapper_26_io_flow = 1'h1; // @[package.scala 95:18:@39072.4]
  assign RetimeWrapper_26_io_in = _T_162 & _T_167; // @[package.scala 94:16:@39071.4]
  assign RetimeWrapper_27_clock = clock; // @[:@39077.4]
  assign RetimeWrapper_27_reset = reset; // @[:@39078.4]
  assign RetimeWrapper_27_io_flow = 1'h1; // @[package.scala 95:18:@39080.4]
  assign RetimeWrapper_27_io_in = reset; // @[package.scala 94:16:@39079.4]
  assign NBufCtr_clock = clock; // @[:@39118.4]
  assign NBufCtr_reset = reset; // @[:@39119.4]
  assign NBufCtr_io_input_countUp = 1'h0; // @[NBuffers.scala 43:24:@39126.4]
  assign NBufCtr_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 42:23:@39125.4]
  assign NBufCtr_1_clock = clock; // @[:@39129.4]
  assign NBufCtr_1_reset = reset; // @[:@39130.4]
  assign NBufCtr_1_io_input_countUp = 1'h0; // @[NBuffers.scala 43:24:@39137.4]
  assign NBufCtr_1_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 42:23:@39136.4]
  assign statesInR_0_clock = clock; // @[:@39140.4]
  assign statesInR_0_reset = reset; // @[:@39141.4]
  assign statesInR_0_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@39148.4]
  assign statesInR_0_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@39147.4]
  assign statesInR_1_clock = clock; // @[:@39151.4]
  assign statesInR_1_reset = reset; // @[:@39152.4]
  assign statesInR_1_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@39159.4]
  assign statesInR_1_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@39158.4]
  assign statesInR_2_clock = clock; // @[:@39162.4]
  assign statesInR_2_reset = reset; // @[:@39163.4]
  assign statesInR_2_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@39170.4]
  assign statesInR_2_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@39169.4]
  assign statesInR_3_clock = clock; // @[:@39173.4]
  assign statesInR_3_reset = reset; // @[:@39174.4]
  assign statesInR_3_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@39181.4]
  assign statesInR_3_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@39180.4]
  assign statesInR_4_clock = clock; // @[:@39184.4]
  assign statesInR_4_reset = reset; // @[:@39185.4]
  assign statesInR_4_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@39192.4]
  assign statesInR_4_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@39191.4]
  assign statesInR_5_clock = clock; // @[:@39195.4]
  assign statesInR_5_reset = reset; // @[:@39196.4]
  assign statesInR_5_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@39203.4]
  assign statesInR_5_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@39202.4]
  assign statesInR_6_clock = clock; // @[:@39206.4]
  assign statesInR_6_reset = reset; // @[:@39207.4]
  assign statesInR_6_io_input_countUp = 1'h0; // @[NBuffers.scala 53:24:@39214.4]
  assign statesInR_6_io_input_enable = _T_162 & _T_167; // @[NBuffers.scala 52:23:@39213.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_167 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_167 <= 1'h0;
    end else begin
      _T_167 <= _T_164;
    end
  end
endmodule
module x558_tmp_4( // @[:@40785.2]
  input         clock, // @[:@40786.4]
  input         reset, // @[:@40787.4]
  input  [1:0]  io_rPort_0_ofs_0, // @[:@40788.4]
  input         io_rPort_0_en_0, // @[:@40788.4]
  output [31:0] io_rPort_0_output_0, // @[:@40788.4]
  input  [1:0]  io_wPort_1_ofs_0, // @[:@40788.4]
  input  [31:0] io_wPort_1_data_0, // @[:@40788.4]
  input         io_wPort_1_en_0, // @[:@40788.4]
  input  [1:0]  io_wPort_0_ofs_0, // @[:@40788.4]
  input  [31:0] io_wPort_0_data_0, // @[:@40788.4]
  input         io_wPort_0_en_0, // @[:@40788.4]
  input         io_sEn_0, // @[:@40788.4]
  input         io_sEn_1, // @[:@40788.4]
  input         io_sEn_2, // @[:@40788.4]
  input         io_sEn_3, // @[:@40788.4]
  input         io_sEn_4, // @[:@40788.4]
  input         io_sEn_5, // @[:@40788.4]
  input         io_sEn_6, // @[:@40788.4]
  input         io_sDone_0, // @[:@40788.4]
  input         io_sDone_1, // @[:@40788.4]
  input         io_sDone_2, // @[:@40788.4]
  input         io_sDone_3, // @[:@40788.4]
  input         io_sDone_4, // @[:@40788.4]
  input         io_sDone_5, // @[:@40788.4]
  input         io_sDone_6 // @[:@40788.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@40798.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@40798.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@40798.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@40798.4]
  wire  ctrl_io_sEn_2; // @[NBuffers.scala 83:20:@40798.4]
  wire  ctrl_io_sEn_3; // @[NBuffers.scala 83:20:@40798.4]
  wire  ctrl_io_sEn_4; // @[NBuffers.scala 83:20:@40798.4]
  wire  ctrl_io_sEn_5; // @[NBuffers.scala 83:20:@40798.4]
  wire  ctrl_io_sEn_6; // @[NBuffers.scala 83:20:@40798.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@40798.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@40798.4]
  wire  ctrl_io_sDone_2; // @[NBuffers.scala 83:20:@40798.4]
  wire  ctrl_io_sDone_3; // @[NBuffers.scala 83:20:@40798.4]
  wire  ctrl_io_sDone_4; // @[NBuffers.scala 83:20:@40798.4]
  wire  ctrl_io_sDone_5; // @[NBuffers.scala 83:20:@40798.4]
  wire  ctrl_io_sDone_6; // @[NBuffers.scala 83:20:@40798.4]
  wire [3:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@40798.4]
  wire [3:0] ctrl_io_statesInW_1; // @[NBuffers.scala 83:20:@40798.4]
  wire [3:0] ctrl_io_statesInR_6; // @[NBuffers.scala 83:20:@40798.4]
  wire  SRAM_clock; // @[NBuffers.scala 94:23:@40815.4]
  wire  SRAM_reset; // @[NBuffers.scala 94:23:@40815.4]
  wire [1:0] SRAM_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@40815.4]
  wire  SRAM_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@40815.4]
  wire  SRAM_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@40815.4]
  wire [31:0] SRAM_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@40815.4]
  wire [1:0] SRAM_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@40815.4]
  wire [31:0] SRAM_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@40815.4]
  wire  SRAM_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@40815.4]
  wire [1:0] SRAM_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@40815.4]
  wire [31:0] SRAM_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@40815.4]
  wire  SRAM_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@40815.4]
  wire  SRAM_1_clock; // @[NBuffers.scala 94:23:@40838.4]
  wire  SRAM_1_reset; // @[NBuffers.scala 94:23:@40838.4]
  wire [1:0] SRAM_1_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@40838.4]
  wire  SRAM_1_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@40838.4]
  wire  SRAM_1_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@40838.4]
  wire [31:0] SRAM_1_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@40838.4]
  wire [1:0] SRAM_1_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@40838.4]
  wire [31:0] SRAM_1_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@40838.4]
  wire  SRAM_1_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@40838.4]
  wire [1:0] SRAM_1_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@40838.4]
  wire [31:0] SRAM_1_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@40838.4]
  wire  SRAM_1_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@40838.4]
  wire  SRAM_2_clock; // @[NBuffers.scala 94:23:@40861.4]
  wire  SRAM_2_reset; // @[NBuffers.scala 94:23:@40861.4]
  wire [1:0] SRAM_2_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@40861.4]
  wire  SRAM_2_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@40861.4]
  wire  SRAM_2_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@40861.4]
  wire [31:0] SRAM_2_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@40861.4]
  wire [1:0] SRAM_2_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@40861.4]
  wire [31:0] SRAM_2_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@40861.4]
  wire  SRAM_2_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@40861.4]
  wire [1:0] SRAM_2_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@40861.4]
  wire [31:0] SRAM_2_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@40861.4]
  wire  SRAM_2_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@40861.4]
  wire  SRAM_3_clock; // @[NBuffers.scala 94:23:@40884.4]
  wire  SRAM_3_reset; // @[NBuffers.scala 94:23:@40884.4]
  wire [1:0] SRAM_3_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@40884.4]
  wire  SRAM_3_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@40884.4]
  wire  SRAM_3_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@40884.4]
  wire [31:0] SRAM_3_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@40884.4]
  wire [1:0] SRAM_3_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@40884.4]
  wire [31:0] SRAM_3_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@40884.4]
  wire  SRAM_3_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@40884.4]
  wire [1:0] SRAM_3_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@40884.4]
  wire [31:0] SRAM_3_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@40884.4]
  wire  SRAM_3_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@40884.4]
  wire  SRAM_4_clock; // @[NBuffers.scala 94:23:@40907.4]
  wire  SRAM_4_reset; // @[NBuffers.scala 94:23:@40907.4]
  wire [1:0] SRAM_4_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@40907.4]
  wire  SRAM_4_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@40907.4]
  wire  SRAM_4_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@40907.4]
  wire [31:0] SRAM_4_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@40907.4]
  wire [1:0] SRAM_4_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@40907.4]
  wire [31:0] SRAM_4_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@40907.4]
  wire  SRAM_4_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@40907.4]
  wire [1:0] SRAM_4_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@40907.4]
  wire [31:0] SRAM_4_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@40907.4]
  wire  SRAM_4_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@40907.4]
  wire  SRAM_5_clock; // @[NBuffers.scala 94:23:@40930.4]
  wire  SRAM_5_reset; // @[NBuffers.scala 94:23:@40930.4]
  wire [1:0] SRAM_5_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@40930.4]
  wire  SRAM_5_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@40930.4]
  wire  SRAM_5_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@40930.4]
  wire [31:0] SRAM_5_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@40930.4]
  wire [1:0] SRAM_5_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@40930.4]
  wire [31:0] SRAM_5_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@40930.4]
  wire  SRAM_5_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@40930.4]
  wire [1:0] SRAM_5_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@40930.4]
  wire [31:0] SRAM_5_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@40930.4]
  wire  SRAM_5_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@40930.4]
  wire  SRAM_6_clock; // @[NBuffers.scala 94:23:@40953.4]
  wire  SRAM_6_reset; // @[NBuffers.scala 94:23:@40953.4]
  wire [1:0] SRAM_6_io_rPort_0_ofs_0; // @[NBuffers.scala 94:23:@40953.4]
  wire  SRAM_6_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@40953.4]
  wire  SRAM_6_io_rPort_0_backpressure; // @[NBuffers.scala 94:23:@40953.4]
  wire [31:0] SRAM_6_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@40953.4]
  wire [1:0] SRAM_6_io_wPort_1_ofs_0; // @[NBuffers.scala 94:23:@40953.4]
  wire [31:0] SRAM_6_io_wPort_1_data_0; // @[NBuffers.scala 94:23:@40953.4]
  wire  SRAM_6_io_wPort_1_en_0; // @[NBuffers.scala 94:23:@40953.4]
  wire [1:0] SRAM_6_io_wPort_0_ofs_0; // @[NBuffers.scala 94:23:@40953.4]
  wire [31:0] SRAM_6_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@40953.4]
  wire  SRAM_6_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@40953.4]
  wire  _T_148; // @[NBuffers.scala 104:105:@40976.4]
  wire  _T_152; // @[NBuffers.scala 104:105:@40986.4]
  wire  _T_156; // @[NBuffers.scala 108:92:@40996.4]
  wire  _T_159; // @[NBuffers.scala 104:105:@41002.4]
  wire  _T_163; // @[NBuffers.scala 104:105:@41012.4]
  wire  _T_167; // @[NBuffers.scala 108:92:@41022.4]
  wire  _T_170; // @[NBuffers.scala 104:105:@41028.4]
  wire  _T_174; // @[NBuffers.scala 104:105:@41038.4]
  wire  _T_178; // @[NBuffers.scala 108:92:@41048.4]
  wire  _T_181; // @[NBuffers.scala 104:105:@41054.4]
  wire  _T_185; // @[NBuffers.scala 104:105:@41064.4]
  wire  _T_189; // @[NBuffers.scala 108:92:@41074.4]
  wire  _T_192; // @[NBuffers.scala 104:105:@41080.4]
  wire  _T_196; // @[NBuffers.scala 104:105:@41090.4]
  wire  _T_200; // @[NBuffers.scala 108:92:@41100.4]
  wire  _T_203; // @[NBuffers.scala 104:105:@41106.4]
  wire  _T_207; // @[NBuffers.scala 104:105:@41116.4]
  wire  _T_211; // @[NBuffers.scala 108:92:@41126.4]
  wire  _T_214; // @[NBuffers.scala 104:105:@41132.4]
  wire  _T_218; // @[NBuffers.scala 104:105:@41142.4]
  wire  _T_222; // @[NBuffers.scala 108:92:@41152.4]
  wire [31:0] _T_240; // @[Mux.scala 19:72:@41165.4]
  wire [31:0] _T_242; // @[Mux.scala 19:72:@41166.4]
  wire [31:0] _T_244; // @[Mux.scala 19:72:@41167.4]
  wire [31:0] _T_246; // @[Mux.scala 19:72:@41168.4]
  wire [31:0] _T_248; // @[Mux.scala 19:72:@41169.4]
  wire [31:0] _T_250; // @[Mux.scala 19:72:@41170.4]
  wire [31:0] _T_252; // @[Mux.scala 19:72:@41171.4]
  wire [31:0] _T_253; // @[Mux.scala 19:72:@41172.4]
  wire [31:0] _T_254; // @[Mux.scala 19:72:@41173.4]
  wire [31:0] _T_255; // @[Mux.scala 19:72:@41174.4]
  wire [31:0] _T_256; // @[Mux.scala 19:72:@41175.4]
  wire [31:0] _T_257; // @[Mux.scala 19:72:@41176.4]
  NBufController_9 ctrl ( // @[NBuffers.scala 83:20:@40798.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sEn_2(ctrl_io_sEn_2),
    .io_sEn_3(ctrl_io_sEn_3),
    .io_sEn_4(ctrl_io_sEn_4),
    .io_sEn_5(ctrl_io_sEn_5),
    .io_sEn_6(ctrl_io_sEn_6),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_sDone_2(ctrl_io_sDone_2),
    .io_sDone_3(ctrl_io_sDone_3),
    .io_sDone_4(ctrl_io_sDone_4),
    .io_sDone_5(ctrl_io_sDone_5),
    .io_sDone_6(ctrl_io_sDone_6),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInW_1(ctrl_io_statesInW_1),
    .io_statesInR_6(ctrl_io_statesInR_6)
  );
  SRAM_10 SRAM ( // @[NBuffers.scala 94:23:@40815.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_rPort_0_ofs_0(SRAM_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_1 ( // @[NBuffers.scala 94:23:@40838.4]
    .clock(SRAM_1_clock),
    .reset(SRAM_1_reset),
    .io_rPort_0_ofs_0(SRAM_1_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_1_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_1_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_1_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_1_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_1_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_1_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_1_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_1_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_2 ( // @[NBuffers.scala 94:23:@40861.4]
    .clock(SRAM_2_clock),
    .reset(SRAM_2_reset),
    .io_rPort_0_ofs_0(SRAM_2_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_2_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_2_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_2_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_2_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_2_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_2_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_2_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_2_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_2_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_3 ( // @[NBuffers.scala 94:23:@40884.4]
    .clock(SRAM_3_clock),
    .reset(SRAM_3_reset),
    .io_rPort_0_ofs_0(SRAM_3_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_3_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_3_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_3_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_3_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_3_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_3_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_3_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_3_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_3_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_4 ( // @[NBuffers.scala 94:23:@40907.4]
    .clock(SRAM_4_clock),
    .reset(SRAM_4_reset),
    .io_rPort_0_ofs_0(SRAM_4_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_4_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_4_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_4_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_4_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_4_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_4_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_4_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_4_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_4_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_5 ( // @[NBuffers.scala 94:23:@40930.4]
    .clock(SRAM_5_clock),
    .reset(SRAM_5_reset),
    .io_rPort_0_ofs_0(SRAM_5_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_5_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_5_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_5_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_5_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_5_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_5_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_5_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_5_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_5_io_wPort_0_en_0)
  );
  SRAM_10 SRAM_6 ( // @[NBuffers.scala 94:23:@40953.4]
    .clock(SRAM_6_clock),
    .reset(SRAM_6_reset),
    .io_rPort_0_ofs_0(SRAM_6_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(SRAM_6_io_rPort_0_en_0),
    .io_rPort_0_backpressure(SRAM_6_io_rPort_0_backpressure),
    .io_rPort_0_output_0(SRAM_6_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(SRAM_6_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(SRAM_6_io_wPort_1_data_0),
    .io_wPort_1_en_0(SRAM_6_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(SRAM_6_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(SRAM_6_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_6_io_wPort_0_en_0)
  );
  assign _T_148 = ctrl_io_statesInW_0 == 4'h0; // @[NBuffers.scala 104:105:@40976.4]
  assign _T_152 = ctrl_io_statesInW_1 == 4'h0; // @[NBuffers.scala 104:105:@40986.4]
  assign _T_156 = ctrl_io_statesInR_6 == 4'h0; // @[NBuffers.scala 108:92:@40996.4]
  assign _T_159 = ctrl_io_statesInW_0 == 4'h1; // @[NBuffers.scala 104:105:@41002.4]
  assign _T_163 = ctrl_io_statesInW_1 == 4'h1; // @[NBuffers.scala 104:105:@41012.4]
  assign _T_167 = ctrl_io_statesInR_6 == 4'h1; // @[NBuffers.scala 108:92:@41022.4]
  assign _T_170 = ctrl_io_statesInW_0 == 4'h2; // @[NBuffers.scala 104:105:@41028.4]
  assign _T_174 = ctrl_io_statesInW_1 == 4'h2; // @[NBuffers.scala 104:105:@41038.4]
  assign _T_178 = ctrl_io_statesInR_6 == 4'h2; // @[NBuffers.scala 108:92:@41048.4]
  assign _T_181 = ctrl_io_statesInW_0 == 4'h3; // @[NBuffers.scala 104:105:@41054.4]
  assign _T_185 = ctrl_io_statesInW_1 == 4'h3; // @[NBuffers.scala 104:105:@41064.4]
  assign _T_189 = ctrl_io_statesInR_6 == 4'h3; // @[NBuffers.scala 108:92:@41074.4]
  assign _T_192 = ctrl_io_statesInW_0 == 4'h4; // @[NBuffers.scala 104:105:@41080.4]
  assign _T_196 = ctrl_io_statesInW_1 == 4'h4; // @[NBuffers.scala 104:105:@41090.4]
  assign _T_200 = ctrl_io_statesInR_6 == 4'h4; // @[NBuffers.scala 108:92:@41100.4]
  assign _T_203 = ctrl_io_statesInW_0 == 4'h5; // @[NBuffers.scala 104:105:@41106.4]
  assign _T_207 = ctrl_io_statesInW_1 == 4'h5; // @[NBuffers.scala 104:105:@41116.4]
  assign _T_211 = ctrl_io_statesInR_6 == 4'h5; // @[NBuffers.scala 108:92:@41126.4]
  assign _T_214 = ctrl_io_statesInW_0 == 4'h6; // @[NBuffers.scala 104:105:@41132.4]
  assign _T_218 = ctrl_io_statesInW_1 == 4'h6; // @[NBuffers.scala 104:105:@41142.4]
  assign _T_222 = ctrl_io_statesInR_6 == 4'h6; // @[NBuffers.scala 108:92:@41152.4]
  assign _T_240 = _T_156 ? SRAM_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@41165.4]
  assign _T_242 = _T_167 ? SRAM_1_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@41166.4]
  assign _T_244 = _T_178 ? SRAM_2_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@41167.4]
  assign _T_246 = _T_189 ? SRAM_3_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@41168.4]
  assign _T_248 = _T_200 ? SRAM_4_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@41169.4]
  assign _T_250 = _T_211 ? SRAM_5_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@41170.4]
  assign _T_252 = _T_222 ? SRAM_6_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@41171.4]
  assign _T_253 = _T_240 | _T_242; // @[Mux.scala 19:72:@41172.4]
  assign _T_254 = _T_253 | _T_244; // @[Mux.scala 19:72:@41173.4]
  assign _T_255 = _T_254 | _T_246; // @[Mux.scala 19:72:@41174.4]
  assign _T_256 = _T_255 | _T_248; // @[Mux.scala 19:72:@41175.4]
  assign _T_257 = _T_256 | _T_250; // @[Mux.scala 19:72:@41176.4]
  assign io_rPort_0_output_0 = _T_257 | _T_252; // @[NBuffers.scala 115:66:@41180.4]
  assign ctrl_clock = clock; // @[:@40799.4]
  assign ctrl_reset = reset; // @[:@40800.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@40801.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@40803.4]
  assign ctrl_io_sEn_2 = io_sEn_2; // @[NBuffers.scala 85:20:@40805.4]
  assign ctrl_io_sEn_3 = io_sEn_3; // @[NBuffers.scala 85:20:@40807.4]
  assign ctrl_io_sEn_4 = io_sEn_4; // @[NBuffers.scala 85:20:@40809.4]
  assign ctrl_io_sEn_5 = io_sEn_5; // @[NBuffers.scala 85:20:@40811.4]
  assign ctrl_io_sEn_6 = io_sEn_6; // @[NBuffers.scala 85:20:@40813.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@40802.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@40804.4]
  assign ctrl_io_sDone_2 = io_sDone_2; // @[NBuffers.scala 86:22:@40806.4]
  assign ctrl_io_sDone_3 = io_sDone_3; // @[NBuffers.scala 86:22:@40808.4]
  assign ctrl_io_sDone_4 = io_sDone_4; // @[NBuffers.scala 86:22:@40810.4]
  assign ctrl_io_sDone_5 = io_sDone_5; // @[NBuffers.scala 86:22:@40812.4]
  assign ctrl_io_sDone_6 = io_sDone_6; // @[NBuffers.scala 86:22:@40814.4]
  assign SRAM_clock = clock; // @[:@40816.4]
  assign SRAM_reset = reset; // @[:@40817.4]
  assign SRAM_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@40998.4]
  assign SRAM_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_156; // @[MemPrimitives.scala 43:33:@41000.4]
  assign SRAM_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@41001.4]
  assign SRAM_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@40988.4]
  assign SRAM_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@40989.4]
  assign SRAM_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_152; // @[MemPrimitives.scala 37:29:@40995.4]
  assign SRAM_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@40978.4]
  assign SRAM_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@40979.4]
  assign SRAM_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_148; // @[MemPrimitives.scala 37:29:@40985.4]
  assign SRAM_1_clock = clock; // @[:@40839.4]
  assign SRAM_1_reset = reset; // @[:@40840.4]
  assign SRAM_1_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@41024.4]
  assign SRAM_1_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_167; // @[MemPrimitives.scala 43:33:@41026.4]
  assign SRAM_1_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@41027.4]
  assign SRAM_1_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@41014.4]
  assign SRAM_1_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@41015.4]
  assign SRAM_1_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_163; // @[MemPrimitives.scala 37:29:@41021.4]
  assign SRAM_1_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@41004.4]
  assign SRAM_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@41005.4]
  assign SRAM_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_159; // @[MemPrimitives.scala 37:29:@41011.4]
  assign SRAM_2_clock = clock; // @[:@40862.4]
  assign SRAM_2_reset = reset; // @[:@40863.4]
  assign SRAM_2_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@41050.4]
  assign SRAM_2_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_178; // @[MemPrimitives.scala 43:33:@41052.4]
  assign SRAM_2_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@41053.4]
  assign SRAM_2_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@41040.4]
  assign SRAM_2_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@41041.4]
  assign SRAM_2_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_174; // @[MemPrimitives.scala 37:29:@41047.4]
  assign SRAM_2_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@41030.4]
  assign SRAM_2_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@41031.4]
  assign SRAM_2_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_170; // @[MemPrimitives.scala 37:29:@41037.4]
  assign SRAM_3_clock = clock; // @[:@40885.4]
  assign SRAM_3_reset = reset; // @[:@40886.4]
  assign SRAM_3_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@41076.4]
  assign SRAM_3_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_189; // @[MemPrimitives.scala 43:33:@41078.4]
  assign SRAM_3_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@41079.4]
  assign SRAM_3_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@41066.4]
  assign SRAM_3_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@41067.4]
  assign SRAM_3_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_185; // @[MemPrimitives.scala 37:29:@41073.4]
  assign SRAM_3_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@41056.4]
  assign SRAM_3_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@41057.4]
  assign SRAM_3_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_181; // @[MemPrimitives.scala 37:29:@41063.4]
  assign SRAM_4_clock = clock; // @[:@40908.4]
  assign SRAM_4_reset = reset; // @[:@40909.4]
  assign SRAM_4_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@41102.4]
  assign SRAM_4_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_200; // @[MemPrimitives.scala 43:33:@41104.4]
  assign SRAM_4_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@41105.4]
  assign SRAM_4_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@41092.4]
  assign SRAM_4_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@41093.4]
  assign SRAM_4_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_196; // @[MemPrimitives.scala 37:29:@41099.4]
  assign SRAM_4_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@41082.4]
  assign SRAM_4_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@41083.4]
  assign SRAM_4_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_192; // @[MemPrimitives.scala 37:29:@41089.4]
  assign SRAM_5_clock = clock; // @[:@40931.4]
  assign SRAM_5_reset = reset; // @[:@40932.4]
  assign SRAM_5_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@41128.4]
  assign SRAM_5_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_211; // @[MemPrimitives.scala 43:33:@41130.4]
  assign SRAM_5_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@41131.4]
  assign SRAM_5_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@41118.4]
  assign SRAM_5_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@41119.4]
  assign SRAM_5_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_207; // @[MemPrimitives.scala 37:29:@41125.4]
  assign SRAM_5_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@41108.4]
  assign SRAM_5_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@41109.4]
  assign SRAM_5_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_203; // @[MemPrimitives.scala 37:29:@41115.4]
  assign SRAM_6_clock = clock; // @[:@40954.4]
  assign SRAM_6_reset = reset; // @[:@40955.4]
  assign SRAM_6_io_rPort_0_ofs_0 = io_rPort_0_ofs_0; // @[MemPrimitives.scala 42:33:@41154.4]
  assign SRAM_6_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_222; // @[MemPrimitives.scala 43:33:@41156.4]
  assign SRAM_6_io_rPort_0_backpressure = 1'h1; // @[MemPrimitives.scala 44:33:@41157.4]
  assign SRAM_6_io_wPort_1_ofs_0 = io_wPort_1_ofs_0; // @[MemPrimitives.scala 32:29:@41144.4]
  assign SRAM_6_io_wPort_1_data_0 = io_wPort_1_data_0; // @[MemPrimitives.scala 33:29:@41145.4]
  assign SRAM_6_io_wPort_1_en_0 = io_wPort_1_en_0 & _T_218; // @[MemPrimitives.scala 37:29:@41151.4]
  assign SRAM_6_io_wPort_0_ofs_0 = io_wPort_0_ofs_0; // @[MemPrimitives.scala 32:29:@41134.4]
  assign SRAM_6_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@41135.4]
  assign SRAM_6_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_214; // @[MemPrimitives.scala 37:29:@41141.4]
endmodule
module RetimeWrapper_451( // @[:@41383.2]
  input   clock, // @[:@41384.4]
  input   reset, // @[:@41385.4]
  input   io_flow, // @[:@41386.4]
  input   io_in, // @[:@41386.4]
  output  io_out // @[:@41386.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@41388.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@41388.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@41388.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@41388.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@41388.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@41388.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@41388.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@41401.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@41400.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@41399.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@41398.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@41397.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@41395.4]
endmodule
module x579_inr_Foreach_sm( // @[:@41531.2]
  input   clock, // @[:@41532.4]
  input   reset, // @[:@41533.4]
  input   io_enable, // @[:@41534.4]
  output  io_done, // @[:@41534.4]
  input   io_ctrDone, // @[:@41534.4]
  output  io_datapathEn, // @[:@41534.4]
  output  io_ctrInc, // @[:@41534.4]
  output  io_ctrRst, // @[:@41534.4]
  input   io_parentAck, // @[:@41534.4]
  input   io_backpressure, // @[:@41534.4]
  input   io_break // @[:@41534.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@41536.4]
  wire  active_reset; // @[Controllers.scala 261:22:@41536.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@41536.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@41536.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@41536.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@41536.4]
  wire  done_clock; // @[Controllers.scala 262:20:@41539.4]
  wire  done_reset; // @[Controllers.scala 262:20:@41539.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@41539.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@41539.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@41539.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@41539.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@41573.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@41573.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@41573.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@41573.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@41573.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@41595.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@41595.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@41595.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@41595.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@41595.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@41607.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@41607.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@41607.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@41607.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@41607.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@41615.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@41615.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@41615.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@41615.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@41615.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@41631.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@41631.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@41631.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@41631.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@41631.4]
  wire  _T_80; // @[Controllers.scala 264:48:@41544.4]
  wire  _T_81; // @[Controllers.scala 264:46:@41545.4]
  wire  _T_82; // @[Controllers.scala 264:62:@41546.4]
  wire  _T_100; // @[package.scala 100:49:@41564.4]
  reg  _T_103; // @[package.scala 48:56:@41565.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@41578.4 package.scala 96:25:@41579.4]
  wire  _T_110; // @[package.scala 100:49:@41580.4]
  reg  _T_113; // @[package.scala 48:56:@41581.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@41583.4]
  wire  _T_118; // @[Controllers.scala 283:41:@41588.4]
  wire  _T_124; // @[package.scala 96:25:@41600.4 package.scala 96:25:@41601.4]
  wire  _T_126; // @[package.scala 100:49:@41602.4]
  reg  _T_129; // @[package.scala 48:56:@41603.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@41627.4]
  reg  _T_153; // @[package.scala 48:56:@41628.4]
  reg [31:0] _RAND_3;
  SRFF active ( // @[Controllers.scala 261:22:@41536.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@41539.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_451 RetimeWrapper ( // @[package.scala 93:22:@41573.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_451 RetimeWrapper_1 ( // @[package.scala 93:22:@41595.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@41607.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@41615.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_4 ( // @[package.scala 93:22:@41631.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@41544.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@41545.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@41546.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@41564.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@41578.4 package.scala 96:25:@41579.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@41580.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@41583.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@41588.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@41600.4 package.scala 96:25:@41601.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@41602.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@41627.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@41606.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@41591.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@41594.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@41586.4]
  assign active_clock = clock; // @[:@41537.4]
  assign active_reset = reset; // @[:@41538.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@41549.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@41553.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@41554.4]
  assign done_clock = clock; // @[:@41540.4]
  assign done_reset = reset; // @[:@41541.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@41569.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@41562.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@41563.4]
  assign RetimeWrapper_clock = clock; // @[:@41574.4]
  assign RetimeWrapper_reset = reset; // @[:@41575.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@41577.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@41576.4]
  assign RetimeWrapper_1_clock = clock; // @[:@41596.4]
  assign RetimeWrapper_1_reset = reset; // @[:@41597.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@41599.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@41598.4]
  assign RetimeWrapper_2_clock = clock; // @[:@41608.4]
  assign RetimeWrapper_2_reset = reset; // @[:@41609.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@41611.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@41610.4]
  assign RetimeWrapper_3_clock = clock; // @[:@41616.4]
  assign RetimeWrapper_3_reset = reset; // @[:@41617.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@41619.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@41618.4]
  assign RetimeWrapper_4_clock = clock; // @[:@41632.4]
  assign RetimeWrapper_4_reset = reset; // @[:@41633.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@41635.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@41634.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox_50( // @[:@42820.2]
  input  [31:0] io_a, // @[:@42823.4]
  output [32:0] io_b // @[:@42823.4]
);
  wire [21:0] tmp_frac; // @[Converter.scala 52:23:@42831.4]
  wire  _T_19; // @[implicits.scala 70:16:@42833.4]
  wire [9:0] _T_20; // @[Converter.scala 84:75:@42835.4]
  wire [10:0] new_dec; // @[Cat.scala 30:58:@42836.4]
  assign tmp_frac = io_a[21:0]; // @[Converter.scala 52:23:@42831.4]
  assign _T_19 = io_a[31]; // @[implicits.scala 70:16:@42833.4]
  assign _T_20 = io_a[31:22]; // @[Converter.scala 84:75:@42835.4]
  assign new_dec = {_T_19,_T_20}; // @[Cat.scala 30:58:@42836.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@42839.4]
endmodule
module __37( // @[:@42841.2]
  input  [31:0] io_b, // @[:@42844.4]
  output [32:0] io_result // @[:@42844.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@42849.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@42849.4]
  fix2fixBox_50 fix2fixBox ( // @[BigIPZynq.scala 219:30:@42849.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@42857.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@42852.4]
endmodule
module fix2fixBox_52( // @[:@42930.2]
  input         clock, // @[:@42931.4]
  input         reset, // @[:@42932.4]
  input  [32:0] io_a, // @[:@42933.4]
  input         io_flow, // @[:@42933.4]
  output [31:0] io_b // @[:@42933.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@42947.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@42947.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@42947.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@42947.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@42947.4]
  wire [21:0] tmp_frac; // @[Converter.scala 52:23:@42941.4]
  wire [9:0] new_dec; // @[Converter.scala 63:26:@42944.4]
  RetimeWrapper_31 RetimeWrapper ( // @[package.scala 93:22:@42947.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign tmp_frac = io_a[21:0]; // @[Converter.scala 52:23:@42941.4]
  assign new_dec = io_a[31:22]; // @[Converter.scala 63:26:@42944.4]
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 94:38:@42954.4]
  assign RetimeWrapper_clock = clock; // @[:@42948.4]
  assign RetimeWrapper_reset = reset; // @[:@42949.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@42951.4]
  assign RetimeWrapper_io_in = {new_dec,tmp_frac}; // @[package.scala 94:16:@42950.4]
endmodule
module x573_sub( // @[:@42956.2]
  input         clock, // @[:@42957.4]
  input         reset, // @[:@42958.4]
  input  [31:0] io_a, // @[:@42959.4]
  input  [31:0] io_b, // @[:@42959.4]
  output [31:0] io_result // @[:@42959.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@42967.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@42967.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@42974.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@42974.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@42993.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@42993.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@42993.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@42993.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@42993.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@42972.4 Math.scala 724:14:@42973.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@42979.4 Math.scala 724:14:@42980.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@42981.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@42982.4]
  __37 _ ( // @[Math.scala 720:24:@42967.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __37 __1 ( // @[Math.scala 720:24:@42974.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_52 fix2fixBox ( // @[Math.scala 182:30:@42993.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@42972.4 Math.scala 724:14:@42973.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@42979.4 Math.scala 724:14:@42980.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@42981.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@42982.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@43001.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@42970.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@42977.4]
  assign fix2fixBox_clock = clock; // @[:@42994.4]
  assign fix2fixBox_reset = reset; // @[:@42995.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@42996.4]
  assign fix2fixBox_io_flow = 1'h1; // @[Math.scala 186:26:@42999.4]
endmodule
module RetimeWrapper_474( // @[:@43015.2]
  input         clock, // @[:@43016.4]
  input         reset, // @[:@43017.4]
  input  [31:0] io_in, // @[:@43018.4]
  output [31:0] io_out // @[:@43018.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@43020.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@43020.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@43020.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@43020.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@43020.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@43020.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@43020.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@43033.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@43032.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@43031.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@43030.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@43029.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@43027.4]
endmodule
module x579_inr_Foreach_kernelx579_inr_Foreach_concrete1( // @[:@43451.2]
  input         clock, // @[:@43452.4]
  input         reset, // @[:@43453.4]
  output [1:0]  io_in_x555_tmp_1_wPort_0_ofs_0, // @[:@43454.4]
  output [31:0] io_in_x555_tmp_1_wPort_0_data_0, // @[:@43454.4]
  output        io_in_x555_tmp_1_wPort_0_en_0, // @[:@43454.4]
  output        io_in_x555_tmp_1_sEn_0, // @[:@43454.4]
  output        io_in_x555_tmp_1_sDone_0, // @[:@43454.4]
  input  [31:0] io_in_b550_number, // @[:@43454.4]
  output [8:0]  io_in_x472_A_sram_1_rPort_0_ofs_0, // @[:@43454.4]
  output        io_in_x472_A_sram_1_rPort_0_en_0, // @[:@43454.4]
  input  [31:0] io_in_x472_A_sram_1_rPort_0_output_0, // @[:@43454.4]
  input  [31:0] io_in_b542_number, // @[:@43454.4]
  output [8:0]  io_in_x471_A_sram_0_rPort_0_ofs_0, // @[:@43454.4]
  output        io_in_x471_A_sram_0_rPort_0_en_0, // @[:@43454.4]
  input  [31:0] io_in_x471_A_sram_0_rPort_0_output_0, // @[:@43454.4]
  output [1:0]  io_in_x554_tmp_0_wPort_0_ofs_0, // @[:@43454.4]
  output [31:0] io_in_x554_tmp_0_wPort_0_data_0, // @[:@43454.4]
  output        io_in_x554_tmp_0_wPort_0_en_0, // @[:@43454.4]
  output        io_in_x554_tmp_0_sEn_0, // @[:@43454.4]
  output        io_in_x554_tmp_0_sDone_0, // @[:@43454.4]
  output [1:0]  io_in_x558_tmp_4_wPort_0_ofs_0, // @[:@43454.4]
  output [31:0] io_in_x558_tmp_4_wPort_0_data_0, // @[:@43454.4]
  output        io_in_x558_tmp_4_wPort_0_en_0, // @[:@43454.4]
  output        io_in_x558_tmp_4_sEn_0, // @[:@43454.4]
  output        io_in_x558_tmp_4_sDone_0, // @[:@43454.4]
  input         io_in_b552, // @[:@43454.4]
  output [1:0]  io_in_x557_tmp_3_wPort_0_ofs_0, // @[:@43454.4]
  output [31:0] io_in_x557_tmp_3_wPort_0_data_0, // @[:@43454.4]
  output        io_in_x557_tmp_3_wPort_0_en_0, // @[:@43454.4]
  output        io_in_x557_tmp_3_sEn_0, // @[:@43454.4]
  output        io_in_x557_tmp_3_sDone_0, // @[:@43454.4]
  output [1:0]  io_in_x556_tmp_2_wPort_0_ofs_0, // @[:@43454.4]
  output [31:0] io_in_x556_tmp_2_wPort_0_data_0, // @[:@43454.4]
  output        io_in_x556_tmp_2_wPort_0_en_0, // @[:@43454.4]
  output        io_in_x556_tmp_2_sEn_0, // @[:@43454.4]
  output        io_in_x556_tmp_2_sDone_0, // @[:@43454.4]
  input         io_in_b543, // @[:@43454.4]
  input         io_sigsIn_done, // @[:@43454.4]
  input         io_sigsIn_datapathEn, // @[:@43454.4]
  input         io_sigsIn_baseEn, // @[:@43454.4]
  input         io_sigsIn_break, // @[:@43454.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@43454.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@43454.4]
  input         io_rr // @[:@43454.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@43711.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@43711.4]
  wire  x745_sum_1_clock; // @[Math.scala 150:24:@43726.4]
  wire  x745_sum_1_reset; // @[Math.scala 150:24:@43726.4]
  wire [31:0] x745_sum_1_io_a; // @[Math.scala 150:24:@43726.4]
  wire [31:0] x745_sum_1_io_b; // @[Math.scala 150:24:@43726.4]
  wire  x745_sum_1_io_flow; // @[Math.scala 150:24:@43726.4]
  wire [31:0] x745_sum_1_io_result; // @[Math.scala 150:24:@43726.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@43737.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@43737.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@43737.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@43737.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@43737.4]
  wire  x565_sum_1_clock; // @[Math.scala 150:24:@43746.4]
  wire  x565_sum_1_reset; // @[Math.scala 150:24:@43746.4]
  wire [31:0] x565_sum_1_io_a; // @[Math.scala 150:24:@43746.4]
  wire [31:0] x565_sum_1_io_b; // @[Math.scala 150:24:@43746.4]
  wire  x565_sum_1_io_flow; // @[Math.scala 150:24:@43746.4]
  wire [31:0] x565_sum_1_io_result; // @[Math.scala 150:24:@43746.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@43757.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@43757.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@43757.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@43757.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@43757.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@43767.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@43767.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@43767.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@43767.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@43767.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@43777.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@43777.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@43777.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@43777.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@43777.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@43789.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@43789.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@43789.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@43789.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@43789.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@43801.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@43801.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@43801.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@43801.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@43801.4]
  wire  x747_sum_1_clock; // @[Math.scala 150:24:@43827.4]
  wire  x747_sum_1_reset; // @[Math.scala 150:24:@43827.4]
  wire [31:0] x747_sum_1_io_a; // @[Math.scala 150:24:@43827.4]
  wire [31:0] x747_sum_1_io_b; // @[Math.scala 150:24:@43827.4]
  wire  x747_sum_1_io_flow; // @[Math.scala 150:24:@43827.4]
  wire [31:0] x747_sum_1_io_result; // @[Math.scala 150:24:@43827.4]
  wire  x570_sum_1_clock; // @[Math.scala 150:24:@43837.4]
  wire  x570_sum_1_reset; // @[Math.scala 150:24:@43837.4]
  wire [31:0] x570_sum_1_io_a; // @[Math.scala 150:24:@43837.4]
  wire [31:0] x570_sum_1_io_b; // @[Math.scala 150:24:@43837.4]
  wire  x570_sum_1_io_flow; // @[Math.scala 150:24:@43837.4]
  wire [31:0] x570_sum_1_io_result; // @[Math.scala 150:24:@43837.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@43850.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@43850.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@43850.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@43850.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@43850.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@43862.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@43862.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@43862.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@43862.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@43862.4]
  wire  x573_sub_1_clock; // @[Math.scala 191:24:@43883.4]
  wire  x573_sub_1_reset; // @[Math.scala 191:24:@43883.4]
  wire [31:0] x573_sub_1_io_a; // @[Math.scala 191:24:@43883.4]
  wire [31:0] x573_sub_1_io_b; // @[Math.scala 191:24:@43883.4]
  wire [31:0] x573_sub_1_io_result; // @[Math.scala 191:24:@43883.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@43894.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@43894.4]
  wire [31:0] RetimeWrapper_8_io_in; // @[package.scala 93:22:@43894.4]
  wire [31:0] RetimeWrapper_8_io_out; // @[package.scala 93:22:@43894.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@43904.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@43904.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@43904.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@43904.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@43904.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@43914.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@43914.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@43914.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@43914.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@43914.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@43924.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@43924.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@43924.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@43924.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@43924.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@43938.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@43938.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@43938.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@43938.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@43938.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@43964.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@43964.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@43964.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@43964.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@43964.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@43990.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@43990.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@43990.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@43990.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@43990.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@44016.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@44016.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@44016.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@44016.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@44016.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@44042.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@44042.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@44042.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@44042.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@44042.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@44063.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@44063.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@44063.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@44063.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@44063.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@44074.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@44074.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@44074.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@44074.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@44074.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@44085.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@44085.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@44085.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@44085.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@44085.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@44096.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@44096.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@44096.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@44096.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@44096.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@44107.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@44107.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@44107.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@44107.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@44107.4]
  wire [32:0] _GEN_0; // @[Math.scala 461:32:@43722.4]
  wire [32:0] _T_1817; // @[Math.scala 461:32:@43722.4]
  wire  _T_1859; // @[package.scala 96:25:@43794.4 package.scala 96:25:@43795.4]
  wire  _T_1861; // @[implicits.scala 56:10:@43796.4]
  wire  _T_1862; // @[sm_x579_inr_Foreach.scala 119:114:@43797.4]
  wire  _T_1863; // @[sm_x579_inr_Foreach.scala 119:111:@43798.4]
  wire  _T_1868; // @[package.scala 96:25:@43806.4 package.scala 96:25:@43807.4]
  wire  _T_1870; // @[implicits.scala 56:10:@43808.4]
  wire  _T_1871; // @[sm_x579_inr_Foreach.scala 119:131:@43809.4]
  wire  x772_b562_D2; // @[package.scala 96:25:@43782.4 package.scala 96:25:@43783.4]
  wire  _T_1872; // @[sm_x579_inr_Foreach.scala 119:228:@43810.4]
  wire  x771_b552_D2; // @[package.scala 96:25:@43772.4 package.scala 96:25:@43773.4]
  wire  _T_1873; // @[sm_x579_inr_Foreach.scala 119:236:@43811.4]
  wire  x770_b543_D2; // @[package.scala 96:25:@43762.4 package.scala 96:25:@43763.4]
  wire [32:0] _GEN_1; // @[Math.scala 461:32:@43823.4]
  wire [32:0] _T_1879; // @[Math.scala 461:32:@43823.4]
  wire  _T_1901; // @[package.scala 96:25:@43855.4 package.scala 96:25:@43856.4]
  wire  _T_1903; // @[implicits.scala 56:10:@43857.4]
  wire  _T_1905; // @[sm_x579_inr_Foreach.scala 134:111:@43859.4]
  wire  _T_1910; // @[package.scala 96:25:@43867.4 package.scala 96:25:@43868.4]
  wire  _T_1912; // @[implicits.scala 56:10:@43869.4]
  wire  _T_1913; // @[sm_x579_inr_Foreach.scala 134:131:@43870.4]
  wire  _T_1914; // @[sm_x579_inr_Foreach.scala 134:228:@43871.4]
  wire  _T_1915; // @[sm_x579_inr_Foreach.scala 134:236:@43872.4]
  wire  _T_1952; // @[package.scala 96:25:@43943.4 package.scala 96:25:@43944.4]
  wire  _T_1954; // @[implicits.scala 56:10:@43945.4]
  wire  _T_1955; // @[sm_x579_inr_Foreach.scala 153:115:@43946.4]
  wire  _T_1957; // @[sm_x579_inr_Foreach.scala 153:212:@43948.4]
  wire  x774_b562_D5; // @[package.scala 96:25:@43909.4 package.scala 96:25:@43910.4]
  wire  _T_1959; // @[sm_x579_inr_Foreach.scala 153:257:@43950.4]
  wire  x775_b552_D5; // @[package.scala 96:25:@43919.4 package.scala 96:25:@43920.4]
  wire  _T_1960; // @[sm_x579_inr_Foreach.scala 153:265:@43951.4]
  wire  x776_b543_D5; // @[package.scala 96:25:@43929.4 package.scala 96:25:@43930.4]
  wire  _T_1972; // @[package.scala 96:25:@43969.4 package.scala 96:25:@43970.4]
  wire  _T_1974; // @[implicits.scala 56:10:@43971.4]
  wire  _T_1975; // @[sm_x579_inr_Foreach.scala 158:115:@43972.4]
  wire  _T_1977; // @[sm_x579_inr_Foreach.scala 158:212:@43974.4]
  wire  _T_1979; // @[sm_x579_inr_Foreach.scala 158:257:@43976.4]
  wire  _T_1980; // @[sm_x579_inr_Foreach.scala 158:265:@43977.4]
  wire  _T_1992; // @[package.scala 96:25:@43995.4 package.scala 96:25:@43996.4]
  wire  _T_1994; // @[implicits.scala 56:10:@43997.4]
  wire  _T_1995; // @[sm_x579_inr_Foreach.scala 163:115:@43998.4]
  wire  _T_1997; // @[sm_x579_inr_Foreach.scala 163:212:@44000.4]
  wire  _T_1999; // @[sm_x579_inr_Foreach.scala 163:257:@44002.4]
  wire  _T_2000; // @[sm_x579_inr_Foreach.scala 163:265:@44003.4]
  wire  _T_2012; // @[package.scala 96:25:@44021.4 package.scala 96:25:@44022.4]
  wire  _T_2014; // @[implicits.scala 56:10:@44023.4]
  wire  _T_2015; // @[sm_x579_inr_Foreach.scala 168:115:@44024.4]
  wire  _T_2017; // @[sm_x579_inr_Foreach.scala 168:212:@44026.4]
  wire  _T_2019; // @[sm_x579_inr_Foreach.scala 168:257:@44028.4]
  wire  _T_2020; // @[sm_x579_inr_Foreach.scala 168:265:@44029.4]
  wire  _T_2032; // @[package.scala 96:25:@44047.4 package.scala 96:25:@44048.4]
  wire  _T_2034; // @[implicits.scala 56:10:@44049.4]
  wire  _T_2035; // @[sm_x579_inr_Foreach.scala 173:115:@44050.4]
  wire  _T_2037; // @[sm_x579_inr_Foreach.scala 173:212:@44052.4]
  wire  _T_2039; // @[sm_x579_inr_Foreach.scala 173:257:@44054.4]
  wire  _T_2040; // @[sm_x579_inr_Foreach.scala 173:265:@44055.4]
  wire  _T_2045; // @[package.scala 96:25:@44068.4 package.scala 96:25:@44069.4]
  wire  _T_2051; // @[package.scala 96:25:@44079.4 package.scala 96:25:@44080.4]
  wire  _T_2057; // @[package.scala 96:25:@44090.4 package.scala 96:25:@44091.4]
  wire  _T_2063; // @[package.scala 96:25:@44101.4 package.scala 96:25:@44102.4]
  wire  _T_2069; // @[package.scala 96:25:@44112.4 package.scala 96:25:@44113.4]
  wire [31:0] x565_sum_number; // @[Math.scala 154:22:@43752.4 Math.scala 155:14:@43753.4]
  wire [31:0] x570_sum_number; // @[Math.scala 154:22:@43843.4 Math.scala 155:14:@43844.4]
  wire [31:0] x773_b561_D5_number; // @[package.scala 96:25:@43899.4 package.scala 96:25:@43900.4]
  _ _ ( // @[Math.scala 720:24:@43711.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x739_sum x745_sum_1 ( // @[Math.scala 150:24:@43726.4]
    .clock(x745_sum_1_clock),
    .reset(x745_sum_1_reset),
    .io_a(x745_sum_1_io_a),
    .io_b(x745_sum_1_io_b),
    .io_flow(x745_sum_1_io_flow),
    .io_result(x745_sum_1_io_result)
  );
  RetimeWrapper_31 RetimeWrapper ( // @[package.scala 93:22:@43737.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x739_sum x565_sum_1 ( // @[Math.scala 150:24:@43746.4]
    .clock(x565_sum_1_clock),
    .reset(x565_sum_1_reset),
    .io_a(x565_sum_1_io_a),
    .io_b(x565_sum_1_io_b),
    .io_flow(x565_sum_1_io_flow),
    .io_result(x565_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@43757.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@43767.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@43777.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@43789.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@43801.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  x739_sum x747_sum_1 ( // @[Math.scala 150:24:@43827.4]
    .clock(x747_sum_1_clock),
    .reset(x747_sum_1_reset),
    .io_a(x747_sum_1_io_a),
    .io_b(x747_sum_1_io_b),
    .io_flow(x747_sum_1_io_flow),
    .io_result(x747_sum_1_io_result)
  );
  x739_sum x570_sum_1 ( // @[Math.scala 150:24:@43837.4]
    .clock(x570_sum_1_clock),
    .reset(x570_sum_1_reset),
    .io_a(x570_sum_1_io_a),
    .io_b(x570_sum_1_io_b),
    .io_flow(x570_sum_1_io_flow),
    .io_result(x570_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@43850.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@43862.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  x573_sub x573_sub_1 ( // @[Math.scala 191:24:@43883.4]
    .clock(x573_sub_1_clock),
    .reset(x573_sub_1_reset),
    .io_a(x573_sub_1_io_a),
    .io_b(x573_sub_1_io_b),
    .io_result(x573_sub_1_io_result)
  );
  RetimeWrapper_474 RetimeWrapper_8 ( // @[package.scala 93:22:@43894.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_9 ( // @[package.scala 93:22:@43904.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_10 ( // @[package.scala 93:22:@43914.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_11 ( // @[package.scala 93:22:@43924.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_12 ( // @[package.scala 93:22:@43938.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_13 ( // @[package.scala 93:22:@43964.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_14 ( // @[package.scala 93:22:@43990.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_15 ( // @[package.scala 93:22:@44016.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_16 ( // @[package.scala 93:22:@44042.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper RetimeWrapper_17 ( // @[package.scala 93:22:@44063.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 ( // @[package.scala 93:22:@44074.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper RetimeWrapper_19 ( // @[package.scala 93:22:@44085.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper RetimeWrapper_20 ( // @[package.scala 93:22:@44096.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper RetimeWrapper_21 ( // @[package.scala 93:22:@44107.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  assign _GEN_0 = {{1'd0}, io_in_b542_number}; // @[Math.scala 461:32:@43722.4]
  assign _T_1817 = _GEN_0 << 1; // @[Math.scala 461:32:@43722.4]
  assign _T_1859 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@43794.4 package.scala 96:25:@43795.4]
  assign _T_1861 = io_rr ? _T_1859 : 1'h0; // @[implicits.scala 56:10:@43796.4]
  assign _T_1862 = ~ io_sigsIn_break; // @[sm_x579_inr_Foreach.scala 119:114:@43797.4]
  assign _T_1863 = _T_1861 & _T_1862; // @[sm_x579_inr_Foreach.scala 119:111:@43798.4]
  assign _T_1868 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@43806.4 package.scala 96:25:@43807.4]
  assign _T_1870 = io_rr ? _T_1868 : 1'h0; // @[implicits.scala 56:10:@43808.4]
  assign _T_1871 = _T_1863 & _T_1870; // @[sm_x579_inr_Foreach.scala 119:131:@43809.4]
  assign x772_b562_D2 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@43782.4 package.scala 96:25:@43783.4]
  assign _T_1872 = _T_1871 & x772_b562_D2; // @[sm_x579_inr_Foreach.scala 119:228:@43810.4]
  assign x771_b552_D2 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@43772.4 package.scala 96:25:@43773.4]
  assign _T_1873 = _T_1872 & x771_b552_D2; // @[sm_x579_inr_Foreach.scala 119:236:@43811.4]
  assign x770_b543_D2 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@43762.4 package.scala 96:25:@43763.4]
  assign _GEN_1 = {{1'd0}, io_in_b550_number}; // @[Math.scala 461:32:@43823.4]
  assign _T_1879 = _GEN_1 << 1; // @[Math.scala 461:32:@43823.4]
  assign _T_1901 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@43855.4 package.scala 96:25:@43856.4]
  assign _T_1903 = io_rr ? _T_1901 : 1'h0; // @[implicits.scala 56:10:@43857.4]
  assign _T_1905 = _T_1903 & _T_1862; // @[sm_x579_inr_Foreach.scala 134:111:@43859.4]
  assign _T_1910 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@43867.4 package.scala 96:25:@43868.4]
  assign _T_1912 = io_rr ? _T_1910 : 1'h0; // @[implicits.scala 56:10:@43869.4]
  assign _T_1913 = _T_1905 & _T_1912; // @[sm_x579_inr_Foreach.scala 134:131:@43870.4]
  assign _T_1914 = _T_1913 & x772_b562_D2; // @[sm_x579_inr_Foreach.scala 134:228:@43871.4]
  assign _T_1915 = _T_1914 & x771_b552_D2; // @[sm_x579_inr_Foreach.scala 134:236:@43872.4]
  assign _T_1952 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@43943.4 package.scala 96:25:@43944.4]
  assign _T_1954 = io_rr ? _T_1952 : 1'h0; // @[implicits.scala 56:10:@43945.4]
  assign _T_1955 = _T_1862 & _T_1954; // @[sm_x579_inr_Foreach.scala 153:115:@43946.4]
  assign _T_1957 = _T_1955 & _T_1862; // @[sm_x579_inr_Foreach.scala 153:212:@43948.4]
  assign x774_b562_D5 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@43909.4 package.scala 96:25:@43910.4]
  assign _T_1959 = _T_1957 & x774_b562_D5; // @[sm_x579_inr_Foreach.scala 153:257:@43950.4]
  assign x775_b552_D5 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@43919.4 package.scala 96:25:@43920.4]
  assign _T_1960 = _T_1959 & x775_b552_D5; // @[sm_x579_inr_Foreach.scala 153:265:@43951.4]
  assign x776_b543_D5 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@43929.4 package.scala 96:25:@43930.4]
  assign _T_1972 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@43969.4 package.scala 96:25:@43970.4]
  assign _T_1974 = io_rr ? _T_1972 : 1'h0; // @[implicits.scala 56:10:@43971.4]
  assign _T_1975 = _T_1862 & _T_1974; // @[sm_x579_inr_Foreach.scala 158:115:@43972.4]
  assign _T_1977 = _T_1975 & _T_1862; // @[sm_x579_inr_Foreach.scala 158:212:@43974.4]
  assign _T_1979 = _T_1977 & x774_b562_D5; // @[sm_x579_inr_Foreach.scala 158:257:@43976.4]
  assign _T_1980 = _T_1979 & x775_b552_D5; // @[sm_x579_inr_Foreach.scala 158:265:@43977.4]
  assign _T_1992 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@43995.4 package.scala 96:25:@43996.4]
  assign _T_1994 = io_rr ? _T_1992 : 1'h0; // @[implicits.scala 56:10:@43997.4]
  assign _T_1995 = _T_1862 & _T_1994; // @[sm_x579_inr_Foreach.scala 163:115:@43998.4]
  assign _T_1997 = _T_1995 & _T_1862; // @[sm_x579_inr_Foreach.scala 163:212:@44000.4]
  assign _T_1999 = _T_1997 & x774_b562_D5; // @[sm_x579_inr_Foreach.scala 163:257:@44002.4]
  assign _T_2000 = _T_1999 & x775_b552_D5; // @[sm_x579_inr_Foreach.scala 163:265:@44003.4]
  assign _T_2012 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@44021.4 package.scala 96:25:@44022.4]
  assign _T_2014 = io_rr ? _T_2012 : 1'h0; // @[implicits.scala 56:10:@44023.4]
  assign _T_2015 = _T_1862 & _T_2014; // @[sm_x579_inr_Foreach.scala 168:115:@44024.4]
  assign _T_2017 = _T_2015 & _T_1862; // @[sm_x579_inr_Foreach.scala 168:212:@44026.4]
  assign _T_2019 = _T_2017 & x774_b562_D5; // @[sm_x579_inr_Foreach.scala 168:257:@44028.4]
  assign _T_2020 = _T_2019 & x775_b552_D5; // @[sm_x579_inr_Foreach.scala 168:265:@44029.4]
  assign _T_2032 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@44047.4 package.scala 96:25:@44048.4]
  assign _T_2034 = io_rr ? _T_2032 : 1'h0; // @[implicits.scala 56:10:@44049.4]
  assign _T_2035 = _T_1862 & _T_2034; // @[sm_x579_inr_Foreach.scala 173:115:@44050.4]
  assign _T_2037 = _T_2035 & _T_1862; // @[sm_x579_inr_Foreach.scala 173:212:@44052.4]
  assign _T_2039 = _T_2037 & x774_b562_D5; // @[sm_x579_inr_Foreach.scala 173:257:@44054.4]
  assign _T_2040 = _T_2039 & x775_b552_D5; // @[sm_x579_inr_Foreach.scala 173:265:@44055.4]
  assign _T_2045 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@44068.4 package.scala 96:25:@44069.4]
  assign _T_2051 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@44079.4 package.scala 96:25:@44080.4]
  assign _T_2057 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@44090.4 package.scala 96:25:@44091.4]
  assign _T_2063 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@44101.4 package.scala 96:25:@44102.4]
  assign _T_2069 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@44112.4 package.scala 96:25:@44113.4]
  assign x565_sum_number = x565_sum_1_io_result; // @[Math.scala 154:22:@43752.4 Math.scala 155:14:@43753.4]
  assign x570_sum_number = x570_sum_1_io_result; // @[Math.scala 154:22:@43843.4 Math.scala 155:14:@43844.4]
  assign x773_b561_D5_number = RetimeWrapper_8_io_out; // @[package.scala 96:25:@43899.4 package.scala 96:25:@43900.4]
  assign io_in_x555_tmp_1_wPort_0_ofs_0 = x773_b561_D5_number[1:0]; // @[MemInterfaceType.scala 89:54:@43954.4]
  assign io_in_x555_tmp_1_wPort_0_data_0 = x573_sub_1_io_result; // @[MemInterfaceType.scala 90:56:@43955.4]
  assign io_in_x555_tmp_1_wPort_0_en_0 = _T_1960 & x776_b543_D5; // @[MemInterfaceType.scala 93:57:@43957.4]
  assign io_in_x555_tmp_1_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@44082.4]
  assign io_in_x555_tmp_1_sDone_0 = io_rr ? _T_2051 : 1'h0; // @[MemInterfaceType.scala 197:17:@44083.4]
  assign io_in_x472_A_sram_1_rPort_0_ofs_0 = x570_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@43876.4]
  assign io_in_x472_A_sram_1_rPort_0_en_0 = _T_1915 & x770_b543_D2; // @[MemInterfaceType.scala 110:79:@43878.4]
  assign io_in_x471_A_sram_0_rPort_0_ofs_0 = x565_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@43815.4]
  assign io_in_x471_A_sram_0_rPort_0_en_0 = _T_1873 & x770_b543_D2; // @[MemInterfaceType.scala 110:79:@43817.4]
  assign io_in_x554_tmp_0_wPort_0_ofs_0 = x773_b561_D5_number[1:0]; // @[MemInterfaceType.scala 89:54:@43980.4]
  assign io_in_x554_tmp_0_wPort_0_data_0 = x573_sub_1_io_result; // @[MemInterfaceType.scala 90:56:@43981.4]
  assign io_in_x554_tmp_0_wPort_0_en_0 = _T_1980 & x776_b543_D5; // @[MemInterfaceType.scala 93:57:@43983.4]
  assign io_in_x554_tmp_0_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@44071.4]
  assign io_in_x554_tmp_0_sDone_0 = io_rr ? _T_2045 : 1'h0; // @[MemInterfaceType.scala 197:17:@44072.4]
  assign io_in_x558_tmp_4_wPort_0_ofs_0 = x773_b561_D5_number[1:0]; // @[MemInterfaceType.scala 89:54:@44006.4]
  assign io_in_x558_tmp_4_wPort_0_data_0 = x573_sub_1_io_result; // @[MemInterfaceType.scala 90:56:@44007.4]
  assign io_in_x558_tmp_4_wPort_0_en_0 = _T_2000 & x776_b543_D5; // @[MemInterfaceType.scala 93:57:@44009.4]
  assign io_in_x558_tmp_4_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@44115.4]
  assign io_in_x558_tmp_4_sDone_0 = io_rr ? _T_2069 : 1'h0; // @[MemInterfaceType.scala 197:17:@44116.4]
  assign io_in_x557_tmp_3_wPort_0_ofs_0 = x773_b561_D5_number[1:0]; // @[MemInterfaceType.scala 89:54:@44032.4]
  assign io_in_x557_tmp_3_wPort_0_data_0 = x573_sub_1_io_result; // @[MemInterfaceType.scala 90:56:@44033.4]
  assign io_in_x557_tmp_3_wPort_0_en_0 = _T_2020 & x776_b543_D5; // @[MemInterfaceType.scala 93:57:@44035.4]
  assign io_in_x557_tmp_3_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@44104.4]
  assign io_in_x557_tmp_3_sDone_0 = io_rr ? _T_2063 : 1'h0; // @[MemInterfaceType.scala 197:17:@44105.4]
  assign io_in_x556_tmp_2_wPort_0_ofs_0 = x773_b561_D5_number[1:0]; // @[MemInterfaceType.scala 89:54:@44058.4]
  assign io_in_x556_tmp_2_wPort_0_data_0 = x573_sub_1_io_result; // @[MemInterfaceType.scala 90:56:@44059.4]
  assign io_in_x556_tmp_2_wPort_0_en_0 = _T_2040 & x776_b543_D5; // @[MemInterfaceType.scala 93:57:@44061.4]
  assign io_in_x556_tmp_2_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@44093.4]
  assign io_in_x556_tmp_2_sDone_0 = io_rr ? _T_2057 : 1'h0; // @[MemInterfaceType.scala 197:17:@44094.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@43714.4]
  assign x745_sum_1_clock = clock; // @[:@43727.4]
  assign x745_sum_1_reset = reset; // @[:@43728.4]
  assign x745_sum_1_io_a = _T_1817[31:0]; // @[Math.scala 151:17:@43729.4]
  assign x745_sum_1_io_b = io_in_b542_number; // @[Math.scala 152:17:@43730.4]
  assign x745_sum_1_io_flow = 1'h1; // @[Math.scala 153:20:@43731.4]
  assign RetimeWrapper_clock = clock; // @[:@43738.4]
  assign RetimeWrapper_reset = reset; // @[:@43739.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@43741.4]
  assign RetimeWrapper_io_in = __io_result; // @[package.scala 94:16:@43740.4]
  assign x565_sum_1_clock = clock; // @[:@43747.4]
  assign x565_sum_1_reset = reset; // @[:@43748.4]
  assign x565_sum_1_io_a = x745_sum_1_io_result; // @[Math.scala 151:17:@43749.4]
  assign x565_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@43750.4]
  assign x565_sum_1_io_flow = 1'h1; // @[Math.scala 153:20:@43751.4]
  assign RetimeWrapper_1_clock = clock; // @[:@43758.4]
  assign RetimeWrapper_1_reset = reset; // @[:@43759.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@43761.4]
  assign RetimeWrapper_1_io_in = io_in_b543; // @[package.scala 94:16:@43760.4]
  assign RetimeWrapper_2_clock = clock; // @[:@43768.4]
  assign RetimeWrapper_2_reset = reset; // @[:@43769.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@43771.4]
  assign RetimeWrapper_2_io_in = io_in_b552; // @[package.scala 94:16:@43770.4]
  assign RetimeWrapper_3_clock = clock; // @[:@43778.4]
  assign RetimeWrapper_3_reset = reset; // @[:@43779.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@43781.4]
  assign RetimeWrapper_3_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@43780.4]
  assign RetimeWrapper_4_clock = clock; // @[:@43790.4]
  assign RetimeWrapper_4_reset = reset; // @[:@43791.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@43793.4]
  assign RetimeWrapper_4_io_in = 1'h1; // @[package.scala 94:16:@43792.4]
  assign RetimeWrapper_5_clock = clock; // @[:@43802.4]
  assign RetimeWrapper_5_reset = reset; // @[:@43803.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@43805.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@43804.4]
  assign x747_sum_1_clock = clock; // @[:@43828.4]
  assign x747_sum_1_reset = reset; // @[:@43829.4]
  assign x747_sum_1_io_a = _T_1879[31:0]; // @[Math.scala 151:17:@43830.4]
  assign x747_sum_1_io_b = io_in_b550_number; // @[Math.scala 152:17:@43831.4]
  assign x747_sum_1_io_flow = 1'h1; // @[Math.scala 153:20:@43832.4]
  assign x570_sum_1_clock = clock; // @[:@43838.4]
  assign x570_sum_1_reset = reset; // @[:@43839.4]
  assign x570_sum_1_io_a = x747_sum_1_io_result; // @[Math.scala 151:17:@43840.4]
  assign x570_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@43841.4]
  assign x570_sum_1_io_flow = 1'h1; // @[Math.scala 153:20:@43842.4]
  assign RetimeWrapper_6_clock = clock; // @[:@43851.4]
  assign RetimeWrapper_6_reset = reset; // @[:@43852.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@43854.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@43853.4]
  assign RetimeWrapper_7_clock = clock; // @[:@43863.4]
  assign RetimeWrapper_7_reset = reset; // @[:@43864.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@43866.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@43865.4]
  assign x573_sub_1_clock = clock; // @[:@43884.4]
  assign x573_sub_1_reset = reset; // @[:@43885.4]
  assign x573_sub_1_io_a = io_in_x471_A_sram_0_rPort_0_output_0; // @[Math.scala 192:17:@43886.4]
  assign x573_sub_1_io_b = io_in_x472_A_sram_1_rPort_0_output_0; // @[Math.scala 193:17:@43887.4]
  assign RetimeWrapper_8_clock = clock; // @[:@43895.4]
  assign RetimeWrapper_8_reset = reset; // @[:@43896.4]
  assign RetimeWrapper_8_io_in = __io_result; // @[package.scala 94:16:@43897.4]
  assign RetimeWrapper_9_clock = clock; // @[:@43905.4]
  assign RetimeWrapper_9_reset = reset; // @[:@43906.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@43908.4]
  assign RetimeWrapper_9_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@43907.4]
  assign RetimeWrapper_10_clock = clock; // @[:@43915.4]
  assign RetimeWrapper_10_reset = reset; // @[:@43916.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@43918.4]
  assign RetimeWrapper_10_io_in = io_in_b552; // @[package.scala 94:16:@43917.4]
  assign RetimeWrapper_11_clock = clock; // @[:@43925.4]
  assign RetimeWrapper_11_reset = reset; // @[:@43926.4]
  assign RetimeWrapper_11_io_flow = 1'h1; // @[package.scala 95:18:@43928.4]
  assign RetimeWrapper_11_io_in = io_in_b543; // @[package.scala 94:16:@43927.4]
  assign RetimeWrapper_12_clock = clock; // @[:@43939.4]
  assign RetimeWrapper_12_reset = reset; // @[:@43940.4]
  assign RetimeWrapper_12_io_flow = 1'h1; // @[package.scala 95:18:@43942.4]
  assign RetimeWrapper_12_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@43941.4]
  assign RetimeWrapper_13_clock = clock; // @[:@43965.4]
  assign RetimeWrapper_13_reset = reset; // @[:@43966.4]
  assign RetimeWrapper_13_io_flow = 1'h1; // @[package.scala 95:18:@43968.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@43967.4]
  assign RetimeWrapper_14_clock = clock; // @[:@43991.4]
  assign RetimeWrapper_14_reset = reset; // @[:@43992.4]
  assign RetimeWrapper_14_io_flow = 1'h1; // @[package.scala 95:18:@43994.4]
  assign RetimeWrapper_14_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@43993.4]
  assign RetimeWrapper_15_clock = clock; // @[:@44017.4]
  assign RetimeWrapper_15_reset = reset; // @[:@44018.4]
  assign RetimeWrapper_15_io_flow = 1'h1; // @[package.scala 95:18:@44020.4]
  assign RetimeWrapper_15_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44019.4]
  assign RetimeWrapper_16_clock = clock; // @[:@44043.4]
  assign RetimeWrapper_16_reset = reset; // @[:@44044.4]
  assign RetimeWrapper_16_io_flow = 1'h1; // @[package.scala 95:18:@44046.4]
  assign RetimeWrapper_16_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@44045.4]
  assign RetimeWrapper_17_clock = clock; // @[:@44064.4]
  assign RetimeWrapper_17_reset = reset; // @[:@44065.4]
  assign RetimeWrapper_17_io_flow = 1'h1; // @[package.scala 95:18:@44067.4]
  assign RetimeWrapper_17_io_in = io_sigsIn_done; // @[package.scala 94:16:@44066.4]
  assign RetimeWrapper_18_clock = clock; // @[:@44075.4]
  assign RetimeWrapper_18_reset = reset; // @[:@44076.4]
  assign RetimeWrapper_18_io_flow = 1'h1; // @[package.scala 95:18:@44078.4]
  assign RetimeWrapper_18_io_in = io_sigsIn_done; // @[package.scala 94:16:@44077.4]
  assign RetimeWrapper_19_clock = clock; // @[:@44086.4]
  assign RetimeWrapper_19_reset = reset; // @[:@44087.4]
  assign RetimeWrapper_19_io_flow = 1'h1; // @[package.scala 95:18:@44089.4]
  assign RetimeWrapper_19_io_in = io_sigsIn_done; // @[package.scala 94:16:@44088.4]
  assign RetimeWrapper_20_clock = clock; // @[:@44097.4]
  assign RetimeWrapper_20_reset = reset; // @[:@44098.4]
  assign RetimeWrapper_20_io_flow = 1'h1; // @[package.scala 95:18:@44100.4]
  assign RetimeWrapper_20_io_in = io_sigsIn_done; // @[package.scala 94:16:@44099.4]
  assign RetimeWrapper_21_clock = clock; // @[:@44108.4]
  assign RetimeWrapper_21_reset = reset; // @[:@44109.4]
  assign RetimeWrapper_21_io_flow = 1'h1; // @[package.scala 95:18:@44111.4]
  assign RetimeWrapper_21_io_in = io_sigsIn_done; // @[package.scala 94:16:@44110.4]
endmodule
module RetimeWrapper_500( // @[:@44592.2]
  input         clock, // @[:@44593.4]
  input         reset, // @[:@44594.4]
  input         io_flow, // @[:@44595.4]
  input  [31:0] io_in, // @[:@44595.4]
  output [31:0] io_out // @[:@44595.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@44597.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@44597.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@44597.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@44597.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@44597.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@44597.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@44597.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@44610.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@44609.4]
  assign sr_init = 32'h2; // @[RetimeShiftRegister.scala 19:16:@44608.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@44607.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@44606.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@44604.4]
endmodule
module NBufCtr_66( // @[:@44612.2]
  input         clock, // @[:@44613.4]
  input         reset, // @[:@44614.4]
  input         io_input_enable, // @[:@44615.4]
  output [31:0] io_output_count // @[:@44615.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@44652.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@44652.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@44652.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@44652.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@44652.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@44657.4 package.scala 96:25:@44658.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@44618.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@44619.4]
  wire  _T_21; // @[Counter.scala 49:55:@44620.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@44621.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@44622.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@44623.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@44624.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@44625.4]
  wire  _T_33; // @[Counter.scala 51:52:@44629.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@44630.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@44631.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@44632.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@44633.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@44634.4]
  RetimeWrapper_500 RetimeWrapper ( // @[package.scala 93:22:@44652.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@44657.4 package.scala 96:25:@44658.4]
  assign _T_18 = {{1'd0}, _T_66}; // @[Counter.scala 49:32:@44618.4]
  assign _T_19 = _T_18[31:0]; // @[Counter.scala 49:32:@44619.4]
  assign _T_21 = _T_19 >= 32'h3; // @[Counter.scala 49:55:@44620.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@44621.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh3); // @[Counter.scala 49:91:@44622.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh3); // @[Counter.scala 49:91:@44623.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@44624.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@44625.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@44629.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@44630.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@44631.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@44632.4]
  assign _T_39 = _T_33 ? 32'h2 : _T_38; // @[Counter.scala 51:47:@44633.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@44634.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@44660.4]
  assign RetimeWrapper_clock = clock; // @[:@44653.4]
  assign RetimeWrapper_reset = reset; // @[:@44654.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@44656.4]
  assign RetimeWrapper_io_in = reset ? 32'h2 : _T_40; // @[package.scala 94:16:@44655.4]
endmodule
module NBufCtr_68( // @[:@44776.2]
  input         clock, // @[:@44777.4]
  input         reset, // @[:@44778.4]
  input         io_input_enable, // @[:@44779.4]
  output [31:0] io_output_count // @[:@44779.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@44816.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@44816.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@44816.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@44816.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@44816.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@44821.4 package.scala 96:25:@44822.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@44782.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@44783.4]
  wire  _T_21; // @[Counter.scala 49:55:@44784.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@44785.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@44786.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@44787.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@44788.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@44789.4]
  wire  _T_33; // @[Counter.scala 51:52:@44793.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@44794.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@44795.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@44796.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@44797.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@44798.4]
  RetimeWrapper_500 RetimeWrapper ( // @[package.scala 93:22:@44816.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@44821.4 package.scala 96:25:@44822.4]
  assign _T_18 = _T_66 + 32'h1; // @[Counter.scala 49:32:@44782.4]
  assign _T_19 = _T_66 + 32'h1; // @[Counter.scala 49:32:@44783.4]
  assign _T_21 = _T_19 >= 32'h3; // @[Counter.scala 49:55:@44784.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@44785.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh2); // @[Counter.scala 49:91:@44786.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh2); // @[Counter.scala 49:91:@44787.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@44788.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@44789.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@44793.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@44794.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@44795.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@44796.4]
  assign _T_39 = _T_33 ? 32'h2 : _T_38; // @[Counter.scala 51:47:@44797.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@44798.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@44824.4]
  assign RetimeWrapper_clock = clock; // @[:@44817.4]
  assign RetimeWrapper_reset = reset; // @[:@44818.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@44820.4]
  assign RetimeWrapper_io_in = reset ? 32'h2 : _T_40; // @[package.scala 94:16:@44819.4]
endmodule
module NBufCtr_69( // @[:@44858.2]
  input         clock, // @[:@44859.4]
  input         reset, // @[:@44860.4]
  input         io_input_enable, // @[:@44861.4]
  output [31:0] io_output_count // @[:@44861.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@44898.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@44898.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@44898.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@44898.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@44898.4]
  wire [31:0] _T_66; // @[package.scala 96:25:@44903.4 package.scala 96:25:@44904.4]
  wire [32:0] _T_18; // @[Counter.scala 49:32:@44864.4]
  wire [31:0] _T_19; // @[Counter.scala 49:32:@44865.4]
  wire  _T_21; // @[Counter.scala 49:55:@44866.4]
  wire [31:0] _T_22; // @[Counter.scala 49:84:@44867.4]
  wire [32:0] _T_24; // @[Counter.scala 49:91:@44868.4]
  wire [31:0] _T_25; // @[Counter.scala 49:91:@44869.4]
  wire [31:0] _T_26; // @[Counter.scala 49:91:@44870.4]
  wire [31:0] _T_27; // @[Counter.scala 49:126:@44871.4]
  wire  _T_33; // @[Counter.scala 51:52:@44875.4]
  wire [32:0] _T_36; // @[Counter.scala 51:103:@44876.4]
  wire [32:0] _T_37; // @[Counter.scala 51:103:@44877.4]
  wire [31:0] _T_38; // @[Counter.scala 51:103:@44878.4]
  wire [31:0] _T_39; // @[Counter.scala 51:47:@44879.4]
  wire [31:0] _T_40; // @[Counter.scala 51:26:@44880.4]
  RetimeWrapper_500 RetimeWrapper ( // @[package.scala 93:22:@44898.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_66 = RetimeWrapper_io_out; // @[package.scala 96:25:@44903.4 package.scala 96:25:@44904.4]
  assign _T_18 = _T_66 + 32'h2; // @[Counter.scala 49:32:@44864.4]
  assign _T_19 = _T_66 + 32'h2; // @[Counter.scala 49:32:@44865.4]
  assign _T_21 = _T_19 >= 32'h3; // @[Counter.scala 49:55:@44866.4]
  assign _T_22 = $signed(_T_66); // @[Counter.scala 49:84:@44867.4]
  assign _T_24 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 49:91:@44868.4]
  assign _T_25 = $signed(_T_22) + $signed(-32'sh1); // @[Counter.scala 49:91:@44869.4]
  assign _T_26 = $signed(_T_25); // @[Counter.scala 49:91:@44870.4]
  assign _T_27 = $unsigned(_T_26); // @[Counter.scala 49:126:@44871.4]
  assign _T_33 = _T_66 == 32'h0; // @[Counter.scala 51:52:@44875.4]
  assign _T_36 = _T_66 - 32'h1; // @[Counter.scala 51:103:@44876.4]
  assign _T_37 = $unsigned(_T_36); // @[Counter.scala 51:103:@44877.4]
  assign _T_38 = _T_37[31:0]; // @[Counter.scala 51:103:@44878.4]
  assign _T_39 = _T_33 ? 32'h2 : _T_38; // @[Counter.scala 51:47:@44879.4]
  assign _T_40 = io_input_enable ? _T_39 : _T_66; // @[Counter.scala 51:26:@44880.4]
  assign io_output_count = _T_21 ? _T_27 : _T_19; // @[Counter.scala 55:21:@44906.4]
  assign RetimeWrapper_clock = clock; // @[:@44899.4]
  assign RetimeWrapper_reset = reset; // @[:@44900.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@44902.4]
  assign RetimeWrapper_io_in = reset ? 32'h2 : _T_40; // @[package.scala 94:16:@44901.4]
endmodule
module NBufController_10( // @[:@44908.2]
  input        clock, // @[:@44909.4]
  input        reset, // @[:@44910.4]
  input        io_sEn_0, // @[:@44911.4]
  input        io_sEn_1, // @[:@44911.4]
  input        io_sEn_2, // @[:@44911.4]
  input        io_sDone_0, // @[:@44911.4]
  input        io_sDone_1, // @[:@44911.4]
  input        io_sDone_2, // @[:@44911.4]
  output [2:0] io_statesInW_0, // @[:@44911.4]
  output [2:0] io_statesInR_1, // @[:@44911.4]
  output [2:0] io_statesInR_2 // @[:@44911.4]
);
  wire  sEn_latch_0_clock; // @[NBuffers.scala 21:52:@44913.4]
  wire  sEn_latch_0_reset; // @[NBuffers.scala 21:52:@44913.4]
  wire  sEn_latch_0_io_input_set; // @[NBuffers.scala 21:52:@44913.4]
  wire  sEn_latch_0_io_input_reset; // @[NBuffers.scala 21:52:@44913.4]
  wire  sEn_latch_0_io_input_asyn_reset; // @[NBuffers.scala 21:52:@44913.4]
  wire  sEn_latch_0_io_output; // @[NBuffers.scala 21:52:@44913.4]
  wire  sEn_latch_1_clock; // @[NBuffers.scala 21:52:@44916.4]
  wire  sEn_latch_1_reset; // @[NBuffers.scala 21:52:@44916.4]
  wire  sEn_latch_1_io_input_set; // @[NBuffers.scala 21:52:@44916.4]
  wire  sEn_latch_1_io_input_reset; // @[NBuffers.scala 21:52:@44916.4]
  wire  sEn_latch_1_io_input_asyn_reset; // @[NBuffers.scala 21:52:@44916.4]
  wire  sEn_latch_1_io_output; // @[NBuffers.scala 21:52:@44916.4]
  wire  sEn_latch_2_clock; // @[NBuffers.scala 21:52:@44919.4]
  wire  sEn_latch_2_reset; // @[NBuffers.scala 21:52:@44919.4]
  wire  sEn_latch_2_io_input_set; // @[NBuffers.scala 21:52:@44919.4]
  wire  sEn_latch_2_io_input_reset; // @[NBuffers.scala 21:52:@44919.4]
  wire  sEn_latch_2_io_input_asyn_reset; // @[NBuffers.scala 21:52:@44919.4]
  wire  sEn_latch_2_io_output; // @[NBuffers.scala 21:52:@44919.4]
  wire  sDone_latch_0_clock; // @[NBuffers.scala 22:54:@44922.4]
  wire  sDone_latch_0_reset; // @[NBuffers.scala 22:54:@44922.4]
  wire  sDone_latch_0_io_input_set; // @[NBuffers.scala 22:54:@44922.4]
  wire  sDone_latch_0_io_input_reset; // @[NBuffers.scala 22:54:@44922.4]
  wire  sDone_latch_0_io_input_asyn_reset; // @[NBuffers.scala 22:54:@44922.4]
  wire  sDone_latch_0_io_output; // @[NBuffers.scala 22:54:@44922.4]
  wire  sDone_latch_1_clock; // @[NBuffers.scala 22:54:@44925.4]
  wire  sDone_latch_1_reset; // @[NBuffers.scala 22:54:@44925.4]
  wire  sDone_latch_1_io_input_set; // @[NBuffers.scala 22:54:@44925.4]
  wire  sDone_latch_1_io_input_reset; // @[NBuffers.scala 22:54:@44925.4]
  wire  sDone_latch_1_io_input_asyn_reset; // @[NBuffers.scala 22:54:@44925.4]
  wire  sDone_latch_1_io_output; // @[NBuffers.scala 22:54:@44925.4]
  wire  sDone_latch_2_clock; // @[NBuffers.scala 22:54:@44928.4]
  wire  sDone_latch_2_reset; // @[NBuffers.scala 22:54:@44928.4]
  wire  sDone_latch_2_io_input_set; // @[NBuffers.scala 22:54:@44928.4]
  wire  sDone_latch_2_io_input_reset; // @[NBuffers.scala 22:54:@44928.4]
  wire  sDone_latch_2_io_input_asyn_reset; // @[NBuffers.scala 22:54:@44928.4]
  wire  sDone_latch_2_io_output; // @[NBuffers.scala 22:54:@44928.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@44935.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@44935.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@44935.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@44935.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@44935.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@44943.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@44943.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@44943.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@44943.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@44943.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@44952.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@44952.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@44952.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@44952.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@44952.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@44960.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@44960.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@44960.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@44960.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@44960.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@44971.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@44971.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@44971.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@44971.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@44971.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@44979.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@44979.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@44979.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@44979.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@44979.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@44988.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@44988.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@44988.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@44988.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@44988.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@44996.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@44996.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@44996.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@44996.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@44996.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@45007.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@45007.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@45007.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@45007.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@45007.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@45015.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@45015.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@45015.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@45015.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@45015.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@45024.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@45024.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@45024.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@45024.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@45024.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@45032.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@45032.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@45032.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@45032.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@45032.4]
  wire  NBufCtr_clock; // @[NBuffers.scala 40:19:@45057.4]
  wire  NBufCtr_reset; // @[NBuffers.scala 40:19:@45057.4]
  wire  NBufCtr_io_input_enable; // @[NBuffers.scala 40:19:@45057.4]
  wire [31:0] NBufCtr_io_output_count; // @[NBuffers.scala 40:19:@45057.4]
  wire  statesInR_0_clock; // @[NBuffers.scala 50:19:@45068.4]
  wire  statesInR_0_reset; // @[NBuffers.scala 50:19:@45068.4]
  wire  statesInR_0_io_input_enable; // @[NBuffers.scala 50:19:@45068.4]
  wire [31:0] statesInR_0_io_output_count; // @[NBuffers.scala 50:19:@45068.4]
  wire  statesInR_1_clock; // @[NBuffers.scala 50:19:@45079.4]
  wire  statesInR_1_reset; // @[NBuffers.scala 50:19:@45079.4]
  wire  statesInR_1_io_input_enable; // @[NBuffers.scala 50:19:@45079.4]
  wire [31:0] statesInR_1_io_output_count; // @[NBuffers.scala 50:19:@45079.4]
  wire  statesInR_2_clock; // @[NBuffers.scala 50:19:@45090.4]
  wire  statesInR_2_reset; // @[NBuffers.scala 50:19:@45090.4]
  wire  statesInR_2_io_input_enable; // @[NBuffers.scala 50:19:@45090.4]
  wire [31:0] statesInR_2_io_output_count; // @[NBuffers.scala 50:19:@45090.4]
  wire  _T_33; // @[NBuffers.scala 26:46:@44932.4]
  wire  _T_48; // @[NBuffers.scala 26:46:@44968.4]
  wire  _T_63; // @[NBuffers.scala 26:46:@45004.4]
  wire  _T_77; // @[NBuffers.scala 33:64:@45040.4]
  wire  anyEnabled; // @[NBuffers.scala 33:64:@45041.4]
  wire  _T_78; // @[NBuffers.scala 34:124:@45042.4]
  wire  _T_79; // @[NBuffers.scala 34:104:@45043.4]
  wire  _T_80; // @[NBuffers.scala 34:124:@45044.4]
  wire  _T_81; // @[NBuffers.scala 34:104:@45045.4]
  wire  _T_82; // @[NBuffers.scala 34:124:@45046.4]
  wire  _T_83; // @[NBuffers.scala 34:104:@45047.4]
  wire  _T_84; // @[NBuffers.scala 34:150:@45048.4]
  wire  _T_85; // @[NBuffers.scala 34:150:@45049.4]
  wire  _T_86; // @[NBuffers.scala 34:154:@45050.4]
  wire  _T_88; // @[package.scala 100:49:@45051.4]
  reg  _T_91; // @[package.scala 48:56:@45052.4]
  reg [31:0] _RAND_0;
  SRFF sEn_latch_0 ( // @[NBuffers.scala 21:52:@44913.4]
    .clock(sEn_latch_0_clock),
    .reset(sEn_latch_0_reset),
    .io_input_set(sEn_latch_0_io_input_set),
    .io_input_reset(sEn_latch_0_io_input_reset),
    .io_input_asyn_reset(sEn_latch_0_io_input_asyn_reset),
    .io_output(sEn_latch_0_io_output)
  );
  SRFF sEn_latch_1 ( // @[NBuffers.scala 21:52:@44916.4]
    .clock(sEn_latch_1_clock),
    .reset(sEn_latch_1_reset),
    .io_input_set(sEn_latch_1_io_input_set),
    .io_input_reset(sEn_latch_1_io_input_reset),
    .io_input_asyn_reset(sEn_latch_1_io_input_asyn_reset),
    .io_output(sEn_latch_1_io_output)
  );
  SRFF sEn_latch_2 ( // @[NBuffers.scala 21:52:@44919.4]
    .clock(sEn_latch_2_clock),
    .reset(sEn_latch_2_reset),
    .io_input_set(sEn_latch_2_io_input_set),
    .io_input_reset(sEn_latch_2_io_input_reset),
    .io_input_asyn_reset(sEn_latch_2_io_input_asyn_reset),
    .io_output(sEn_latch_2_io_output)
  );
  SRFF sDone_latch_0 ( // @[NBuffers.scala 22:54:@44922.4]
    .clock(sDone_latch_0_clock),
    .reset(sDone_latch_0_reset),
    .io_input_set(sDone_latch_0_io_input_set),
    .io_input_reset(sDone_latch_0_io_input_reset),
    .io_input_asyn_reset(sDone_latch_0_io_input_asyn_reset),
    .io_output(sDone_latch_0_io_output)
  );
  SRFF sDone_latch_1 ( // @[NBuffers.scala 22:54:@44925.4]
    .clock(sDone_latch_1_clock),
    .reset(sDone_latch_1_reset),
    .io_input_set(sDone_latch_1_io_input_set),
    .io_input_reset(sDone_latch_1_io_input_reset),
    .io_input_asyn_reset(sDone_latch_1_io_input_asyn_reset),
    .io_output(sDone_latch_1_io_output)
  );
  SRFF sDone_latch_2 ( // @[NBuffers.scala 22:54:@44928.4]
    .clock(sDone_latch_2_clock),
    .reset(sDone_latch_2_reset),
    .io_input_set(sDone_latch_2_io_input_set),
    .io_input_reset(sDone_latch_2_io_input_reset),
    .io_input_asyn_reset(sDone_latch_2_io_input_asyn_reset),
    .io_output(sDone_latch_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@44935.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@44943.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@44952.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@44960.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@44971.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@44979.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@44988.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@44996.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@45007.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@45015.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@45024.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 ( // @[package.scala 93:22:@45032.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  NBufCtr_66 NBufCtr ( // @[NBuffers.scala 40:19:@45057.4]
    .clock(NBufCtr_clock),
    .reset(NBufCtr_reset),
    .io_input_enable(NBufCtr_io_input_enable),
    .io_output_count(NBufCtr_io_output_count)
  );
  NBufCtr_66 statesInR_0 ( // @[NBuffers.scala 50:19:@45068.4]
    .clock(statesInR_0_clock),
    .reset(statesInR_0_reset),
    .io_input_enable(statesInR_0_io_input_enable),
    .io_output_count(statesInR_0_io_output_count)
  );
  NBufCtr_68 statesInR_1 ( // @[NBuffers.scala 50:19:@45079.4]
    .clock(statesInR_1_clock),
    .reset(statesInR_1_reset),
    .io_input_enable(statesInR_1_io_input_enable),
    .io_output_count(statesInR_1_io_output_count)
  );
  NBufCtr_69 statesInR_2 ( // @[NBuffers.scala 50:19:@45090.4]
    .clock(statesInR_2_clock),
    .reset(statesInR_2_reset),
    .io_input_enable(statesInR_2_io_input_enable),
    .io_output_count(statesInR_2_io_output_count)
  );
  assign _T_33 = io_sDone_0 == 1'h0; // @[NBuffers.scala 26:46:@44932.4]
  assign _T_48 = io_sDone_1 == 1'h0; // @[NBuffers.scala 26:46:@44968.4]
  assign _T_63 = io_sDone_2 == 1'h0; // @[NBuffers.scala 26:46:@45004.4]
  assign _T_77 = sEn_latch_0_io_output | sEn_latch_1_io_output; // @[NBuffers.scala 33:64:@45040.4]
  assign anyEnabled = _T_77 | sEn_latch_2_io_output; // @[NBuffers.scala 33:64:@45041.4]
  assign _T_78 = sDone_latch_0_io_output | io_sDone_0; // @[NBuffers.scala 34:124:@45042.4]
  assign _T_79 = sEn_latch_0_io_output == _T_78; // @[NBuffers.scala 34:104:@45043.4]
  assign _T_80 = sDone_latch_1_io_output | io_sDone_1; // @[NBuffers.scala 34:124:@45044.4]
  assign _T_81 = sEn_latch_1_io_output == _T_80; // @[NBuffers.scala 34:104:@45045.4]
  assign _T_82 = sDone_latch_2_io_output | io_sDone_2; // @[NBuffers.scala 34:124:@45046.4]
  assign _T_83 = sEn_latch_2_io_output == _T_82; // @[NBuffers.scala 34:104:@45047.4]
  assign _T_84 = _T_79 & _T_81; // @[NBuffers.scala 34:150:@45048.4]
  assign _T_85 = _T_84 & _T_83; // @[NBuffers.scala 34:150:@45049.4]
  assign _T_86 = _T_85 & anyEnabled; // @[NBuffers.scala 34:154:@45050.4]
  assign _T_88 = _T_86 == 1'h0; // @[package.scala 100:49:@45051.4]
  assign io_statesInW_0 = NBufCtr_io_output_count[2:0]; // @[NBuffers.scala 44:21:@45067.4]
  assign io_statesInR_1 = statesInR_1_io_output_count[2:0]; // @[NBuffers.scala 54:21:@45089.4]
  assign io_statesInR_2 = statesInR_2_io_output_count[2:0]; // @[NBuffers.scala 54:21:@45100.4]
  assign sEn_latch_0_clock = clock; // @[:@44914.4]
  assign sEn_latch_0_reset = reset; // @[:@44915.4]
  assign sEn_latch_0_io_input_set = io_sEn_0 & _T_33; // @[NBuffers.scala 26:31:@44934.4]
  assign sEn_latch_0_io_input_reset = RetimeWrapper_io_out; // @[NBuffers.scala 27:33:@44942.4]
  assign sEn_latch_0_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[NBuffers.scala 28:38:@44950.4]
  assign sEn_latch_1_clock = clock; // @[:@44917.4]
  assign sEn_latch_1_reset = reset; // @[:@44918.4]
  assign sEn_latch_1_io_input_set = io_sEn_1 & _T_48; // @[NBuffers.scala 26:31:@44970.4]
  assign sEn_latch_1_io_input_reset = RetimeWrapper_4_io_out; // @[NBuffers.scala 27:33:@44978.4]
  assign sEn_latch_1_io_input_asyn_reset = RetimeWrapper_5_io_out; // @[NBuffers.scala 28:38:@44986.4]
  assign sEn_latch_2_clock = clock; // @[:@44920.4]
  assign sEn_latch_2_reset = reset; // @[:@44921.4]
  assign sEn_latch_2_io_input_set = io_sEn_2 & _T_63; // @[NBuffers.scala 26:31:@45006.4]
  assign sEn_latch_2_io_input_reset = RetimeWrapper_8_io_out; // @[NBuffers.scala 27:33:@45014.4]
  assign sEn_latch_2_io_input_asyn_reset = RetimeWrapper_9_io_out; // @[NBuffers.scala 28:38:@45022.4]
  assign sDone_latch_0_clock = clock; // @[:@44923.4]
  assign sDone_latch_0_reset = reset; // @[:@44924.4]
  assign sDone_latch_0_io_input_set = io_sDone_0; // @[NBuffers.scala 29:33:@44951.4]
  assign sDone_latch_0_io_input_reset = RetimeWrapper_2_io_out; // @[NBuffers.scala 30:35:@44959.4]
  assign sDone_latch_0_io_input_asyn_reset = RetimeWrapper_3_io_out; // @[NBuffers.scala 31:40:@44967.4]
  assign sDone_latch_1_clock = clock; // @[:@44926.4]
  assign sDone_latch_1_reset = reset; // @[:@44927.4]
  assign sDone_latch_1_io_input_set = io_sDone_1; // @[NBuffers.scala 29:33:@44987.4]
  assign sDone_latch_1_io_input_reset = RetimeWrapper_6_io_out; // @[NBuffers.scala 30:35:@44995.4]
  assign sDone_latch_1_io_input_asyn_reset = RetimeWrapper_7_io_out; // @[NBuffers.scala 31:40:@45003.4]
  assign sDone_latch_2_clock = clock; // @[:@44929.4]
  assign sDone_latch_2_reset = reset; // @[:@44930.4]
  assign sDone_latch_2_io_input_set = io_sDone_2; // @[NBuffers.scala 29:33:@45023.4]
  assign sDone_latch_2_io_input_reset = RetimeWrapper_10_io_out; // @[NBuffers.scala 30:35:@45031.4]
  assign sDone_latch_2_io_input_asyn_reset = RetimeWrapper_11_io_out; // @[NBuffers.scala 31:40:@45039.4]
  assign RetimeWrapper_clock = clock; // @[:@44936.4]
  assign RetimeWrapper_reset = reset; // @[:@44937.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@44939.4]
  assign RetimeWrapper_io_in = _T_86 & _T_91; // @[package.scala 94:16:@44938.4]
  assign RetimeWrapper_1_clock = clock; // @[:@44944.4]
  assign RetimeWrapper_1_reset = reset; // @[:@44945.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@44947.4]
  assign RetimeWrapper_1_io_in = reset; // @[package.scala 94:16:@44946.4]
  assign RetimeWrapper_2_clock = clock; // @[:@44953.4]
  assign RetimeWrapper_2_reset = reset; // @[:@44954.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@44956.4]
  assign RetimeWrapper_2_io_in = _T_86 & _T_91; // @[package.scala 94:16:@44955.4]
  assign RetimeWrapper_3_clock = clock; // @[:@44961.4]
  assign RetimeWrapper_3_reset = reset; // @[:@44962.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@44964.4]
  assign RetimeWrapper_3_io_in = reset; // @[package.scala 94:16:@44963.4]
  assign RetimeWrapper_4_clock = clock; // @[:@44972.4]
  assign RetimeWrapper_4_reset = reset; // @[:@44973.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@44975.4]
  assign RetimeWrapper_4_io_in = _T_86 & _T_91; // @[package.scala 94:16:@44974.4]
  assign RetimeWrapper_5_clock = clock; // @[:@44980.4]
  assign RetimeWrapper_5_reset = reset; // @[:@44981.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@44983.4]
  assign RetimeWrapper_5_io_in = reset; // @[package.scala 94:16:@44982.4]
  assign RetimeWrapper_6_clock = clock; // @[:@44989.4]
  assign RetimeWrapper_6_reset = reset; // @[:@44990.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@44992.4]
  assign RetimeWrapper_6_io_in = _T_86 & _T_91; // @[package.scala 94:16:@44991.4]
  assign RetimeWrapper_7_clock = clock; // @[:@44997.4]
  assign RetimeWrapper_7_reset = reset; // @[:@44998.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@45000.4]
  assign RetimeWrapper_7_io_in = reset; // @[package.scala 94:16:@44999.4]
  assign RetimeWrapper_8_clock = clock; // @[:@45008.4]
  assign RetimeWrapper_8_reset = reset; // @[:@45009.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@45011.4]
  assign RetimeWrapper_8_io_in = _T_86 & _T_91; // @[package.scala 94:16:@45010.4]
  assign RetimeWrapper_9_clock = clock; // @[:@45016.4]
  assign RetimeWrapper_9_reset = reset; // @[:@45017.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@45019.4]
  assign RetimeWrapper_9_io_in = reset; // @[package.scala 94:16:@45018.4]
  assign RetimeWrapper_10_clock = clock; // @[:@45025.4]
  assign RetimeWrapper_10_reset = reset; // @[:@45026.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@45028.4]
  assign RetimeWrapper_10_io_in = _T_86 & _T_91; // @[package.scala 94:16:@45027.4]
  assign RetimeWrapper_11_clock = clock; // @[:@45033.4]
  assign RetimeWrapper_11_reset = reset; // @[:@45034.4]
  assign RetimeWrapper_11_io_flow = 1'h1; // @[package.scala 95:18:@45036.4]
  assign RetimeWrapper_11_io_in = reset; // @[package.scala 94:16:@45035.4]
  assign NBufCtr_clock = clock; // @[:@45058.4]
  assign NBufCtr_reset = reset; // @[:@45059.4]
  assign NBufCtr_io_input_enable = _T_86 & _T_91; // @[NBuffers.scala 42:23:@45065.4]
  assign statesInR_0_clock = clock; // @[:@45069.4]
  assign statesInR_0_reset = reset; // @[:@45070.4]
  assign statesInR_0_io_input_enable = _T_86 & _T_91; // @[NBuffers.scala 52:23:@45076.4]
  assign statesInR_1_clock = clock; // @[:@45080.4]
  assign statesInR_1_reset = reset; // @[:@45081.4]
  assign statesInR_1_io_input_enable = _T_86 & _T_91; // @[NBuffers.scala 52:23:@45087.4]
  assign statesInR_2_clock = clock; // @[:@45091.4]
  assign statesInR_2_reset = reset; // @[:@45092.4]
  assign statesInR_2_io_input_enable = _T_86 & _T_91; // @[NBuffers.scala 52:23:@45098.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_91 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_91 <= 1'h0;
    end else begin
      _T_91 <= _T_88;
    end
  end
endmodule
module Mem1D_39( // @[:@45166.2]
  input         clock, // @[:@45167.4]
  input         reset, // @[:@45168.4]
  input         io_r_ofs_0, // @[:@45169.4]
  input         io_r_backpressure, // @[:@45169.4]
  input         io_w_ofs_0, // @[:@45169.4]
  input  [31:0] io_w_data_0, // @[:@45169.4]
  input         io_w_en_0, // @[:@45169.4]
  output [31:0] io_output // @[:@45169.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@45179.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@45179.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@45179.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@45179.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@45179.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@45188.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@45188.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@45188.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@45188.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@45188.4]
  reg [31:0] _T_127; // @[MemPrimitives.scala 746:26:@45173.4]
  reg [31:0] _RAND_0;
  wire  _T_130; // @[MemPrimitives.scala 747:61:@45175.4]
  wire  _T_131; // @[MemPrimitives.scala 747:44:@45176.4]
  wire [31:0] _T_132; // @[MemPrimitives.scala 747:19:@45177.4]
  wire  _T_135; // @[package.scala 96:25:@45184.4 package.scala 96:25:@45185.4]
  wire  _T_137; // @[Mux.scala 46:19:@45186.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@45179.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_31 RetimeWrapper_1 ( // @[package.scala 93:22:@45188.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_130 = io_w_ofs_0 == 1'h0; // @[MemPrimitives.scala 747:61:@45175.4]
  assign _T_131 = io_w_en_0 & _T_130; // @[MemPrimitives.scala 747:44:@45176.4]
  assign _T_132 = _T_131 ? io_w_data_0 : _T_127; // @[MemPrimitives.scala 747:19:@45177.4]
  assign _T_135 = RetimeWrapper_io_out; // @[package.scala 96:25:@45184.4 package.scala 96:25:@45185.4]
  assign _T_137 = 1'h0 == _T_135; // @[Mux.scala 46:19:@45186.4]
  assign io_output = RetimeWrapper_1_io_out; // @[MemPrimitives.scala 751:17:@45195.4]
  assign RetimeWrapper_clock = clock; // @[:@45180.4]
  assign RetimeWrapper_reset = reset; // @[:@45181.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@45183.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@45182.4]
  assign RetimeWrapper_1_clock = clock; // @[:@45189.4]
  assign RetimeWrapper_1_reset = reset; // @[:@45190.4]
  assign RetimeWrapper_1_io_flow = io_r_backpressure; // @[package.scala 95:18:@45192.4]
  assign RetimeWrapper_1_io_in = _T_137 ? _T_127 : 32'h0; // @[package.scala 94:16:@45191.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_127 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_127 <= 32'h0;
    end else begin
      if (_T_131) begin
        _T_127 <= io_w_data_0;
      end
    end
  end
endmodule
module StickySelects_38( // @[:@45197.2]
  input   clock, // @[:@45198.4]
  input   reset, // @[:@45199.4]
  input   io_ins_0, // @[:@45200.4]
  input   io_ins_1, // @[:@45200.4]
  output  io_outs_0, // @[:@45200.4]
  output  io_outs_1 // @[:@45200.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@45202.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@45203.4]
  reg [31:0] _RAND_1;
  wire  _T_23; // @[StickySelects.scala 49:53:@45204.4]
  wire  _T_24; // @[StickySelects.scala 49:21:@45205.4]
  wire  _T_25; // @[StickySelects.scala 49:53:@45207.4]
  wire  _T_26; // @[StickySelects.scala 49:21:@45208.4]
  assign _T_23 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@45204.4]
  assign _T_24 = io_ins_1 ? io_ins_0 : _T_23; // @[StickySelects.scala 49:21:@45205.4]
  assign _T_25 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@45207.4]
  assign _T_26 = io_ins_0 ? io_ins_1 : _T_25; // @[StickySelects.scala 49:21:@45208.4]
  assign io_outs_0 = io_ins_1 ? io_ins_0 : _T_23; // @[StickySelects.scala 53:57:@45210.4]
  assign io_outs_1 = io_ins_0 ? io_ins_1 : _T_25; // @[StickySelects.scala 53:57:@45211.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (io_ins_1) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_23;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (io_ins_0) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_25;
      end
    end
  end
endmodule
module SRAM_71( // @[:@45277.2]
  input         clock, // @[:@45278.4]
  input         reset, // @[:@45279.4]
  input         io_rPort_1_en_0, // @[:@45280.4]
  output [31:0] io_rPort_1_output_0, // @[:@45280.4]
  input         io_rPort_0_en_0, // @[:@45280.4]
  output [31:0] io_rPort_0_output_0, // @[:@45280.4]
  input  [31:0] io_wPort_0_data_0, // @[:@45280.4]
  input         io_wPort_0_en_0 // @[:@45280.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@45300.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@45300.4]
  wire  Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@45300.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@45300.4]
  wire  Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@45300.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@45300.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@45300.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@45300.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@45327.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@45327.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@45327.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@45327.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@45327.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@45327.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@45346.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@45346.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@45346.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@45346.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@45346.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@45355.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@45355.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@45355.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@45355.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@45355.4]
  wire [33:0] _T_96; // @[Cat.scala 30:58:@45318.4]
  wire  _T_104; // @[MemPrimitives.scala 126:35:@45332.4]
  wire  _T_105; // @[MemPrimitives.scala 126:35:@45333.4]
  wire [2:0] _T_107; // @[Cat.scala 30:58:@45335.4]
  wire [2:0] _T_109; // @[Cat.scala 30:58:@45337.4]
  wire [2:0] _T_110; // @[Mux.scala 31:69:@45338.4]
  Mem1D_39 Mem1D ( // @[MemPrimitives.scala 64:21:@45300.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  StickySelects_38 StickySelects ( // @[MemPrimitives.scala 124:33:@45327.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@45346.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@45355.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_96 = {io_wPort_0_en_0,io_wPort_0_data_0,1'h0}; // @[Cat.scala 30:58:@45318.4]
  assign _T_104 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@45332.4]
  assign _T_105 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@45333.4]
  assign _T_107 = {_T_104,1'h1,1'h0}; // @[Cat.scala 30:58:@45335.4]
  assign _T_109 = {_T_105,1'h1,1'h0}; // @[Cat.scala 30:58:@45337.4]
  assign _T_110 = _T_104 ? _T_107 : _T_109; // @[Mux.scala 31:69:@45338.4]
  assign io_rPort_1_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@45362.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@45353.4]
  assign Mem1D_clock = clock; // @[:@45301.4]
  assign Mem1D_reset = reset; // @[:@45302.4]
  assign Mem1D_io_r_ofs_0 = _T_110[0]; // @[MemPrimitives.scala 131:28:@45342.4]
  assign Mem1D_io_r_backpressure = _T_110[1]; // @[MemPrimitives.scala 132:32:@45343.4]
  assign Mem1D_io_w_ofs_0 = _T_96[0]; // @[MemPrimitives.scala 94:28:@45322.4]
  assign Mem1D_io_w_data_0 = _T_96[32:1]; // @[MemPrimitives.scala 95:29:@45323.4]
  assign Mem1D_io_w_en_0 = _T_96[33]; // @[MemPrimitives.scala 96:27:@45324.4]
  assign StickySelects_clock = clock; // @[:@45328.4]
  assign StickySelects_reset = reset; // @[:@45329.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@45330.4]
  assign StickySelects_io_ins_1 = io_rPort_1_en_0; // @[MemPrimitives.scala 125:64:@45331.4]
  assign RetimeWrapper_clock = clock; // @[:@45347.4]
  assign RetimeWrapper_reset = reset; // @[:@45348.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@45350.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@45349.4]
  assign RetimeWrapper_1_clock = clock; // @[:@45356.4]
  assign RetimeWrapper_1_reset = reset; // @[:@45357.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@45359.4]
  assign RetimeWrapper_1_io_in = io_rPort_1_en_0; // @[package.scala 94:16:@45358.4]
endmodule
module x580_r_0( // @[:@45888.2]
  input         clock, // @[:@45889.4]
  input         reset, // @[:@45890.4]
  input         io_rPort_1_en_0, // @[:@45891.4]
  output [31:0] io_rPort_1_output_0, // @[:@45891.4]
  input         io_rPort_0_en_0, // @[:@45891.4]
  output [31:0] io_rPort_0_output_0, // @[:@45891.4]
  input  [31:0] io_wPort_0_data_0, // @[:@45891.4]
  input         io_wPort_0_en_0, // @[:@45891.4]
  input         io_sEn_0, // @[:@45891.4]
  input         io_sEn_1, // @[:@45891.4]
  input         io_sEn_2, // @[:@45891.4]
  input         io_sDone_0, // @[:@45891.4]
  input         io_sDone_1, // @[:@45891.4]
  input         io_sDone_2 // @[:@45891.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@45901.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@45901.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@45901.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@45901.4]
  wire  ctrl_io_sEn_2; // @[NBuffers.scala 83:20:@45901.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@45901.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@45901.4]
  wire  ctrl_io_sDone_2; // @[NBuffers.scala 83:20:@45901.4]
  wire [2:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@45901.4]
  wire [2:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@45901.4]
  wire [2:0] ctrl_io_statesInR_2; // @[NBuffers.scala 83:20:@45901.4]
  wire  SRAM_clock; // @[NBuffers.scala 94:23:@45910.4]
  wire  SRAM_reset; // @[NBuffers.scala 94:23:@45910.4]
  wire  SRAM_io_rPort_1_en_0; // @[NBuffers.scala 94:23:@45910.4]
  wire [31:0] SRAM_io_rPort_1_output_0; // @[NBuffers.scala 94:23:@45910.4]
  wire  SRAM_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@45910.4]
  wire [31:0] SRAM_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@45910.4]
  wire [31:0] SRAM_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@45910.4]
  wire  SRAM_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@45910.4]
  wire  SRAM_1_clock; // @[NBuffers.scala 94:23:@45931.4]
  wire  SRAM_1_reset; // @[NBuffers.scala 94:23:@45931.4]
  wire  SRAM_1_io_rPort_1_en_0; // @[NBuffers.scala 94:23:@45931.4]
  wire [31:0] SRAM_1_io_rPort_1_output_0; // @[NBuffers.scala 94:23:@45931.4]
  wire  SRAM_1_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@45931.4]
  wire [31:0] SRAM_1_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@45931.4]
  wire [31:0] SRAM_1_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@45931.4]
  wire  SRAM_1_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@45931.4]
  wire  SRAM_2_clock; // @[NBuffers.scala 94:23:@45952.4]
  wire  SRAM_2_reset; // @[NBuffers.scala 94:23:@45952.4]
  wire  SRAM_2_io_rPort_1_en_0; // @[NBuffers.scala 94:23:@45952.4]
  wire [31:0] SRAM_2_io_rPort_1_output_0; // @[NBuffers.scala 94:23:@45952.4]
  wire  SRAM_2_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@45952.4]
  wire [31:0] SRAM_2_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@45952.4]
  wire [31:0] SRAM_2_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@45952.4]
  wire  SRAM_2_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@45952.4]
  wire  _T_140; // @[NBuffers.scala 104:105:@45973.4]
  wire  _T_144; // @[NBuffers.scala 108:92:@45983.4]
  wire  _T_147; // @[NBuffers.scala 108:92:@45989.4]
  wire  _T_150; // @[NBuffers.scala 104:105:@45995.4]
  wire  _T_154; // @[NBuffers.scala 108:92:@46005.4]
  wire  _T_157; // @[NBuffers.scala 108:92:@46011.4]
  wire  _T_160; // @[NBuffers.scala 104:105:@46017.4]
  wire  _T_164; // @[NBuffers.scala 108:92:@46027.4]
  wire  _T_167; // @[NBuffers.scala 108:92:@46033.4]
  wire [31:0] _T_177; // @[Mux.scala 19:72:@46042.4]
  wire [31:0] _T_179; // @[Mux.scala 19:72:@46043.4]
  wire [31:0] _T_181; // @[Mux.scala 19:72:@46044.4]
  wire [31:0] _T_182; // @[Mux.scala 19:72:@46045.4]
  wire [31:0] _T_194; // @[Mux.scala 19:72:@46053.4]
  wire [31:0] _T_196; // @[Mux.scala 19:72:@46054.4]
  wire [31:0] _T_198; // @[Mux.scala 19:72:@46055.4]
  wire [31:0] _T_199; // @[Mux.scala 19:72:@46056.4]
  NBufController_10 ctrl ( // @[NBuffers.scala 83:20:@45901.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sEn_2(ctrl_io_sEn_2),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_sDone_2(ctrl_io_sDone_2),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1),
    .io_statesInR_2(ctrl_io_statesInR_2)
  );
  SRAM_71 SRAM ( // @[NBuffers.scala 94:23:@45910.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_rPort_1_en_0(SRAM_io_rPort_1_en_0),
    .io_rPort_1_output_0(SRAM_io_rPort_1_output_0),
    .io_rPort_0_en_0(SRAM_io_rPort_0_en_0),
    .io_rPort_0_output_0(SRAM_io_rPort_0_output_0),
    .io_wPort_0_data_0(SRAM_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_io_wPort_0_en_0)
  );
  SRAM_71 SRAM_1 ( // @[NBuffers.scala 94:23:@45931.4]
    .clock(SRAM_1_clock),
    .reset(SRAM_1_reset),
    .io_rPort_1_en_0(SRAM_1_io_rPort_1_en_0),
    .io_rPort_1_output_0(SRAM_1_io_rPort_1_output_0),
    .io_rPort_0_en_0(SRAM_1_io_rPort_0_en_0),
    .io_rPort_0_output_0(SRAM_1_io_rPort_0_output_0),
    .io_wPort_0_data_0(SRAM_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_1_io_wPort_0_en_0)
  );
  SRAM_71 SRAM_2 ( // @[NBuffers.scala 94:23:@45952.4]
    .clock(SRAM_2_clock),
    .reset(SRAM_2_reset),
    .io_rPort_1_en_0(SRAM_2_io_rPort_1_en_0),
    .io_rPort_1_output_0(SRAM_2_io_rPort_1_output_0),
    .io_rPort_0_en_0(SRAM_2_io_rPort_0_en_0),
    .io_rPort_0_output_0(SRAM_2_io_rPort_0_output_0),
    .io_wPort_0_data_0(SRAM_2_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_2_io_wPort_0_en_0)
  );
  assign _T_140 = ctrl_io_statesInW_0 == 3'h0; // @[NBuffers.scala 104:105:@45973.4]
  assign _T_144 = ctrl_io_statesInR_1 == 3'h0; // @[NBuffers.scala 108:92:@45983.4]
  assign _T_147 = ctrl_io_statesInR_2 == 3'h0; // @[NBuffers.scala 108:92:@45989.4]
  assign _T_150 = ctrl_io_statesInW_0 == 3'h1; // @[NBuffers.scala 104:105:@45995.4]
  assign _T_154 = ctrl_io_statesInR_1 == 3'h1; // @[NBuffers.scala 108:92:@46005.4]
  assign _T_157 = ctrl_io_statesInR_2 == 3'h1; // @[NBuffers.scala 108:92:@46011.4]
  assign _T_160 = ctrl_io_statesInW_0 == 3'h2; // @[NBuffers.scala 104:105:@46017.4]
  assign _T_164 = ctrl_io_statesInR_1 == 3'h2; // @[NBuffers.scala 108:92:@46027.4]
  assign _T_167 = ctrl_io_statesInR_2 == 3'h2; // @[NBuffers.scala 108:92:@46033.4]
  assign _T_177 = _T_144 ? SRAM_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@46042.4]
  assign _T_179 = _T_154 ? SRAM_1_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@46043.4]
  assign _T_181 = _T_164 ? SRAM_2_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@46044.4]
  assign _T_182 = _T_177 | _T_179; // @[Mux.scala 19:72:@46045.4]
  assign _T_194 = _T_147 ? SRAM_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@46053.4]
  assign _T_196 = _T_157 ? SRAM_1_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@46054.4]
  assign _T_198 = _T_167 ? SRAM_2_io_rPort_1_output_0 : 32'h0; // @[Mux.scala 19:72:@46055.4]
  assign _T_199 = _T_194 | _T_196; // @[Mux.scala 19:72:@46056.4]
  assign io_rPort_1_output_0 = _T_199 | _T_198; // @[NBuffers.scala 115:66:@46060.4]
  assign io_rPort_0_output_0 = _T_182 | _T_181; // @[NBuffers.scala 115:66:@46049.4]
  assign ctrl_clock = clock; // @[:@45902.4]
  assign ctrl_reset = reset; // @[:@45903.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@45904.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@45906.4]
  assign ctrl_io_sEn_2 = io_sEn_2; // @[NBuffers.scala 85:20:@45908.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@45905.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@45907.4]
  assign ctrl_io_sDone_2 = io_sDone_2; // @[NBuffers.scala 86:22:@45909.4]
  assign SRAM_clock = clock; // @[:@45911.4]
  assign SRAM_reset = reset; // @[:@45912.4]
  assign SRAM_io_rPort_1_en_0 = io_rPort_1_en_0 & _T_147; // @[MemPrimitives.scala 43:33:@45993.4]
  assign SRAM_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_144; // @[MemPrimitives.scala 43:33:@45987.4]
  assign SRAM_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@45976.4]
  assign SRAM_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_140; // @[MemPrimitives.scala 37:29:@45982.4]
  assign SRAM_1_clock = clock; // @[:@45932.4]
  assign SRAM_1_reset = reset; // @[:@45933.4]
  assign SRAM_1_io_rPort_1_en_0 = io_rPort_1_en_0 & _T_157; // @[MemPrimitives.scala 43:33:@46015.4]
  assign SRAM_1_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_154; // @[MemPrimitives.scala 43:33:@46009.4]
  assign SRAM_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@45998.4]
  assign SRAM_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_150; // @[MemPrimitives.scala 37:29:@46004.4]
  assign SRAM_2_clock = clock; // @[:@45953.4]
  assign SRAM_2_reset = reset; // @[:@45954.4]
  assign SRAM_2_io_rPort_1_en_0 = io_rPort_1_en_0 & _T_167; // @[MemPrimitives.scala 43:33:@46037.4]
  assign SRAM_2_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_164; // @[MemPrimitives.scala 43:33:@46031.4]
  assign SRAM_2_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@46020.4]
  assign SRAM_2_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_160; // @[MemPrimitives.scala 37:29:@46026.4]
endmodule
module RetimeWrapper_516( // @[:@46100.2]
  input   clock, // @[:@46101.4]
  input   reset, // @[:@46102.4]
  input   io_in, // @[:@46103.4]
  output  io_out // @[:@46103.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@46105.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@46105.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@46105.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@46105.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@46105.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@46105.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@46105.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@46118.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@46117.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@46116.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@46115.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@46114.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@46112.4]
endmodule
module RetimeWrapper_520( // @[:@46228.2]
  input   clock, // @[:@46229.4]
  input   reset, // @[:@46230.4]
  input   io_flow, // @[:@46231.4]
  input   io_in, // @[:@46231.4]
  output  io_out // @[:@46231.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@46233.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@46233.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@46233.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@46233.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@46233.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@46233.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@46233.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@46246.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@46245.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@46244.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@46243.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@46242.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@46240.4]
endmodule
module x593_inr_UnitPipe_sm( // @[:@46248.2]
  input   clock, // @[:@46249.4]
  input   reset, // @[:@46250.4]
  input   io_enable, // @[:@46251.4]
  output  io_done, // @[:@46251.4]
  input   io_ctrDone, // @[:@46251.4]
  output  io_datapathEn, // @[:@46251.4]
  output  io_ctrInc, // @[:@46251.4]
  input   io_parentAck, // @[:@46251.4]
  input   io_backpressure, // @[:@46251.4]
  input   io_break // @[:@46251.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@46253.4]
  wire  active_reset; // @[Controllers.scala 261:22:@46253.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@46253.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@46253.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@46253.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@46253.4]
  wire  done_clock; // @[Controllers.scala 262:20:@46256.4]
  wire  done_reset; // @[Controllers.scala 262:20:@46256.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@46256.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@46256.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@46256.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@46256.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@46290.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@46290.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@46290.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@46290.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@46312.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@46312.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@46312.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@46312.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@46324.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@46324.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@46324.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@46324.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@46324.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@46332.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@46332.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@46332.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@46332.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@46332.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@46348.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@46348.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@46348.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@46348.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@46348.4]
  wire  _T_80; // @[Controllers.scala 264:48:@46261.4]
  wire  _T_81; // @[Controllers.scala 264:46:@46262.4]
  wire  _T_82; // @[Controllers.scala 264:62:@46263.4]
  wire  _T_100; // @[package.scala 100:49:@46281.4]
  reg  _T_103; // @[package.scala 48:56:@46282.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@46305.4]
  wire  _T_124; // @[package.scala 96:25:@46317.4 package.scala 96:25:@46318.4]
  wire  _T_126; // @[package.scala 100:49:@46319.4]
  reg  _T_129; // @[package.scala 48:56:@46320.4]
  reg [31:0] _RAND_1;
  wire  _T_150; // @[package.scala 100:49:@46344.4]
  reg  _T_153; // @[package.scala 48:56:@46345.4]
  reg [31:0] _RAND_2;
  SRFF active ( // @[Controllers.scala 261:22:@46253.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@46256.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_516 RetimeWrapper ( // @[package.scala 93:22:@46290.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_516 RetimeWrapper_1 ( // @[package.scala 93:22:@46312.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@46324.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@46332.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_520 RetimeWrapper_4 ( // @[package.scala 93:22:@46348.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@46261.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@46262.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@46263.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@46281.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@46305.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@46317.4 package.scala 96:25:@46318.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@46319.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@46344.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@46323.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@46308.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@46311.4]
  assign active_clock = clock; // @[:@46254.4]
  assign active_reset = reset; // @[:@46255.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@46266.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@46270.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@46271.4]
  assign done_clock = clock; // @[:@46257.4]
  assign done_reset = reset; // @[:@46258.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@46286.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@46279.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@46280.4]
  assign RetimeWrapper_clock = clock; // @[:@46291.4]
  assign RetimeWrapper_reset = reset; // @[:@46292.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@46293.4]
  assign RetimeWrapper_1_clock = clock; // @[:@46313.4]
  assign RetimeWrapper_1_reset = reset; // @[:@46314.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@46315.4]
  assign RetimeWrapper_2_clock = clock; // @[:@46325.4]
  assign RetimeWrapper_2_reset = reset; // @[:@46326.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@46328.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@46327.4]
  assign RetimeWrapper_3_clock = clock; // @[:@46333.4]
  assign RetimeWrapper_3_reset = reset; // @[:@46334.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@46336.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@46335.4]
  assign RetimeWrapper_4_clock = clock; // @[:@46349.4]
  assign RetimeWrapper_4_reset = reset; // @[:@46350.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@46352.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@46351.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_153 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module Multiplier( // @[:@46507.2]
  input         clock, // @[:@46508.4]
  input         io_flow, // @[:@46510.4]
  input  [53:0] io_a, // @[:@46510.4]
  input  [53:0] io_b, // @[:@46510.4]
  output [53:0] io_out // @[:@46510.4]
);
  wire [53:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@46512.4]
  wire [53:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@46512.4]
  wire [53:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@46512.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@46512.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@46512.4]
  mul_54_54_54_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@46512.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@46522.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@46520.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@46519.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@46521.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@46518.4]
endmodule
module fix2fixBox_53( // @[:@46588.2]
  input  [53:0] io_a, // @[:@46591.4]
  output [31:0] io_b // @[:@46591.4]
);
  wire [21:0] tmp_frac; // @[Converter.scala 38:42:@46599.4]
  wire [9:0] new_dec; // @[Converter.scala 88:34:@46602.4]
  assign tmp_frac = io_a[43:22]; // @[Converter.scala 38:42:@46599.4]
  assign new_dec = io_a[53:44]; // @[Converter.scala 88:34:@46602.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@46605.4]
endmodule
module x586_mul( // @[:@46607.2]
  input         clock, // @[:@46608.4]
  input         reset, // @[:@46609.4]
  input  [31:0] io_a, // @[:@46610.4]
  input  [31:0] io_b, // @[:@46610.4]
  input         io_flow, // @[:@46610.4]
  output [31:0] io_result // @[:@46610.4]
);
  wire  x586_mul_clock; // @[BigIPZynq.scala 63:21:@46625.4]
  wire  x586_mul_io_flow; // @[BigIPZynq.scala 63:21:@46625.4]
  wire [53:0] x586_mul_io_a; // @[BigIPZynq.scala 63:21:@46625.4]
  wire [53:0] x586_mul_io_b; // @[BigIPZynq.scala 63:21:@46625.4]
  wire [53:0] x586_mul_io_out; // @[BigIPZynq.scala 63:21:@46625.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@46636.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@46636.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@46636.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@46636.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@46636.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@46647.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@46647.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@46647.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@46647.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@46647.4]
  wire [53:0] fix2fixBox_io_a; // @[Math.scala 253:30:@46654.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@46654.4]
  wire  _T_16; // @[FixedPoint.scala 50:25:@46617.4]
  wire [21:0] _T_20; // @[Bitwise.scala 72:12:@46619.4]
  wire  _T_22; // @[FixedPoint.scala 50:25:@46621.4]
  wire [21:0] _T_26; // @[Bitwise.scala 72:12:@46623.4]
  wire  _T_31; // @[Math.scala 251:56:@46635.4]
  Multiplier x586_mul ( // @[BigIPZynq.scala 63:21:@46625.4]
    .clock(x586_mul_clock),
    .io_flow(x586_mul_io_flow),
    .io_a(x586_mul_io_a),
    .io_b(x586_mul_io_b),
    .io_out(x586_mul_io_out)
  );
  RetimeWrapper_451 RetimeWrapper ( // @[package.scala 93:22:@46636.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_451 RetimeWrapper_1 ( // @[package.scala 93:22:@46647.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  fix2fixBox_53 fix2fixBox ( // @[Math.scala 253:30:@46654.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_16 = io_a[31]; // @[FixedPoint.scala 50:25:@46617.4]
  assign _T_20 = _T_16 ? 22'h3fffff : 22'h0; // @[Bitwise.scala 72:12:@46619.4]
  assign _T_22 = io_b[31]; // @[FixedPoint.scala 50:25:@46621.4]
  assign _T_26 = _T_22 ? 22'h3fffff : 22'h0; // @[Bitwise.scala 72:12:@46623.4]
  assign _T_31 = _T_16 ^ _T_22; // @[Math.scala 251:56:@46635.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@46662.4]
  assign x586_mul_clock = clock; // @[:@46626.4]
  assign x586_mul_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@46630.4]
  assign x586_mul_io_a = {_T_20,io_a}; // @[BigIPZynq.scala 64:14:@46628.4]
  assign x586_mul_io_b = {_T_26,io_b}; // @[BigIPZynq.scala 65:14:@46629.4]
  assign RetimeWrapper_clock = clock; // @[:@46637.4]
  assign RetimeWrapper_reset = reset; // @[:@46638.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@46640.4]
  assign RetimeWrapper_io_in = _T_16 ^ _T_22; // @[package.scala 94:16:@46639.4]
  assign RetimeWrapper_1_clock = clock; // @[:@46648.4]
  assign RetimeWrapper_1_reset = reset; // @[:@46649.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@46651.4]
  assign RetimeWrapper_1_io_in = _T_31 == 1'h0; // @[package.scala 94:16:@46650.4]
  assign fix2fixBox_io_a = x586_mul_io_out; // @[Math.scala 254:23:@46657.4]
endmodule
module RetimeWrapper_527( // @[:@46676.2]
  input         clock, // @[:@46677.4]
  input         reset, // @[:@46678.4]
  input         io_flow, // @[:@46679.4]
  input  [31:0] io_in, // @[:@46679.4]
  output [31:0] io_out // @[:@46679.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@46681.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@46681.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@46681.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@46681.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@46681.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@46681.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@46681.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@46694.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@46693.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@46692.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@46691.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@46690.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@46688.4]
endmodule
module fix2fixBox_57( // @[:@46973.2]
  input  [32:0] io_a, // @[:@46976.4]
  output [31:0] io_b // @[:@46976.4]
);
  wire [21:0] tmp_frac; // @[Converter.scala 52:23:@46984.4]
  wire [9:0] new_dec; // @[Converter.scala 63:26:@46987.4]
  assign tmp_frac = io_a[21:0]; // @[Converter.scala 52:23:@46984.4]
  assign new_dec = io_a[31:22]; // @[Converter.scala 63:26:@46987.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@46990.4]
endmodule
module add( // @[:@46992.2]
  input  [31:0] io_a, // @[:@46995.4]
  input  [31:0] io_b, // @[:@46995.4]
  output [31:0] io_result // @[:@46995.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@47003.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@47003.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@47010.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@47010.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@47028.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@47028.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@47008.4 Math.scala 724:14:@47009.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@47015.4 Math.scala 724:14:@47016.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@47017.4]
  __37 _ ( // @[Math.scala 720:24:@47003.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __37 __1 ( // @[Math.scala 720:24:@47010.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_57 fix2fixBox ( // @[Math.scala 141:30:@47028.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@47008.4 Math.scala 724:14:@47009.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@47015.4 Math.scala 724:14:@47016.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@47017.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@47036.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@47006.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@47013.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@47031.4]
endmodule
module x748( // @[:@47038.2]
  input         clock, // @[:@47039.4]
  input         reset, // @[:@47040.4]
  input  [31:0] io_m0, // @[:@47041.4]
  input  [31:0] io_m1, // @[:@47041.4]
  input  [31:0] io_add, // @[:@47041.4]
  output [31:0] io_result // @[:@47041.4]
);
  wire  fmamul_x748_clock; // @[Math.scala 262:24:@47049.4]
  wire  fmamul_x748_reset; // @[Math.scala 262:24:@47049.4]
  wire [31:0] fmamul_x748_io_a; // @[Math.scala 262:24:@47049.4]
  wire [31:0] fmamul_x748_io_b; // @[Math.scala 262:24:@47049.4]
  wire  fmamul_x748_io_flow; // @[Math.scala 262:24:@47049.4]
  wire [31:0] fmamul_x748_io_result; // @[Math.scala 262:24:@47049.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@47057.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@47057.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@47057.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@47057.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@47057.4]
  wire [31:0] add_1_io_a; // @[Math.scala 150:24:@47067.4]
  wire [31:0] add_1_io_b; // @[Math.scala 150:24:@47067.4]
  wire [31:0] add_1_io_result; // @[Math.scala 150:24:@47067.4]
  x586_mul fmamul_x748 ( // @[Math.scala 262:24:@47049.4]
    .clock(fmamul_x748_clock),
    .reset(fmamul_x748_reset),
    .io_a(fmamul_x748_io_a),
    .io_b(fmamul_x748_io_b),
    .io_flow(fmamul_x748_io_flow),
    .io_result(fmamul_x748_io_result)
  );
  RetimeWrapper_527 RetimeWrapper ( // @[package.scala 93:22:@47057.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  add add_1 ( // @[Math.scala 150:24:@47067.4]
    .io_a(add_1_io_a),
    .io_b(add_1_io_b),
    .io_result(add_1_io_result)
  );
  assign io_result = add_1_io_result; // @[Math.scala 857:17:@47075.4]
  assign fmamul_x748_clock = clock; // @[:@47050.4]
  assign fmamul_x748_reset = reset; // @[:@47051.4]
  assign fmamul_x748_io_a = io_m0; // @[Math.scala 263:17:@47052.4]
  assign fmamul_x748_io_b = io_m1; // @[Math.scala 264:17:@47053.4]
  assign fmamul_x748_io_flow = 1'h1; // @[Math.scala 265:20:@47054.4]
  assign RetimeWrapper_clock = clock; // @[:@47058.4]
  assign RetimeWrapper_reset = reset; // @[:@47059.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@47061.4]
  assign RetimeWrapper_io_in = io_add; // @[package.scala 94:16:@47060.4]
  assign add_1_io_a = fmamul_x748_io_result; // @[Math.scala 151:17:@47070.4]
  assign add_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@47071.4]
endmodule
module fix2fixBox_58( // @[:@47077.2]
  input  [31:0] io_a, // @[:@47080.4]
  output [31:0] io_b // @[:@47080.4]
);
  wire [21:0] tmp_frac; // @[Converter.scala 52:23:@47088.4]
  wire [9:0] new_dec; // @[Converter.scala 88:34:@47091.4]
  assign tmp_frac = io_a[21:0]; // @[Converter.scala 52:23:@47088.4]
  assign new_dec = io_a[31:22]; // @[Converter.scala 88:34:@47091.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@47094.4]
endmodule
module cast_x748( // @[:@47096.2]
  input  [31:0] io_b, // @[:@47099.4]
  output [31:0] io_result // @[:@47099.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@47104.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@47104.4]
  fix2fixBox_58 fix2fixBox ( // @[BigIPZynq.scala 219:30:@47104.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@47112.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@47107.4]
endmodule
module RetimeWrapper_531( // @[:@47126.2]
  input         clock, // @[:@47127.4]
  input         reset, // @[:@47128.4]
  input  [31:0] io_in, // @[:@47129.4]
  output [31:0] io_out // @[:@47129.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@47131.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@47131.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@47131.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@47131.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@47131.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@47131.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(12)) sr ( // @[RetimeShiftRegister.scala 15:20:@47131.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@47144.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@47143.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@47142.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@47141.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@47140.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@47138.4]
endmodule
module x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1( // @[:@47788.2]
  input         clock, // @[:@47789.4]
  input         reset, // @[:@47790.4]
  output        io_in_x555_tmp_1_rPort_0_en_0, // @[:@47791.4]
  input  [31:0] io_in_x555_tmp_1_rPort_0_output_0, // @[:@47791.4]
  output        io_in_x555_tmp_1_sEn_1, // @[:@47791.4]
  output        io_in_x555_tmp_1_sDone_1, // @[:@47791.4]
  output        io_in_x554_tmp_0_rPort_0_en_0, // @[:@47791.4]
  input  [31:0] io_in_x554_tmp_0_rPort_0_output_0, // @[:@47791.4]
  output        io_in_x554_tmp_0_sEn_1, // @[:@47791.4]
  output        io_in_x554_tmp_0_sDone_1, // @[:@47791.4]
  output        io_in_x558_tmp_4_sEn_1, // @[:@47791.4]
  output        io_in_x558_tmp_4_sDone_1, // @[:@47791.4]
  output        io_in_x557_tmp_3_sEn_1, // @[:@47791.4]
  output        io_in_x557_tmp_3_sDone_1, // @[:@47791.4]
  output [31:0] io_in_x580_r_0_wPort_0_data_0, // @[:@47791.4]
  output        io_in_x580_r_0_wPort_0_en_0, // @[:@47791.4]
  output        io_in_x580_r_0_sEn_0, // @[:@47791.4]
  output        io_in_x580_r_0_sDone_0, // @[:@47791.4]
  output        io_in_x556_tmp_2_rPort_0_en_0, // @[:@47791.4]
  input  [31:0] io_in_x556_tmp_2_rPort_0_output_0, // @[:@47791.4]
  output        io_in_x556_tmp_2_sEn_1, // @[:@47791.4]
  output        io_in_x556_tmp_2_sDone_1, // @[:@47791.4]
  input         io_sigsIn_done, // @[:@47791.4]
  input         io_sigsIn_datapathEn, // @[:@47791.4]
  input         io_sigsIn_baseEn, // @[:@47791.4]
  input         io_sigsIn_break, // @[:@47791.4]
  input         io_rr // @[:@47791.4]
);
  wire  x586_mul_1_clock; // @[Math.scala 262:24:@48098.4]
  wire  x586_mul_1_reset; // @[Math.scala 262:24:@48098.4]
  wire [31:0] x586_mul_1_io_a; // @[Math.scala 262:24:@48098.4]
  wire [31:0] x586_mul_1_io_b; // @[Math.scala 262:24:@48098.4]
  wire  x586_mul_1_io_flow; // @[Math.scala 262:24:@48098.4]
  wire [31:0] x586_mul_1_io_result; // @[Math.scala 262:24:@48098.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@48109.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@48109.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@48109.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@48109.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@48109.4]
  wire  x748_1_clock; // @[Math.scala 860:24:@48118.4]
  wire  x748_1_reset; // @[Math.scala 860:24:@48118.4]
  wire [31:0] x748_1_io_m0; // @[Math.scala 860:24:@48118.4]
  wire [31:0] x748_1_io_m1; // @[Math.scala 860:24:@48118.4]
  wire [31:0] x748_1_io_add; // @[Math.scala 860:24:@48118.4]
  wire [31:0] x748_1_io_result; // @[Math.scala 860:24:@48118.4]
  wire [31:0] cast_x748_io_b; // @[Math.scala 720:24:@48127.4]
  wire [31:0] cast_x748_io_result; // @[Math.scala 720:24:@48127.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@48159.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@48159.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@48159.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@48159.4]
  wire  x749_1_clock; // @[Math.scala 860:24:@48168.4]
  wire  x749_1_reset; // @[Math.scala 860:24:@48168.4]
  wire [31:0] x749_1_io_m0; // @[Math.scala 860:24:@48168.4]
  wire [31:0] x749_1_io_m1; // @[Math.scala 860:24:@48168.4]
  wire [31:0] x749_1_io_add; // @[Math.scala 860:24:@48168.4]
  wire [31:0] x749_1_io_result; // @[Math.scala 860:24:@48168.4]
  wire [31:0] cast_x749_io_b; // @[Math.scala 720:24:@48177.4]
  wire [31:0] cast_x749_io_result; // @[Math.scala 720:24:@48177.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@48193.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@48193.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@48193.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@48193.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@48193.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@48212.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@48212.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@48212.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@48212.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@48212.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@48223.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@48223.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@48223.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@48223.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@48223.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@48234.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@48234.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@48234.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@48234.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@48234.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@48245.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@48245.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@48245.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@48245.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@48245.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@48256.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@48256.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@48256.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@48256.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@48256.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@48267.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@48267.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@48267.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@48267.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@48267.4]
  wire  _T_1839; // @[sm_x593_inr_UnitPipe.scala 89:114:@48060.4]
  wire  _T_1840; // @[sm_x593_inr_UnitPipe.scala 89:111:@48061.4]
  wire  _T_1845; // @[implicits.scala 56:10:@48064.4]
  wire  _T_1950; // @[package.scala 96:25:@48198.4 package.scala 96:25:@48199.4]
  wire  _T_1952; // @[implicits.scala 56:10:@48200.4]
  wire  _T_1953; // @[sm_x593_inr_UnitPipe.scala 126:113:@48201.4]
  wire  _T_1962; // @[package.scala 96:25:@48217.4 package.scala 96:25:@48218.4]
  wire  _T_1968; // @[package.scala 96:25:@48228.4 package.scala 96:25:@48229.4]
  wire  _T_1974; // @[package.scala 96:25:@48239.4 package.scala 96:25:@48240.4]
  wire  _T_1980; // @[package.scala 96:25:@48250.4 package.scala 96:25:@48251.4]
  wire  _T_1986; // @[package.scala 96:25:@48261.4 package.scala 96:25:@48262.4]
  wire  _T_1992; // @[package.scala 96:25:@48272.4 package.scala 96:25:@48273.4]
  x586_mul x586_mul_1 ( // @[Math.scala 262:24:@48098.4]
    .clock(x586_mul_1_clock),
    .reset(x586_mul_1_reset),
    .io_a(x586_mul_1_io_a),
    .io_b(x586_mul_1_io_b),
    .io_flow(x586_mul_1_io_flow),
    .io_result(x586_mul_1_io_result)
  );
  RetimeWrapper_527 RetimeWrapper ( // @[package.scala 93:22:@48109.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x748 x748_1 ( // @[Math.scala 860:24:@48118.4]
    .clock(x748_1_clock),
    .reset(x748_1_reset),
    .io_m0(x748_1_io_m0),
    .io_m1(x748_1_io_m1),
    .io_add(x748_1_io_add),
    .io_result(x748_1_io_result)
  );
  cast_x748 cast_x748 ( // @[Math.scala 720:24:@48127.4]
    .io_b(cast_x748_io_b),
    .io_result(cast_x748_io_result)
  );
  RetimeWrapper_531 RetimeWrapper_1 ( // @[package.scala 93:22:@48159.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x748 x749_1 ( // @[Math.scala 860:24:@48168.4]
    .clock(x749_1_clock),
    .reset(x749_1_reset),
    .io_m0(x749_1_io_m0),
    .io_m1(x749_1_io_m1),
    .io_add(x749_1_io_add),
    .io_result(x749_1_io_result)
  );
  cast_x748 cast_x749 ( // @[Math.scala 720:24:@48177.4]
    .io_b(cast_x749_io_b),
    .io_result(cast_x749_io_result)
  );
  RetimeWrapper_520 RetimeWrapper_2 ( // @[package.scala 93:22:@48193.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@48212.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@48223.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@48234.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@48245.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@48256.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@48267.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  assign _T_1839 = ~ io_sigsIn_break; // @[sm_x593_inr_UnitPipe.scala 89:114:@48060.4]
  assign _T_1840 = io_rr & _T_1839; // @[sm_x593_inr_UnitPipe.scala 89:111:@48061.4]
  assign _T_1845 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 56:10:@48064.4]
  assign _T_1950 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@48198.4 package.scala 96:25:@48199.4]
  assign _T_1952 = io_rr ? _T_1950 : 1'h0; // @[implicits.scala 56:10:@48200.4]
  assign _T_1953 = _T_1839 & _T_1952; // @[sm_x593_inr_UnitPipe.scala 126:113:@48201.4]
  assign _T_1962 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@48217.4 package.scala 96:25:@48218.4]
  assign _T_1968 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@48228.4 package.scala 96:25:@48229.4]
  assign _T_1974 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@48239.4 package.scala 96:25:@48240.4]
  assign _T_1980 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@48250.4 package.scala 96:25:@48251.4]
  assign _T_1986 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@48261.4 package.scala 96:25:@48262.4]
  assign _T_1992 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@48272.4 package.scala 96:25:@48273.4]
  assign io_in_x555_tmp_1_rPort_0_en_0 = _T_1840 & _T_1845; // @[MemInterfaceType.scala 110:79:@48093.4]
  assign io_in_x555_tmp_1_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@48231.4]
  assign io_in_x555_tmp_1_sDone_1 = io_rr ? _T_1968 : 1'h0; // @[MemInterfaceType.scala 197:17:@48232.4]
  assign io_in_x554_tmp_0_rPort_0_en_0 = _T_1840 & _T_1845; // @[MemInterfaceType.scala 110:79:@48071.4]
  assign io_in_x554_tmp_0_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@48220.4]
  assign io_in_x554_tmp_0_sDone_1 = io_rr ? _T_1962 : 1'h0; // @[MemInterfaceType.scala 197:17:@48221.4]
  assign io_in_x558_tmp_4_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@48264.4]
  assign io_in_x558_tmp_4_sDone_1 = io_rr ? _T_1986 : 1'h0; // @[MemInterfaceType.scala 197:17:@48265.4]
  assign io_in_x557_tmp_3_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@48253.4]
  assign io_in_x557_tmp_3_sDone_1 = io_rr ? _T_1980 : 1'h0; // @[MemInterfaceType.scala 197:17:@48254.4]
  assign io_in_x580_r_0_wPort_0_data_0 = cast_x749_io_result; // @[MemInterfaceType.scala 90:56:@48208.4]
  assign io_in_x580_r_0_wPort_0_en_0 = _T_1953 & _T_1839; // @[MemInterfaceType.scala 93:57:@48210.4]
  assign io_in_x580_r_0_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@48275.4]
  assign io_in_x580_r_0_sDone_0 = io_rr ? _T_1992 : 1'h0; // @[MemInterfaceType.scala 197:17:@48276.4]
  assign io_in_x556_tmp_2_rPort_0_en_0 = _T_1840 & _T_1845; // @[MemInterfaceType.scala 110:79:@48153.4]
  assign io_in_x556_tmp_2_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@48242.4]
  assign io_in_x556_tmp_2_sDone_1 = io_rr ? _T_1974 : 1'h0; // @[MemInterfaceType.scala 197:17:@48243.4]
  assign x586_mul_1_clock = clock; // @[:@48099.4]
  assign x586_mul_1_reset = reset; // @[:@48100.4]
  assign x586_mul_1_io_a = io_in_x555_tmp_1_rPort_0_output_0; // @[Math.scala 263:17:@48101.4]
  assign x586_mul_1_io_b = io_in_x555_tmp_1_rPort_0_output_0; // @[Math.scala 264:17:@48102.4]
  assign x586_mul_1_io_flow = 1'h1; // @[Math.scala 265:20:@48103.4]
  assign RetimeWrapper_clock = clock; // @[:@48110.4]
  assign RetimeWrapper_reset = reset; // @[:@48111.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@48113.4]
  assign RetimeWrapper_io_in = io_in_x554_tmp_0_rPort_0_output_0; // @[package.scala 94:16:@48112.4]
  assign x748_1_clock = clock; // @[:@48119.4]
  assign x748_1_reset = reset; // @[:@48120.4]
  assign x748_1_io_m0 = RetimeWrapper_io_out; // @[Math.scala 861:18:@48121.4]
  assign x748_1_io_m1 = RetimeWrapper_io_out; // @[Math.scala 862:18:@48122.4]
  assign x748_1_io_add = x586_mul_1_io_result; // @[Math.scala 863:19:@48123.4]
  assign cast_x748_io_b = x748_1_io_result; // @[Math.scala 721:17:@48130.4]
  assign RetimeWrapper_1_clock = clock; // @[:@48160.4]
  assign RetimeWrapper_1_reset = reset; // @[:@48161.4]
  assign RetimeWrapper_1_io_in = io_in_x556_tmp_2_rPort_0_output_0; // @[package.scala 94:16:@48162.4]
  assign x749_1_clock = clock; // @[:@48169.4]
  assign x749_1_reset = reset; // @[:@48170.4]
  assign x749_1_io_m0 = RetimeWrapper_1_io_out; // @[Math.scala 861:18:@48171.4]
  assign x749_1_io_m1 = RetimeWrapper_1_io_out; // @[Math.scala 862:18:@48172.4]
  assign x749_1_io_add = cast_x748_io_result; // @[Math.scala 863:19:@48173.4]
  assign cast_x749_io_b = x749_1_io_result; // @[Math.scala 721:17:@48180.4]
  assign RetimeWrapper_2_clock = clock; // @[:@48194.4]
  assign RetimeWrapper_2_reset = reset; // @[:@48195.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@48197.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@48196.4]
  assign RetimeWrapper_3_clock = clock; // @[:@48213.4]
  assign RetimeWrapper_3_reset = reset; // @[:@48214.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@48216.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_done; // @[package.scala 94:16:@48215.4]
  assign RetimeWrapper_4_clock = clock; // @[:@48224.4]
  assign RetimeWrapper_4_reset = reset; // @[:@48225.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@48227.4]
  assign RetimeWrapper_4_io_in = io_sigsIn_done; // @[package.scala 94:16:@48226.4]
  assign RetimeWrapper_5_clock = clock; // @[:@48235.4]
  assign RetimeWrapper_5_reset = reset; // @[:@48236.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@48238.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_done; // @[package.scala 94:16:@48237.4]
  assign RetimeWrapper_6_clock = clock; // @[:@48246.4]
  assign RetimeWrapper_6_reset = reset; // @[:@48247.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@48249.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_done; // @[package.scala 94:16:@48248.4]
  assign RetimeWrapper_7_clock = clock; // @[:@48257.4]
  assign RetimeWrapper_7_reset = reset; // @[:@48258.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@48260.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_done; // @[package.scala 94:16:@48259.4]
  assign RetimeWrapper_8_clock = clock; // @[:@48268.4]
  assign RetimeWrapper_8_reset = reset; // @[:@48269.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@48271.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_done; // @[package.scala 94:16:@48270.4]
endmodule
module SRAM_74( // @[:@49103.2]
  input         clock, // @[:@49104.4]
  input         reset, // @[:@49105.4]
  input         io_rPort_0_en_0, // @[:@49106.4]
  output [31:0] io_rPort_0_output_0, // @[:@49106.4]
  input  [31:0] io_wPort_0_data_0, // @[:@49106.4]
  input         io_wPort_0_en_0 // @[:@49106.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@49121.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@49121.4]
  wire  Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@49121.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@49121.4]
  wire  Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@49121.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@49121.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@49121.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@49121.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@49147.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@49147.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@49161.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@49161.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@49161.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@49161.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@49161.4]
  wire [33:0] _T_70; // @[Cat.scala 30:58:@49139.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@49151.4]
  wire [2:0] _T_78; // @[Cat.scala 30:58:@49153.4]
  Mem1D_39 Mem1D ( // @[MemPrimitives.scala 64:21:@49121.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@49147.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@49161.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_70 = {io_wPort_0_en_0,io_wPort_0_data_0,1'h0}; // @[Cat.scala 30:58:@49139.4]
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@49151.4]
  assign _T_78 = {_T_76,1'h1,1'h0}; // @[Cat.scala 30:58:@49153.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@49168.4]
  assign Mem1D_clock = clock; // @[:@49122.4]
  assign Mem1D_reset = reset; // @[:@49123.4]
  assign Mem1D_io_r_ofs_0 = _T_78[0]; // @[MemPrimitives.scala 131:28:@49157.4]
  assign Mem1D_io_r_backpressure = _T_78[1]; // @[MemPrimitives.scala 132:32:@49158.4]
  assign Mem1D_io_w_ofs_0 = _T_70[0]; // @[MemPrimitives.scala 94:28:@49143.4]
  assign Mem1D_io_w_data_0 = _T_70[32:1]; // @[MemPrimitives.scala 95:29:@49144.4]
  assign Mem1D_io_w_en_0 = _T_70[33]; // @[MemPrimitives.scala 96:27:@49145.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@49150.4]
  assign RetimeWrapper_clock = clock; // @[:@49162.4]
  assign RetimeWrapper_reset = reset; // @[:@49163.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@49165.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@49164.4]
endmodule
module x594_force_0( // @[:@49371.2]
  input         clock, // @[:@49372.4]
  input         reset, // @[:@49373.4]
  input         io_rPort_0_en_0, // @[:@49374.4]
  output [31:0] io_rPort_0_output_0, // @[:@49374.4]
  input  [31:0] io_wPort_0_data_0, // @[:@49374.4]
  input         io_wPort_0_en_0, // @[:@49374.4]
  input         io_sEn_0, // @[:@49374.4]
  input         io_sEn_1, // @[:@49374.4]
  input         io_sDone_0, // @[:@49374.4]
  input         io_sDone_1 // @[:@49374.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@49383.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@49383.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@49383.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@49383.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@49383.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@49383.4]
  wire [2:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@49383.4]
  wire [2:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@49383.4]
  wire  SRAM_clock; // @[NBuffers.scala 94:23:@49390.4]
  wire  SRAM_reset; // @[NBuffers.scala 94:23:@49390.4]
  wire  SRAM_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@49390.4]
  wire [31:0] SRAM_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@49390.4]
  wire [31:0] SRAM_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@49390.4]
  wire  SRAM_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@49390.4]
  wire  SRAM_1_clock; // @[NBuffers.scala 94:23:@49406.4]
  wire  SRAM_1_reset; // @[NBuffers.scala 94:23:@49406.4]
  wire  SRAM_1_io_rPort_0_en_0; // @[NBuffers.scala 94:23:@49406.4]
  wire [31:0] SRAM_1_io_rPort_0_output_0; // @[NBuffers.scala 94:23:@49406.4]
  wire [31:0] SRAM_1_io_wPort_0_data_0; // @[NBuffers.scala 94:23:@49406.4]
  wire  SRAM_1_io_wPort_0_en_0; // @[NBuffers.scala 94:23:@49406.4]
  wire  _T_110; // @[NBuffers.scala 104:105:@49422.4]
  wire  _T_114; // @[NBuffers.scala 108:92:@49432.4]
  wire  _T_117; // @[NBuffers.scala 104:105:@49438.4]
  wire  _T_121; // @[NBuffers.scala 108:92:@49448.4]
  wire [31:0] _T_129; // @[Mux.scala 19:72:@49456.4]
  wire [31:0] _T_131; // @[Mux.scala 19:72:@49457.4]
  NBufController ctrl ( // @[NBuffers.scala 83:20:@49383.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1)
  );
  SRAM_74 SRAM ( // @[NBuffers.scala 94:23:@49390.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_rPort_0_en_0(SRAM_io_rPort_0_en_0),
    .io_rPort_0_output_0(SRAM_io_rPort_0_output_0),
    .io_wPort_0_data_0(SRAM_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_io_wPort_0_en_0)
  );
  SRAM_74 SRAM_1 ( // @[NBuffers.scala 94:23:@49406.4]
    .clock(SRAM_1_clock),
    .reset(SRAM_1_reset),
    .io_rPort_0_en_0(SRAM_1_io_rPort_0_en_0),
    .io_rPort_0_output_0(SRAM_1_io_rPort_0_output_0),
    .io_wPort_0_data_0(SRAM_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(SRAM_1_io_wPort_0_en_0)
  );
  assign _T_110 = ctrl_io_statesInW_0 == 3'h0; // @[NBuffers.scala 104:105:@49422.4]
  assign _T_114 = ctrl_io_statesInR_1 == 3'h0; // @[NBuffers.scala 108:92:@49432.4]
  assign _T_117 = ctrl_io_statesInW_0 == 3'h1; // @[NBuffers.scala 104:105:@49438.4]
  assign _T_121 = ctrl_io_statesInR_1 == 3'h1; // @[NBuffers.scala 108:92:@49448.4]
  assign _T_129 = _T_114 ? SRAM_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@49456.4]
  assign _T_131 = _T_121 ? SRAM_1_io_rPort_0_output_0 : 32'h0; // @[Mux.scala 19:72:@49457.4]
  assign io_rPort_0_output_0 = _T_129 | _T_131; // @[NBuffers.scala 115:66:@49461.4]
  assign ctrl_clock = clock; // @[:@49384.4]
  assign ctrl_reset = reset; // @[:@49385.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@49386.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@49388.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@49387.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@49389.4]
  assign SRAM_clock = clock; // @[:@49391.4]
  assign SRAM_reset = reset; // @[:@49392.4]
  assign SRAM_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_114; // @[MemPrimitives.scala 43:33:@49436.4]
  assign SRAM_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@49425.4]
  assign SRAM_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_110; // @[MemPrimitives.scala 37:29:@49431.4]
  assign SRAM_1_clock = clock; // @[:@49407.4]
  assign SRAM_1_reset = reset; // @[:@49408.4]
  assign SRAM_1_io_rPort_0_en_0 = io_rPort_0_en_0 & _T_121; // @[MemPrimitives.scala 43:33:@49452.4]
  assign SRAM_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@49441.4]
  assign SRAM_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_117; // @[MemPrimitives.scala 37:29:@49447.4]
endmodule
module FF_28( // @[:@50154.2]
  input   clock, // @[:@50155.4]
  input   reset, // @[:@50156.4]
  output  io_rPort_1_output_0, // @[:@50157.4]
  output  io_rPort_0_output_0, // @[:@50157.4]
  input   io_wPort_0_data_0, // @[:@50157.4]
  input   io_wPort_0_reset, // @[:@50157.4]
  input   io_wPort_0_en_0 // @[:@50157.4]
);
  reg  ff; // @[MemPrimitives.scala 321:19:@50177.4]
  reg [31:0] _RAND_0;
  wire  _T_94; // @[MemPrimitives.scala 325:32:@50179.4]
  wire  _T_95; // @[MemPrimitives.scala 325:12:@50180.4]
  assign _T_94 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@50179.4]
  assign _T_95 = io_wPort_0_reset ? 1'h0 : _T_94; // @[MemPrimitives.scala 325:12:@50180.4]
  assign io_rPort_1_output_0 = ff; // @[MemPrimitives.scala 326:34:@50183.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@50182.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 1'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 1'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module x595_reg( // @[:@50216.2]
  input   clock, // @[:@50217.4]
  input   reset, // @[:@50218.4]
  output  io_rPort_1_output_0, // @[:@50219.4]
  output  io_rPort_0_output_0, // @[:@50219.4]
  input   io_wPort_0_data_0, // @[:@50219.4]
  input   io_wPort_0_reset, // @[:@50219.4]
  input   io_wPort_0_en_0, // @[:@50219.4]
  input   io_sEn_0, // @[:@50219.4]
  input   io_sEn_1, // @[:@50219.4]
  input   io_sDone_0, // @[:@50219.4]
  input   io_sDone_1 // @[:@50219.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@50229.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@50229.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@50229.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@50229.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@50229.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@50229.4]
  wire [2:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@50229.4]
  wire [2:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@50229.4]
  wire  FF_clock; // @[NBuffers.scala 146:23:@50236.4]
  wire  FF_reset; // @[NBuffers.scala 146:23:@50236.4]
  wire  FF_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@50236.4]
  wire  FF_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@50236.4]
  wire  FF_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@50236.4]
  wire  FF_io_wPort_0_reset; // @[NBuffers.scala 146:23:@50236.4]
  wire  FF_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@50236.4]
  wire  FF_1_clock; // @[NBuffers.scala 146:23:@50257.4]
  wire  FF_1_reset; // @[NBuffers.scala 146:23:@50257.4]
  wire  FF_1_io_rPort_1_output_0; // @[NBuffers.scala 146:23:@50257.4]
  wire  FF_1_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@50257.4]
  wire  FF_1_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@50257.4]
  wire  FF_1_io_wPort_0_reset; // @[NBuffers.scala 146:23:@50257.4]
  wire  FF_1_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@50257.4]
  wire  _T_140; // @[NBuffers.scala 153:105:@50280.4]
  wire  _T_144; // @[NBuffers.scala 157:92:@50290.4]
  wire  _T_150; // @[NBuffers.scala 153:105:@50302.4]
  wire  _T_154; // @[NBuffers.scala 157:92:@50312.4]
  wire  _T_165; // @[Mux.scala 19:72:@50326.4]
  wire  _T_167; // @[Mux.scala 19:72:@50327.4]
  wire  _T_177; // @[Mux.scala 19:72:@50334.4]
  wire  _T_179; // @[Mux.scala 19:72:@50335.4]
  NBufController ctrl ( // @[NBuffers.scala 83:20:@50229.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1)
  );
  FF_28 FF ( // @[NBuffers.scala 146:23:@50236.4]
    .clock(FF_clock),
    .reset(FF_reset),
    .io_rPort_1_output_0(FF_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_io_wPort_0_en_0)
  );
  FF_28 FF_1 ( // @[NBuffers.scala 146:23:@50257.4]
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_rPort_1_output_0(FF_1_io_rPort_1_output_0),
    .io_rPort_0_output_0(FF_1_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_1_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_1_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_1_io_wPort_0_en_0)
  );
  assign _T_140 = ctrl_io_statesInW_0 == 3'h0; // @[NBuffers.scala 153:105:@50280.4]
  assign _T_144 = ctrl_io_statesInR_1 == 3'h0; // @[NBuffers.scala 157:92:@50290.4]
  assign _T_150 = ctrl_io_statesInW_0 == 3'h1; // @[NBuffers.scala 153:105:@50302.4]
  assign _T_154 = ctrl_io_statesInR_1 == 3'h1; // @[NBuffers.scala 157:92:@50312.4]
  assign _T_165 = _T_144 ? FF_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@50326.4]
  assign _T_167 = _T_154 ? FF_1_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@50327.4]
  assign _T_177 = _T_144 ? FF_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@50334.4]
  assign _T_179 = _T_154 ? FF_1_io_rPort_1_output_0 : 1'h0; // @[Mux.scala 19:72:@50335.4]
  assign io_rPort_1_output_0 = _T_177 | _T_179; // @[NBuffers.scala 163:66:@50339.4]
  assign io_rPort_0_output_0 = _T_165 | _T_167; // @[NBuffers.scala 163:66:@50331.4]
  assign ctrl_clock = clock; // @[:@50230.4]
  assign ctrl_reset = reset; // @[:@50231.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@50232.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@50234.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@50233.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@50235.4]
  assign FF_clock = clock; // @[:@50237.4]
  assign FF_reset = reset; // @[:@50238.4]
  assign FF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@50283.4]
  assign FF_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@50284.4]
  assign FF_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_140; // @[MemPrimitives.scala 37:29:@50289.4]
  assign FF_1_clock = clock; // @[:@50258.4]
  assign FF_1_reset = reset; // @[:@50259.4]
  assign FF_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@50305.4]
  assign FF_1_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@50306.4]
  assign FF_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_150; // @[MemPrimitives.scala 37:29:@50311.4]
endmodule
module FF_30( // @[:@51032.2]
  input   clock, // @[:@51033.4]
  input   reset, // @[:@51034.4]
  output  io_rPort_0_output_0, // @[:@51035.4]
  input   io_wPort_0_data_0, // @[:@51035.4]
  input   io_wPort_0_reset, // @[:@51035.4]
  input   io_wPort_0_en_0 // @[:@51035.4]
);
  reg  ff; // @[MemPrimitives.scala 321:19:@51050.4]
  reg [31:0] _RAND_0;
  wire  _T_68; // @[MemPrimitives.scala 325:32:@51052.4]
  wire  _T_69; // @[MemPrimitives.scala 325:12:@51053.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@51052.4]
  assign _T_69 = io_wPort_0_reset ? 1'h0 : _T_68; // @[MemPrimitives.scala 325:12:@51053.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@51055.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 1'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 1'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module x596_reg( // @[:@51082.2]
  input   clock, // @[:@51083.4]
  input   reset, // @[:@51084.4]
  output  io_rPort_0_output_0, // @[:@51085.4]
  input   io_wPort_0_data_0, // @[:@51085.4]
  input   io_wPort_0_reset, // @[:@51085.4]
  input   io_wPort_0_en_0, // @[:@51085.4]
  input   io_sEn_0, // @[:@51085.4]
  input   io_sEn_1, // @[:@51085.4]
  input   io_sDone_0, // @[:@51085.4]
  input   io_sDone_1 // @[:@51085.4]
);
  wire  ctrl_clock; // @[NBuffers.scala 83:20:@51094.4]
  wire  ctrl_reset; // @[NBuffers.scala 83:20:@51094.4]
  wire  ctrl_io_sEn_0; // @[NBuffers.scala 83:20:@51094.4]
  wire  ctrl_io_sEn_1; // @[NBuffers.scala 83:20:@51094.4]
  wire  ctrl_io_sDone_0; // @[NBuffers.scala 83:20:@51094.4]
  wire  ctrl_io_sDone_1; // @[NBuffers.scala 83:20:@51094.4]
  wire [2:0] ctrl_io_statesInW_0; // @[NBuffers.scala 83:20:@51094.4]
  wire [2:0] ctrl_io_statesInR_1; // @[NBuffers.scala 83:20:@51094.4]
  wire  FF_clock; // @[NBuffers.scala 146:23:@51101.4]
  wire  FF_reset; // @[NBuffers.scala 146:23:@51101.4]
  wire  FF_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@51101.4]
  wire  FF_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@51101.4]
  wire  FF_io_wPort_0_reset; // @[NBuffers.scala 146:23:@51101.4]
  wire  FF_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@51101.4]
  wire  FF_1_clock; // @[NBuffers.scala 146:23:@51117.4]
  wire  FF_1_reset; // @[NBuffers.scala 146:23:@51117.4]
  wire  FF_1_io_rPort_0_output_0; // @[NBuffers.scala 146:23:@51117.4]
  wire  FF_1_io_wPort_0_data_0; // @[NBuffers.scala 146:23:@51117.4]
  wire  FF_1_io_wPort_0_reset; // @[NBuffers.scala 146:23:@51117.4]
  wire  FF_1_io_wPort_0_en_0; // @[NBuffers.scala 146:23:@51117.4]
  wire  _T_110; // @[NBuffers.scala 153:105:@51135.4]
  wire  _T_114; // @[NBuffers.scala 157:92:@51145.4]
  wire  _T_117; // @[NBuffers.scala 153:105:@51151.4]
  wire  _T_121; // @[NBuffers.scala 157:92:@51161.4]
  wire  _T_129; // @[Mux.scala 19:72:@51169.4]
  wire  _T_131; // @[Mux.scala 19:72:@51170.4]
  NBufController ctrl ( // @[NBuffers.scala 83:20:@51094.4]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_sEn_0(ctrl_io_sEn_0),
    .io_sEn_1(ctrl_io_sEn_1),
    .io_sDone_0(ctrl_io_sDone_0),
    .io_sDone_1(ctrl_io_sDone_1),
    .io_statesInW_0(ctrl_io_statesInW_0),
    .io_statesInR_1(ctrl_io_statesInR_1)
  );
  FF_30 FF ( // @[NBuffers.scala 146:23:@51101.4]
    .clock(FF_clock),
    .reset(FF_reset),
    .io_rPort_0_output_0(FF_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_io_wPort_0_en_0)
  );
  FF_30 FF_1 ( // @[NBuffers.scala 146:23:@51117.4]
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_rPort_0_output_0(FF_1_io_rPort_0_output_0),
    .io_wPort_0_data_0(FF_1_io_wPort_0_data_0),
    .io_wPort_0_reset(FF_1_io_wPort_0_reset),
    .io_wPort_0_en_0(FF_1_io_wPort_0_en_0)
  );
  assign _T_110 = ctrl_io_statesInW_0 == 3'h0; // @[NBuffers.scala 153:105:@51135.4]
  assign _T_114 = ctrl_io_statesInR_1 == 3'h0; // @[NBuffers.scala 157:92:@51145.4]
  assign _T_117 = ctrl_io_statesInW_0 == 3'h1; // @[NBuffers.scala 153:105:@51151.4]
  assign _T_121 = ctrl_io_statesInR_1 == 3'h1; // @[NBuffers.scala 157:92:@51161.4]
  assign _T_129 = _T_114 ? FF_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@51169.4]
  assign _T_131 = _T_121 ? FF_1_io_rPort_0_output_0 : 1'h0; // @[Mux.scala 19:72:@51170.4]
  assign io_rPort_0_output_0 = _T_129 | _T_131; // @[NBuffers.scala 163:66:@51174.4]
  assign ctrl_clock = clock; // @[:@51095.4]
  assign ctrl_reset = reset; // @[:@51096.4]
  assign ctrl_io_sEn_0 = io_sEn_0; // @[NBuffers.scala 85:20:@51097.4]
  assign ctrl_io_sEn_1 = io_sEn_1; // @[NBuffers.scala 85:20:@51099.4]
  assign ctrl_io_sDone_0 = io_sDone_0; // @[NBuffers.scala 86:22:@51098.4]
  assign ctrl_io_sDone_1 = io_sDone_1; // @[NBuffers.scala 86:22:@51100.4]
  assign FF_clock = clock; // @[:@51102.4]
  assign FF_reset = reset; // @[:@51103.4]
  assign FF_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@51138.4]
  assign FF_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@51139.4]
  assign FF_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_110; // @[MemPrimitives.scala 37:29:@51144.4]
  assign FF_1_clock = clock; // @[:@51118.4]
  assign FF_1_reset = reset; // @[:@51119.4]
  assign FF_1_io_wPort_0_data_0 = io_wPort_0_data_0; // @[MemPrimitives.scala 33:29:@51154.4]
  assign FF_1_io_wPort_0_reset = io_wPort_0_reset; // @[MemPrimitives.scala 34:29:@51155.4]
  assign FF_1_io_wPort_0_en_0 = io_wPort_0_en_0 & _T_117; // @[MemPrimitives.scala 37:29:@51160.4]
endmodule
module x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1( // @[:@51931.2]
  input         clock, // @[:@51932.4]
  input         reset, // @[:@51933.4]
  output        io_in_x555_tmp_1_sEn_2, // @[:@51934.4]
  output        io_in_x555_tmp_1_sDone_2, // @[:@51934.4]
  output        io_in_x554_tmp_0_sEn_2, // @[:@51934.4]
  output        io_in_x554_tmp_0_sDone_2, // @[:@51934.4]
  output        io_in_x558_tmp_4_sEn_2, // @[:@51934.4]
  output        io_in_x558_tmp_4_sDone_2, // @[:@51934.4]
  output        io_in_x557_tmp_3_sEn_2, // @[:@51934.4]
  output        io_in_x557_tmp_3_sDone_2, // @[:@51934.4]
  output        io_in_x580_r_0_rPort_0_en_0, // @[:@51934.4]
  input  [31:0] io_in_x580_r_0_rPort_0_output_0, // @[:@51934.4]
  output        io_in_x580_r_0_sEn_1, // @[:@51934.4]
  output        io_in_x580_r_0_sDone_1, // @[:@51934.4]
  output        io_in_x595_reg_wPort_0_data_0, // @[:@51934.4]
  output        io_in_x595_reg_wPort_0_reset, // @[:@51934.4]
  output        io_in_x595_reg_wPort_0_en_0, // @[:@51934.4]
  output        io_in_x595_reg_reset, // @[:@51934.4]
  output        io_in_x595_reg_sEn_0, // @[:@51934.4]
  output        io_in_x595_reg_sDone_0, // @[:@51934.4]
  output        io_in_x556_tmp_2_sEn_2, // @[:@51934.4]
  output        io_in_x556_tmp_2_sDone_2, // @[:@51934.4]
  output        io_in_x596_reg_wPort_0_data_0, // @[:@51934.4]
  output        io_in_x596_reg_wPort_0_reset, // @[:@51934.4]
  output        io_in_x596_reg_wPort_0_en_0, // @[:@51934.4]
  output        io_in_x596_reg_reset, // @[:@51934.4]
  output        io_in_x596_reg_sEn_0, // @[:@51934.4]
  output        io_in_x596_reg_sDone_0, // @[:@51934.4]
  input         io_sigsIn_done, // @[:@51934.4]
  input         io_sigsIn_datapathEn, // @[:@51934.4]
  input         io_sigsIn_baseEn, // @[:@51934.4]
  input         io_sigsIn_break, // @[:@51934.4]
  input         io_rr // @[:@51934.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@52301.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@52301.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@52301.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@52301.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@52301.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@52321.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@52321.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@52321.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@52321.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@52321.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@52338.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@52338.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@52338.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@52338.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@52338.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@52349.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@52349.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@52349.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@52349.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@52349.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@52360.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@52360.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@52360.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@52360.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@52360.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@52371.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@52371.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@52371.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@52371.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@52371.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@52382.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@52382.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@52382.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@52382.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@52382.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@52393.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@52393.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@52393.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@52393.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@52393.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@52404.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@52404.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@52404.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@52404.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@52404.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@52415.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@52415.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@52415.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@52415.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@52415.4]
  wire  _T_2319; // @[sm_x605_inr_UnitPipe.scala 97:114:@52262.4]
  wire  _T_2320; // @[sm_x605_inr_UnitPipe.scala 97:111:@52263.4]
  wire  _T_2325; // @[implicits.scala 56:10:@52266.4]
  wire [31:0] _T_2337; // @[Math.scala 476:50:@52281.4]
  wire  x599; // @[Math.scala 476:44:@52282.4]
  wire  x600; // @[Math.scala 476:44:@52289.4]
  wire  x601; // @[sm_x605_inr_UnitPipe.scala 107:20:@52292.4]
  wire  _T_2358; // @[package.scala 96:25:@52306.4 package.scala 96:25:@52307.4]
  wire  _T_2360; // @[implicits.scala 56:10:@52308.4]
  wire  _T_2361; // @[sm_x605_inr_UnitPipe.scala 114:133:@52309.4]
  wire  _T_2373; // @[package.scala 96:25:@52326.4 package.scala 96:25:@52327.4]
  wire  _T_2375; // @[implicits.scala 56:10:@52328.4]
  wire  _T_2376; // @[sm_x605_inr_UnitPipe.scala 119:133:@52329.4]
  wire  _T_2385; // @[package.scala 96:25:@52343.4 package.scala 96:25:@52344.4]
  wire  _T_2391; // @[package.scala 96:25:@52354.4 package.scala 96:25:@52355.4]
  wire  _T_2397; // @[package.scala 96:25:@52365.4 package.scala 96:25:@52366.4]
  wire  _T_2403; // @[package.scala 96:25:@52376.4 package.scala 96:25:@52377.4]
  wire  _T_2409; // @[package.scala 96:25:@52387.4 package.scala 96:25:@52388.4]
  wire  _T_2415; // @[package.scala 96:25:@52398.4 package.scala 96:25:@52399.4]
  wire  _T_2421; // @[package.scala 96:25:@52409.4 package.scala 96:25:@52410.4]
  wire  _T_2427; // @[package.scala 96:25:@52420.4 package.scala 96:25:@52421.4]
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@52301.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@52321.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@52338.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@52349.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@52360.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@52371.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@52382.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@52393.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@52404.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@52415.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  assign _T_2319 = ~ io_sigsIn_break; // @[sm_x605_inr_UnitPipe.scala 97:114:@52262.4]
  assign _T_2320 = io_rr & _T_2319; // @[sm_x605_inr_UnitPipe.scala 97:111:@52263.4]
  assign _T_2325 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 56:10:@52266.4]
  assign _T_2337 = $signed(io_in_x580_r_0_rPort_0_output_0); // @[Math.scala 476:50:@52281.4]
  assign x599 = $signed(32'sh0) < $signed(_T_2337); // @[Math.scala 476:44:@52282.4]
  assign x600 = $signed(32'sh400000) < $signed(_T_2337); // @[Math.scala 476:44:@52289.4]
  assign x601 = x599 & x600; // @[sm_x605_inr_UnitPipe.scala 107:20:@52292.4]
  assign _T_2358 = RetimeWrapper_io_out; // @[package.scala 96:25:@52306.4 package.scala 96:25:@52307.4]
  assign _T_2360 = io_rr ? _T_2358 : 1'h0; // @[implicits.scala 56:10:@52308.4]
  assign _T_2361 = _T_2319 & _T_2360; // @[sm_x605_inr_UnitPipe.scala 114:133:@52309.4]
  assign _T_2373 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@52326.4 package.scala 96:25:@52327.4]
  assign _T_2375 = io_rr ? _T_2373 : 1'h0; // @[implicits.scala 56:10:@52328.4]
  assign _T_2376 = _T_2319 & _T_2375; // @[sm_x605_inr_UnitPipe.scala 119:133:@52329.4]
  assign _T_2385 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@52343.4 package.scala 96:25:@52344.4]
  assign _T_2391 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@52354.4 package.scala 96:25:@52355.4]
  assign _T_2397 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@52365.4 package.scala 96:25:@52366.4]
  assign _T_2403 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@52376.4 package.scala 96:25:@52377.4]
  assign _T_2409 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@52387.4 package.scala 96:25:@52388.4]
  assign _T_2415 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@52398.4 package.scala 96:25:@52399.4]
  assign _T_2421 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@52409.4 package.scala 96:25:@52410.4]
  assign _T_2427 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@52420.4 package.scala 96:25:@52421.4]
  assign io_in_x555_tmp_1_sEn_2 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@52357.4]
  assign io_in_x555_tmp_1_sDone_2 = io_rr ? _T_2391 : 1'h0; // @[MemInterfaceType.scala 197:17:@52358.4]
  assign io_in_x554_tmp_0_sEn_2 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@52346.4]
  assign io_in_x554_tmp_0_sDone_2 = io_rr ? _T_2385 : 1'h0; // @[MemInterfaceType.scala 197:17:@52347.4]
  assign io_in_x558_tmp_4_sEn_2 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@52390.4]
  assign io_in_x558_tmp_4_sDone_2 = io_rr ? _T_2409 : 1'h0; // @[MemInterfaceType.scala 197:17:@52391.4]
  assign io_in_x557_tmp_3_sEn_2 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@52379.4]
  assign io_in_x557_tmp_3_sDone_2 = io_rr ? _T_2403 : 1'h0; // @[MemInterfaceType.scala 197:17:@52380.4]
  assign io_in_x580_r_0_rPort_0_en_0 = _T_2320 & _T_2325; // @[MemInterfaceType.scala 110:79:@52273.4]
  assign io_in_x580_r_0_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@52401.4]
  assign io_in_x580_r_0_sDone_1 = io_rr ? _T_2415 : 1'h0; // @[MemInterfaceType.scala 197:17:@52402.4]
  assign io_in_x595_reg_wPort_0_data_0 = x599 & x600; // @[MemInterfaceType.scala 90:56:@52314.4]
  assign io_in_x595_reg_wPort_0_reset = io_in_x595_reg_reset; // @[MemInterfaceType.scala 91:23:@52315.4]
  assign io_in_x595_reg_wPort_0_en_0 = _T_2361 & _T_2319; // @[MemInterfaceType.scala 93:57:@52316.4]
  assign io_in_x595_reg_reset = 1'h0;
  assign io_in_x595_reg_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@52412.4]
  assign io_in_x595_reg_sDone_0 = io_rr ? _T_2421 : 1'h0; // @[MemInterfaceType.scala 197:17:@52413.4]
  assign io_in_x556_tmp_2_sEn_2 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@52368.4]
  assign io_in_x556_tmp_2_sDone_2 = io_rr ? _T_2397 : 1'h0; // @[MemInterfaceType.scala 197:17:@52369.4]
  assign io_in_x596_reg_wPort_0_data_0 = ~ x601; // @[MemInterfaceType.scala 90:56:@52334.4]
  assign io_in_x596_reg_wPort_0_reset = io_in_x596_reg_reset; // @[MemInterfaceType.scala 91:23:@52335.4]
  assign io_in_x596_reg_wPort_0_en_0 = _T_2376 & _T_2319; // @[MemInterfaceType.scala 93:57:@52336.4]
  assign io_in_x596_reg_reset = 1'h0;
  assign io_in_x596_reg_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@52423.4]
  assign io_in_x596_reg_sDone_0 = io_rr ? _T_2427 : 1'h0; // @[MemInterfaceType.scala 197:17:@52424.4]
  assign RetimeWrapper_clock = clock; // @[:@52302.4]
  assign RetimeWrapper_reset = reset; // @[:@52303.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@52305.4]
  assign RetimeWrapper_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@52304.4]
  assign RetimeWrapper_1_clock = clock; // @[:@52322.4]
  assign RetimeWrapper_1_reset = reset; // @[:@52323.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@52325.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@52324.4]
  assign RetimeWrapper_2_clock = clock; // @[:@52339.4]
  assign RetimeWrapper_2_reset = reset; // @[:@52340.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@52342.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_done; // @[package.scala 94:16:@52341.4]
  assign RetimeWrapper_3_clock = clock; // @[:@52350.4]
  assign RetimeWrapper_3_reset = reset; // @[:@52351.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@52353.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_done; // @[package.scala 94:16:@52352.4]
  assign RetimeWrapper_4_clock = clock; // @[:@52361.4]
  assign RetimeWrapper_4_reset = reset; // @[:@52362.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@52364.4]
  assign RetimeWrapper_4_io_in = io_sigsIn_done; // @[package.scala 94:16:@52363.4]
  assign RetimeWrapper_5_clock = clock; // @[:@52372.4]
  assign RetimeWrapper_5_reset = reset; // @[:@52373.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@52375.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_done; // @[package.scala 94:16:@52374.4]
  assign RetimeWrapper_6_clock = clock; // @[:@52383.4]
  assign RetimeWrapper_6_reset = reset; // @[:@52384.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@52386.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_done; // @[package.scala 94:16:@52385.4]
  assign RetimeWrapper_7_clock = clock; // @[:@52394.4]
  assign RetimeWrapper_7_reset = reset; // @[:@52395.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@52397.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_done; // @[package.scala 94:16:@52396.4]
  assign RetimeWrapper_8_clock = clock; // @[:@52405.4]
  assign RetimeWrapper_8_reset = reset; // @[:@52406.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@52408.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_done; // @[package.scala 94:16:@52407.4]
  assign RetimeWrapper_9_clock = clock; // @[:@52416.4]
  assign RetimeWrapper_9_reset = reset; // @[:@52417.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@52419.4]
  assign RetimeWrapper_9_io_in = io_sigsIn_done; // @[package.scala 94:16:@52418.4]
endmodule
module x621_inr_Switch_sm( // @[:@52580.2]
  input   clock, // @[:@52581.4]
  input   reset, // @[:@52582.4]
  input   io_enable, // @[:@52583.4]
  output  io_done, // @[:@52583.4]
  input   io_parentAck, // @[:@52583.4]
  input   io_backpressure, // @[:@52583.4]
  input   io_doneIn_0, // @[:@52583.4]
  input   io_doneIn_1, // @[:@52583.4]
  output  io_childAck_0, // @[:@52583.4]
  output  io_childAck_1, // @[:@52583.4]
  input   io_selectsIn_0, // @[:@52583.4]
  input   io_selectsIn_1, // @[:@52583.4]
  output  io_selectsOut_0, // @[:@52583.4]
  output  io_selectsOut_1 // @[:@52583.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@52585.4]
  wire  active_reset; // @[Controllers.scala 261:22:@52585.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@52585.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@52585.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@52585.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@52585.4]
  wire  done_clock; // @[Controllers.scala 262:20:@52588.4]
  wire  done_reset; // @[Controllers.scala 262:20:@52588.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@52588.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@52588.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@52588.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@52588.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@52641.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@52641.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@52641.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@52641.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@52641.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@52649.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@52649.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@52649.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@52649.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@52649.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@52659.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@52659.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@52659.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@52659.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@52659.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@52667.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@52667.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@52667.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@52667.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@52667.4]
  wire  _T_82; // @[Controllers.scala 264:62:@52595.4]
  wire  _T_103; // @[package.scala 100:49:@52621.4]
  reg  _T_120; // @[package.scala 48:56:@52637.4]
  reg [31:0] _RAND_0;
  wire  _T_125; // @[package.scala 96:25:@52646.4 package.scala 96:25:@52647.4]
  wire  _T_131; // @[package.scala 96:25:@52654.4 package.scala 96:25:@52655.4]
  wire  _T_138; // @[package.scala 96:25:@52664.4 package.scala 96:25:@52665.4]
  wire  _T_144; // @[package.scala 96:25:@52672.4 package.scala 96:25:@52673.4]
  SRFF active ( // @[Controllers.scala 261:22:@52585.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@52588.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@52641.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@52649.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@52659.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@52667.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@52595.4]
  assign _T_103 = done_io_output == 1'h0; // @[package.scala 100:49:@52621.4]
  assign _T_125 = RetimeWrapper_io_out; // @[package.scala 96:25:@52646.4 package.scala 96:25:@52647.4]
  assign _T_131 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@52654.4 package.scala 96:25:@52655.4]
  assign _T_138 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@52664.4 package.scala 96:25:@52665.4]
  assign _T_144 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@52672.4 package.scala 96:25:@52673.4]
  assign io_done = done_io_output & _T_120; // @[Controllers.scala 287:13:@52640.4]
  assign io_childAck_0 = _T_125 | _T_131; // @[Controllers.scala 288:56:@52658.4]
  assign io_childAck_1 = _T_138 | _T_144; // @[Controllers.scala 288:56:@52676.4]
  assign io_selectsOut_0 = io_selectsIn_0 & io_enable; // @[Controllers.scala 271:55:@52616.4]
  assign io_selectsOut_1 = io_selectsIn_1 & io_enable; // @[Controllers.scala 271:55:@52618.4]
  assign active_clock = clock; // @[:@52586.4]
  assign active_reset = reset; // @[:@52587.4]
  assign active_io_input_set = io_enable & _T_82; // @[Controllers.scala 264:23:@52598.4]
  assign active_io_input_reset = io_parentAck; // @[Controllers.scala 265:25:@52602.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@52603.4]
  assign done_clock = clock; // @[:@52589.4]
  assign done_reset = reset; // @[:@52590.4]
  assign done_io_input_set = io_doneIn_0 | io_doneIn_1; // @[Controllers.scala 269:50:@52614.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@52611.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@52612.4]
  assign RetimeWrapper_clock = clock; // @[:@52642.4]
  assign RetimeWrapper_reset = reset; // @[:@52643.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@52645.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@52644.4]
  assign RetimeWrapper_1_clock = clock; // @[:@52650.4]
  assign RetimeWrapper_1_reset = reset; // @[:@52651.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@52653.4]
  assign RetimeWrapper_1_io_in = 1'h0; // @[package.scala 94:16:@52652.4]
  assign RetimeWrapper_2_clock = clock; // @[:@52660.4]
  assign RetimeWrapper_2_reset = reset; // @[:@52661.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@52663.4]
  assign RetimeWrapper_2_io_in = io_doneIn_1; // @[package.scala 94:16:@52662.4]
  assign RetimeWrapper_3_clock = clock; // @[:@52668.4]
  assign RetimeWrapper_3_reset = reset; // @[:@52669.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@52671.4]
  assign RetimeWrapper_3_io_in = 1'h0; // @[package.scala 94:16:@52670.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_120 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_120 <= 1'h0;
    end else begin
      _T_120 <= _T_103;
    end
  end
endmodule
module RetimeWrapper_608( // @[:@52863.2]
  input   clock, // @[:@52864.4]
  input   reset, // @[:@52865.4]
  input   io_flow, // @[:@52866.4]
  input   io_in, // @[:@52866.4]
  output  io_out // @[:@52866.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@52868.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@52868.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@52868.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@52868.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@52868.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@52868.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(103)) sr ( // @[RetimeShiftRegister.scala 15:20:@52868.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@52881.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@52880.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@52879.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@52878.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@52877.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@52875.4]
endmodule
module RetimeWrapper_612( // @[:@52991.2]
  input   clock, // @[:@52992.4]
  input   reset, // @[:@52993.4]
  input   io_flow, // @[:@52994.4]
  input   io_in // @[:@52994.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@52996.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@52996.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@52996.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@52996.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@52996.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@52996.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(102)) sr ( // @[RetimeShiftRegister.scala 15:20:@52996.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@53008.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@53007.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@53006.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@53005.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@53003.4]
endmodule
module x619_inr_SwitchCase_sm( // @[:@53011.2]
  input   clock, // @[:@53012.4]
  input   reset, // @[:@53013.4]
  input   io_enable, // @[:@53014.4]
  output  io_done, // @[:@53014.4]
  input   io_ctrDone, // @[:@53014.4]
  output  io_datapathEn, // @[:@53014.4]
  output  io_ctrInc, // @[:@53014.4]
  input   io_parentAck, // @[:@53014.4]
  input   io_break // @[:@53014.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@53016.4]
  wire  active_reset; // @[Controllers.scala 261:22:@53016.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@53016.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@53016.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@53016.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@53016.4]
  wire  done_clock; // @[Controllers.scala 262:20:@53019.4]
  wire  done_reset; // @[Controllers.scala 262:20:@53019.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@53019.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@53019.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@53019.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@53019.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@53053.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@53053.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@53053.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@53053.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@53053.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@53075.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@53075.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@53075.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@53075.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@53075.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@53087.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@53087.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@53087.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@53087.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@53087.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@53095.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@53095.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@53095.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@53095.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@53095.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@53111.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@53111.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@53111.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@53111.4]
  wire  _T_80; // @[Controllers.scala 264:48:@53024.4]
  wire  _T_81; // @[Controllers.scala 264:46:@53025.4]
  wire  _T_82; // @[Controllers.scala 264:62:@53026.4]
  wire  _T_100; // @[package.scala 100:49:@53044.4]
  reg  _T_103; // @[package.scala 48:56:@53045.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@53068.4]
  wire  _T_124; // @[package.scala 96:25:@53080.4 package.scala 96:25:@53081.4]
  wire  _T_126; // @[package.scala 100:49:@53082.4]
  reg  _T_129; // @[package.scala 48:56:@53083.4]
  reg [31:0] _RAND_1;
  wire  _T_150; // @[package.scala 100:49:@53107.4]
  reg  _T_153; // @[package.scala 48:56:@53108.4]
  reg [31:0] _RAND_2;
  SRFF active ( // @[Controllers.scala 261:22:@53016.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@53019.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_608 RetimeWrapper ( // @[package.scala 93:22:@53053.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_608 RetimeWrapper_1 ( // @[package.scala 93:22:@53075.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@53087.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@53095.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_612 RetimeWrapper_4 ( // @[package.scala 93:22:@53111.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@53024.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@53025.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@53026.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@53044.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@53068.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@53080.4 package.scala 96:25:@53081.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@53082.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@53107.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@53086.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@53071.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@53074.4]
  assign active_clock = clock; // @[:@53017.4]
  assign active_reset = reset; // @[:@53018.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@53029.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@53033.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@53034.4]
  assign done_clock = clock; // @[:@53020.4]
  assign done_reset = reset; // @[:@53021.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@53049.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@53042.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@53043.4]
  assign RetimeWrapper_clock = clock; // @[:@53054.4]
  assign RetimeWrapper_reset = reset; // @[:@53055.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@53057.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@53056.4]
  assign RetimeWrapper_1_clock = clock; // @[:@53076.4]
  assign RetimeWrapper_1_reset = reset; // @[:@53077.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@53079.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@53078.4]
  assign RetimeWrapper_2_clock = clock; // @[:@53088.4]
  assign RetimeWrapper_2_reset = reset; // @[:@53089.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@53091.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@53090.4]
  assign RetimeWrapper_3_clock = clock; // @[:@53096.4]
  assign RetimeWrapper_3_reset = reset; // @[:@53097.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@53099.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@53098.4]
  assign RetimeWrapper_4_clock = clock; // @[:@53112.4]
  assign RetimeWrapper_4_reset = reset; // @[:@53113.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@53115.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@53114.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_153 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox_64( // @[:@53132.2]
  input  [31:0] io_a, // @[:@53135.4]
  output [54:0] io_b // @[:@53135.4]
);
  wire [21:0] _T_18; // @[Converter.scala 48:44:@53143.4]
  wire [44:0] tmp_frac; // @[Cat.scala 30:58:@53144.4]
  wire [9:0] new_dec; // @[Converter.scala 88:34:@53147.4]
  assign _T_18 = io_a[21:0]; // @[Converter.scala 48:44:@53143.4]
  assign tmp_frac = {_T_18,23'h0}; // @[Cat.scala 30:58:@53144.4]
  assign new_dec = io_a[31:22]; // @[Converter.scala 88:34:@53147.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@53150.4]
endmodule
module cast_x611_div( // @[:@53152.2]
  input  [31:0] io_b, // @[:@53155.4]
  output [54:0] io_result // @[:@53155.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@53160.4]
  wire [54:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@53160.4]
  fix2fixBox_64 fix2fixBox ( // @[BigIPZynq.scala 219:30:@53160.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@53168.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@53163.4]
endmodule
module Divider( // @[:@53183.2]
  input         clock, // @[:@53184.4]
  input         io_flow, // @[:@53186.4]
  input  [54:0] io_dividend, // @[:@53186.4]
  input  [31:0] io_divisor, // @[:@53186.4]
  output [54:0] io_out // @[:@53186.4]
);
  wire [54:0] m_m_axis_dout_tdata; // @[ZynqBlackBoxes.scala 26:19:@53188.4]
  wire  m_m_axis_dout_tvalid; // @[ZynqBlackBoxes.scala 26:19:@53188.4]
  wire [31:0] m_s_axis_divisor_tdata; // @[ZynqBlackBoxes.scala 26:19:@53188.4]
  wire  m_s_axis_divisor_tvalid; // @[ZynqBlackBoxes.scala 26:19:@53188.4]
  wire [54:0] m_s_axis_dividend_tdata; // @[ZynqBlackBoxes.scala 26:19:@53188.4]
  wire  m_s_axis_dividend_tvalid; // @[ZynqBlackBoxes.scala 26:19:@53188.4]
  wire  m_aclken; // @[ZynqBlackBoxes.scala 26:19:@53188.4]
  wire  m_aclk; // @[ZynqBlackBoxes.scala 26:19:@53188.4]
  wire [52:0] _T_15; // @[ZynqBlackBoxes.scala 34:37:@53204.4]
  div_55_32_20_Signed_Fractional m ( // @[ZynqBlackBoxes.scala 26:19:@53188.4]
    .m_axis_dout_tdata(m_m_axis_dout_tdata),
    .m_axis_dout_tvalid(m_m_axis_dout_tvalid),
    .s_axis_divisor_tdata(m_s_axis_divisor_tdata),
    .s_axis_divisor_tvalid(m_s_axis_divisor_tvalid),
    .s_axis_dividend_tdata(m_s_axis_dividend_tdata),
    .s_axis_dividend_tvalid(m_s_axis_dividend_tvalid),
    .aclken(m_aclken),
    .aclk(m_aclk)
  );
  assign _T_15 = m_m_axis_dout_tdata[54:2]; // @[ZynqBlackBoxes.scala 34:37:@53204.4]
  assign io_out = {{2'd0}, _T_15}; // @[ZynqBlackBoxes.scala 34:12:@53205.4]
  assign m_s_axis_divisor_tdata = io_divisor; // @[ZynqBlackBoxes.scala 32:31:@53202.4]
  assign m_s_axis_divisor_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 31:32:@53201.4]
  assign m_s_axis_dividend_tdata = io_dividend; // @[ZynqBlackBoxes.scala 30:32:@53200.4]
  assign m_s_axis_dividend_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 29:33:@53199.4]
  assign m_aclken = io_flow; // @[ZynqBlackBoxes.scala 28:17:@53198.4 ZynqBlackBoxes.scala 33:17:@53203.4]
  assign m_aclk = clock; // @[ZynqBlackBoxes.scala 27:15:@53197.4]
endmodule
module fix2fixBox_65( // @[:@53271.2]
  input  [32:0] io_a, // @[:@53274.4]
  output [31:0] io_b // @[:@53274.4]
);
  wire [21:0] tmp_frac; // @[Converter.scala 38:42:@53282.4]
  wire [9:0] new_dec; // @[Converter.scala 88:34:@53285.4]
  assign tmp_frac = io_a[22:1]; // @[Converter.scala 38:42:@53282.4]
  assign new_dec = io_a[32:23]; // @[Converter.scala 88:34:@53285.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@53288.4]
endmodule
module x611_div( // @[:@53290.2]
  input         clock, // @[:@53291.4]
  input         reset, // @[:@53292.4]
  input  [31:0] io_a, // @[:@53293.4]
  input  [31:0] io_b, // @[:@53293.4]
  output [31:0] io_result // @[:@53293.4]
);
  wire [31:0] cast_x611_div_io_b; // @[Math.scala 720:24:@53301.4]
  wire [54:0] cast_x611_div_io_result; // @[Math.scala 720:24:@53301.4]
  wire  x611_div_clock; // @[BigIPZynq.scala 25:21:@53311.4]
  wire  x611_div_io_flow; // @[BigIPZynq.scala 25:21:@53311.4]
  wire [54:0] x611_div_io_dividend; // @[BigIPZynq.scala 25:21:@53311.4]
  wire [31:0] x611_div_io_divisor; // @[BigIPZynq.scala 25:21:@53311.4]
  wire [54:0] x611_div_io_out; // @[BigIPZynq.scala 25:21:@53311.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@53326.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@53326.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@53326.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@53326.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@53326.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@53337.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@53337.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@53337.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@53337.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@53337.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 317:32:@53344.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 317:32:@53344.4]
  wire [54:0] _T_21_number; // @[Math.scala 723:22:@53306.4 Math.scala 724:14:@53307.4]
  wire [54:0] _T_22; // @[FixedPoint.scala 33:34:@53309.4]
  wire [31:0] _T_23; // @[FixedPoint.scala 24:59:@53310.4]
  wire [54:0] _T_26; // @[BigIPZynq.scala 29:16:@53319.4]
  wire [54:0] _T_27; // @[Math.scala 307:88:@53320.4]
  wire  _T_30; // @[FixedPoint.scala 50:25:@53323.4]
  wire  _T_31; // @[FixedPoint.scala 50:25:@53324.4]
  wire  _T_32; // @[Math.scala 315:58:@53325.4]
  cast_x611_div cast_x611_div ( // @[Math.scala 720:24:@53301.4]
    .io_b(cast_x611_div_io_b),
    .io_result(cast_x611_div_io_result)
  );
  Divider x611_div ( // @[BigIPZynq.scala 25:21:@53311.4]
    .clock(x611_div_clock),
    .io_flow(x611_div_io_flow),
    .io_dividend(x611_div_io_dividend),
    .io_divisor(x611_div_io_divisor),
    .io_out(x611_div_io_out)
  );
  RetimeWrapper_520 RetimeWrapper ( // @[package.scala 93:22:@53326.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_520 RetimeWrapper_1 ( // @[package.scala 93:22:@53337.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  fix2fixBox_65 fix2fixBox ( // @[Math.scala 317:32:@53344.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_21_number = cast_x611_div_io_result; // @[Math.scala 723:22:@53306.4 Math.scala 724:14:@53307.4]
  assign _T_22 = $signed(_T_21_number); // @[FixedPoint.scala 33:34:@53309.4]
  assign _T_23 = $signed(io_b); // @[FixedPoint.scala 24:59:@53310.4]
  assign _T_26 = $signed(x611_div_io_out); // @[BigIPZynq.scala 29:16:@53319.4]
  assign _T_27 = $unsigned(_T_26); // @[Math.scala 307:88:@53320.4]
  assign _T_30 = io_a[31]; // @[FixedPoint.scala 50:25:@53323.4]
  assign _T_31 = io_b[31]; // @[FixedPoint.scala 50:25:@53324.4]
  assign _T_32 = _T_30 ^ _T_31; // @[Math.scala 315:58:@53325.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 323:19:@53352.4]
  assign cast_x611_div_io_b = io_a; // @[Math.scala 721:17:@53304.4]
  assign x611_div_clock = clock; // @[:@53312.4]
  assign x611_div_io_flow = 1'h1; // @[BigIPZynq.scala 28:17:@53318.4]
  assign x611_div_io_dividend = $unsigned(_T_22); // @[BigIPZynq.scala 26:21:@53315.4]
  assign x611_div_io_divisor = $unsigned(_T_23); // @[BigIPZynq.scala 27:20:@53317.4]
  assign RetimeWrapper_clock = clock; // @[:@53327.4]
  assign RetimeWrapper_reset = reset; // @[:@53328.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@53330.4]
  assign RetimeWrapper_io_in = _T_30 ^ _T_31; // @[package.scala 94:16:@53329.4]
  assign RetimeWrapper_1_clock = clock; // @[:@53338.4]
  assign RetimeWrapper_1_reset = reset; // @[:@53339.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@53341.4]
  assign RetimeWrapper_1_io_in = _T_32 == 1'h0; // @[package.scala 94:16:@53340.4]
  assign fix2fixBox_io_a = _T_27[32:0]; // @[Math.scala 318:25:@53347.4]
endmodule
module RetimeWrapper_615( // @[:@53366.2]
  input         clock, // @[:@53367.4]
  input         reset, // @[:@53368.4]
  input  [31:0] io_in, // @[:@53369.4]
  output [31:0] io_out // @[:@53369.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@53371.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@53371.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@53371.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@53371.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@53371.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@53371.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@53371.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@53384.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@53383.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@53382.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@53381.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@53380.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@53378.4]
endmodule
module RetimeWrapper_618( // @[:@53620.2]
  input         clock, // @[:@53621.4]
  input         reset, // @[:@53622.4]
  input  [31:0] io_in, // @[:@53623.4]
  output [31:0] io_out // @[:@53623.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@53625.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@53625.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@53625.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@53625.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@53625.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@53625.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(40)) sr ( // @[RetimeShiftRegister.scala 15:20:@53625.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@53638.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@53637.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@53636.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@53635.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@53634.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@53632.4]
endmodule
module RetimeWrapper_621( // @[:@53874.2]
  input         clock, // @[:@53875.4]
  input         reset, // @[:@53876.4]
  input  [31:0] io_in, // @[:@53877.4]
  output [31:0] io_out // @[:@53877.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@53879.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@53879.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@53879.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@53879.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@53879.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@53879.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(60)) sr ( // @[RetimeShiftRegister.scala 15:20:@53879.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@53892.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@53891.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@53890.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@53889.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@53888.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@53886.4]
endmodule
module RetimeWrapper_624( // @[:@54128.2]
  input         clock, // @[:@54129.4]
  input         reset, // @[:@54130.4]
  input  [31:0] io_in, // @[:@54131.4]
  output [31:0] io_out // @[:@54131.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@54133.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@54133.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@54133.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@54133.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@54133.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@54133.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(80)) sr ( // @[RetimeShiftRegister.scala 15:20:@54133.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@54146.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@54145.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@54144.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@54143.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@54142.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@54140.4]
endmodule
module x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1( // @[:@55029.2]
  input         clock, // @[:@55030.4]
  input         reset, // @[:@55031.4]
  output        io_in_x580_r_0_rPort_1_en_0, // @[:@55032.4]
  input  [31:0] io_in_x580_r_0_rPort_1_output_0, // @[:@55032.4]
  input         io_in_x595_reg_rPort_1_output_0, // @[:@55032.4]
  input         io_sigsIn_datapathEn, // @[:@55032.4]
  input         io_sigsIn_break, // @[:@55032.4]
  input         io_rr, // @[:@55032.4]
  output [31:0] io_ret_number // @[:@55032.4]
);
  wire  x611_div_1_clock; // @[Math.scala 327:24:@55149.4]
  wire  x611_div_1_reset; // @[Math.scala 327:24:@55149.4]
  wire [31:0] x611_div_1_io_a; // @[Math.scala 327:24:@55149.4]
  wire [31:0] x611_div_1_io_b; // @[Math.scala 327:24:@55149.4]
  wire [31:0] x611_div_1_io_result; // @[Math.scala 327:24:@55149.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@55160.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@55160.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@55160.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@55160.4]
  wire  x612_div_1_clock; // @[Math.scala 327:24:@55169.4]
  wire  x612_div_1_reset; // @[Math.scala 327:24:@55169.4]
  wire [31:0] x612_div_1_io_a; // @[Math.scala 327:24:@55169.4]
  wire [31:0] x612_div_1_io_b; // @[Math.scala 327:24:@55169.4]
  wire [31:0] x612_div_1_io_result; // @[Math.scala 327:24:@55169.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@55180.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@55180.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@55180.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@55180.4]
  wire  x613_div_1_clock; // @[Math.scala 327:24:@55189.4]
  wire  x613_div_1_reset; // @[Math.scala 327:24:@55189.4]
  wire [31:0] x613_div_1_io_a; // @[Math.scala 327:24:@55189.4]
  wire [31:0] x613_div_1_io_b; // @[Math.scala 327:24:@55189.4]
  wire [31:0] x613_div_1_io_result; // @[Math.scala 327:24:@55189.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@55200.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@55200.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@55200.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@55200.4]
  wire  x614_div_1_clock; // @[Math.scala 327:24:@55209.4]
  wire  x614_div_1_reset; // @[Math.scala 327:24:@55209.4]
  wire [31:0] x614_div_1_io_a; // @[Math.scala 327:24:@55209.4]
  wire [31:0] x614_div_1_io_b; // @[Math.scala 327:24:@55209.4]
  wire [31:0] x614_div_1_io_result; // @[Math.scala 327:24:@55209.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@55220.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@55220.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@55220.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@55220.4]
  wire  x615_div_1_clock; // @[Math.scala 327:24:@55229.4]
  wire  x615_div_1_reset; // @[Math.scala 327:24:@55229.4]
  wire [31:0] x615_div_1_io_a; // @[Math.scala 327:24:@55229.4]
  wire [31:0] x615_div_1_io_b; // @[Math.scala 327:24:@55229.4]
  wire [31:0] x615_div_1_io_result; // @[Math.scala 327:24:@55229.4]
  wire  x616_div_1_clock; // @[Math.scala 327:24:@55241.4]
  wire  x616_div_1_reset; // @[Math.scala 327:24:@55241.4]
  wire [31:0] x616_div_1_io_a; // @[Math.scala 327:24:@55241.4]
  wire [31:0] x616_div_1_io_b; // @[Math.scala 327:24:@55241.4]
  wire [31:0] x616_div_1_io_result; // @[Math.scala 327:24:@55241.4]
  wire  x617_div_1_clock; // @[Math.scala 327:24:@55251.4]
  wire  x617_div_1_reset; // @[Math.scala 327:24:@55251.4]
  wire [31:0] x617_div_1_io_a; // @[Math.scala 327:24:@55251.4]
  wire [31:0] x617_div_1_io_b; // @[Math.scala 327:24:@55251.4]
  wire [31:0] x617_div_1_io_result; // @[Math.scala 327:24:@55251.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@55262.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@55262.4]
  wire [31:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@55262.4]
  wire [31:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@55262.4]
  wire  x618_sub_1_clock; // @[Math.scala 191:24:@55271.4]
  wire  x618_sub_1_reset; // @[Math.scala 191:24:@55271.4]
  wire [31:0] x618_sub_1_io_a; // @[Math.scala 191:24:@55271.4]
  wire [31:0] x618_sub_1_io_b; // @[Math.scala 191:24:@55271.4]
  wire [31:0] x618_sub_1_io_result; // @[Math.scala 191:24:@55271.4]
  wire  _T_664; // @[sm_x619_inr_SwitchCase.scala 66:119:@55113.4]
  wire  _T_665; // @[sm_x619_inr_SwitchCase.scala 66:116:@55114.4]
  wire  _T_670; // @[implicits.scala 56:10:@55117.4]
  wire  x608_rd_x595_shared_en; // @[sm_x619_inr_SwitchCase.scala 66:136:@55118.4]
  x611_div x611_div_1 ( // @[Math.scala 327:24:@55149.4]
    .clock(x611_div_1_clock),
    .reset(x611_div_1_reset),
    .io_a(x611_div_1_io_a),
    .io_b(x611_div_1_io_b),
    .io_result(x611_div_1_io_result)
  );
  RetimeWrapper_615 RetimeWrapper ( // @[package.scala 93:22:@55160.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x611_div x612_div_1 ( // @[Math.scala 327:24:@55169.4]
    .clock(x612_div_1_clock),
    .reset(x612_div_1_reset),
    .io_a(x612_div_1_io_a),
    .io_b(x612_div_1_io_b),
    .io_result(x612_div_1_io_result)
  );
  RetimeWrapper_618 RetimeWrapper_1 ( // @[package.scala 93:22:@55180.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x611_div x613_div_1 ( // @[Math.scala 327:24:@55189.4]
    .clock(x613_div_1_clock),
    .reset(x613_div_1_reset),
    .io_a(x613_div_1_io_a),
    .io_b(x613_div_1_io_b),
    .io_result(x613_div_1_io_result)
  );
  RetimeWrapper_621 RetimeWrapper_2 ( // @[package.scala 93:22:@55200.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x611_div x614_div_1 ( // @[Math.scala 327:24:@55209.4]
    .clock(x614_div_1_clock),
    .reset(x614_div_1_reset),
    .io_a(x614_div_1_io_a),
    .io_b(x614_div_1_io_b),
    .io_result(x614_div_1_io_result)
  );
  RetimeWrapper_624 RetimeWrapper_3 ( // @[package.scala 93:22:@55220.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x611_div x615_div_1 ( // @[Math.scala 327:24:@55229.4]
    .clock(x615_div_1_clock),
    .reset(x615_div_1_reset),
    .io_a(x615_div_1_io_a),
    .io_b(x615_div_1_io_b),
    .io_result(x615_div_1_io_result)
  );
  x611_div x616_div_1 ( // @[Math.scala 327:24:@55241.4]
    .clock(x616_div_1_clock),
    .reset(x616_div_1_reset),
    .io_a(x616_div_1_io_a),
    .io_b(x616_div_1_io_b),
    .io_result(x616_div_1_io_result)
  );
  x611_div x617_div_1 ( // @[Math.scala 327:24:@55251.4]
    .clock(x617_div_1_clock),
    .reset(x617_div_1_reset),
    .io_a(x617_div_1_io_a),
    .io_b(x617_div_1_io_b),
    .io_result(x617_div_1_io_result)
  );
  RetimeWrapper_621 RetimeWrapper_4 ( // @[package.scala 93:22:@55262.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x573_sub x618_sub_1 ( // @[Math.scala 191:24:@55271.4]
    .clock(x618_sub_1_clock),
    .reset(x618_sub_1_reset),
    .io_a(x618_sub_1_io_a),
    .io_b(x618_sub_1_io_b),
    .io_result(x618_sub_1_io_result)
  );
  assign _T_664 = ~ io_sigsIn_break; // @[sm_x619_inr_SwitchCase.scala 66:119:@55113.4]
  assign _T_665 = io_rr & _T_664; // @[sm_x619_inr_SwitchCase.scala 66:116:@55114.4]
  assign _T_670 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 56:10:@55117.4]
  assign x608_rd_x595_shared_en = _T_665 & _T_670; // @[sm_x619_inr_SwitchCase.scala 66:136:@55118.4]
  assign io_in_x580_r_0_rPort_1_en_0 = x608_rd_x595_shared_en & io_in_x595_reg_rPort_1_output_0; // @[MemInterfaceType.scala 110:79:@55142.4]
  assign io_ret_number = x618_sub_1_io_result; // @[sm_x619_inr_SwitchCase.scala 103:16:@55280.4]
  assign x611_div_1_clock = clock; // @[:@55150.4]
  assign x611_div_1_reset = reset; // @[:@55151.4]
  assign x611_div_1_io_a = 32'h19000000; // @[Math.scala 328:17:@55152.4]
  assign x611_div_1_io_b = io_in_x580_r_0_rPort_1_output_0; // @[Math.scala 329:17:@55153.4]
  assign RetimeWrapper_clock = clock; // @[:@55161.4]
  assign RetimeWrapper_reset = reset; // @[:@55162.4]
  assign RetimeWrapper_io_in = io_in_x580_r_0_rPort_1_output_0; // @[package.scala 94:16:@55163.4]
  assign x612_div_1_clock = clock; // @[:@55170.4]
  assign x612_div_1_reset = reset; // @[:@55171.4]
  assign x612_div_1_io_a = x611_div_1_io_result; // @[Math.scala 328:17:@55172.4]
  assign x612_div_1_io_b = RetimeWrapper_io_out; // @[Math.scala 329:17:@55173.4]
  assign RetimeWrapper_1_clock = clock; // @[:@55181.4]
  assign RetimeWrapper_1_reset = reset; // @[:@55182.4]
  assign RetimeWrapper_1_io_in = io_in_x580_r_0_rPort_1_output_0; // @[package.scala 94:16:@55183.4]
  assign x613_div_1_clock = clock; // @[:@55190.4]
  assign x613_div_1_reset = reset; // @[:@55191.4]
  assign x613_div_1_io_a = x612_div_1_io_result; // @[Math.scala 328:17:@55192.4]
  assign x613_div_1_io_b = RetimeWrapper_1_io_out; // @[Math.scala 329:17:@55193.4]
  assign RetimeWrapper_2_clock = clock; // @[:@55201.4]
  assign RetimeWrapper_2_reset = reset; // @[:@55202.4]
  assign RetimeWrapper_2_io_in = io_in_x580_r_0_rPort_1_output_0; // @[package.scala 94:16:@55203.4]
  assign x614_div_1_clock = clock; // @[:@55210.4]
  assign x614_div_1_reset = reset; // @[:@55211.4]
  assign x614_div_1_io_a = x613_div_1_io_result; // @[Math.scala 328:17:@55212.4]
  assign x614_div_1_io_b = RetimeWrapper_2_io_out; // @[Math.scala 329:17:@55213.4]
  assign RetimeWrapper_3_clock = clock; // @[:@55221.4]
  assign RetimeWrapper_3_reset = reset; // @[:@55222.4]
  assign RetimeWrapper_3_io_in = io_in_x580_r_0_rPort_1_output_0; // @[package.scala 94:16:@55223.4]
  assign x615_div_1_clock = clock; // @[:@55230.4]
  assign x615_div_1_reset = reset; // @[:@55231.4]
  assign x615_div_1_io_a = x614_div_1_io_result; // @[Math.scala 328:17:@55232.4]
  assign x615_div_1_io_b = RetimeWrapper_3_io_out; // @[Math.scala 329:17:@55233.4]
  assign x616_div_1_clock = clock; // @[:@55242.4]
  assign x616_div_1_reset = reset; // @[:@55243.4]
  assign x616_div_1_io_a = 32'h2800000; // @[Math.scala 328:17:@55244.4]
  assign x616_div_1_io_b = io_in_x580_r_0_rPort_1_output_0; // @[Math.scala 329:17:@55245.4]
  assign x617_div_1_clock = clock; // @[:@55252.4]
  assign x617_div_1_reset = reset; // @[:@55253.4]
  assign x617_div_1_io_a = x616_div_1_io_result; // @[Math.scala 328:17:@55254.4]
  assign x617_div_1_io_b = RetimeWrapper_io_out; // @[Math.scala 329:17:@55255.4]
  assign RetimeWrapper_4_clock = clock; // @[:@55263.4]
  assign RetimeWrapper_4_reset = reset; // @[:@55264.4]
  assign RetimeWrapper_4_io_in = x617_div_1_io_result; // @[package.scala 94:16:@55265.4]
  assign x618_sub_1_clock = clock; // @[:@55272.4]
  assign x618_sub_1_reset = reset; // @[:@55273.4]
  assign x618_sub_1_io_a = x615_div_1_io_result; // @[Math.scala 192:17:@55274.4]
  assign x618_sub_1_io_b = RetimeWrapper_4_io_out; // @[Math.scala 193:17:@55275.4]
endmodule
module x621_inr_Switch_kernelx621_inr_Switch_concrete1( // @[:@55862.2]
  input         clock, // @[:@55863.4]
  input         reset, // @[:@55864.4]
  output        io_in_x555_tmp_1_sEn_3, // @[:@55865.4]
  output        io_in_x555_tmp_1_sDone_3, // @[:@55865.4]
  output        io_in_x554_tmp_0_sEn_3, // @[:@55865.4]
  output        io_in_x554_tmp_0_sDone_3, // @[:@55865.4]
  output        io_in_x558_tmp_4_sEn_3, // @[:@55865.4]
  output        io_in_x558_tmp_4_sDone_3, // @[:@55865.4]
  input         io_in_x736_rd_x596, // @[:@55865.4]
  output        io_in_x557_tmp_3_sEn_3, // @[:@55865.4]
  output        io_in_x557_tmp_3_sDone_3, // @[:@55865.4]
  output        io_in_x580_r_0_rPort_1_en_0, // @[:@55865.4]
  input  [31:0] io_in_x580_r_0_rPort_1_output_0, // @[:@55865.4]
  output        io_in_x580_r_0_sEn_2, // @[:@55865.4]
  output        io_in_x580_r_0_sDone_2, // @[:@55865.4]
  input         io_in_x595_reg_rPort_1_output_0, // @[:@55865.4]
  output        io_in_x595_reg_sEn_1, // @[:@55865.4]
  output        io_in_x595_reg_sDone_1, // @[:@55865.4]
  output        io_in_x556_tmp_2_sEn_3, // @[:@55865.4]
  output        io_in_x556_tmp_2_sDone_3, // @[:@55865.4]
  input         io_in_x735_rd_x595, // @[:@55865.4]
  output        io_in_x596_reg_sEn_1, // @[:@55865.4]
  output        io_in_x596_reg_sDone_1, // @[:@55865.4]
  input         io_sigsIn_done, // @[:@55865.4]
  input         io_sigsIn_baseEn, // @[:@55865.4]
  input         io_sigsIn_smSelectsOut_0, // @[:@55865.4]
  input         io_sigsIn_smSelectsOut_1, // @[:@55865.4]
  input         io_sigsIn_smChildAcks_0, // @[:@55865.4]
  input         io_sigsIn_smChildAcks_1, // @[:@55865.4]
  output        io_sigsOut_smDoneIn_0, // @[:@55865.4]
  output        io_sigsOut_smDoneIn_1, // @[:@55865.4]
  input         io_rr, // @[:@55865.4]
  output [31:0] io_ret_number // @[:@55865.4]
);
  wire  x619_inr_SwitchCase_sm_clock; // @[sm_x619_inr_SwitchCase.scala 32:18:@56224.4]
  wire  x619_inr_SwitchCase_sm_reset; // @[sm_x619_inr_SwitchCase.scala 32:18:@56224.4]
  wire  x619_inr_SwitchCase_sm_io_enable; // @[sm_x619_inr_SwitchCase.scala 32:18:@56224.4]
  wire  x619_inr_SwitchCase_sm_io_done; // @[sm_x619_inr_SwitchCase.scala 32:18:@56224.4]
  wire  x619_inr_SwitchCase_sm_io_ctrDone; // @[sm_x619_inr_SwitchCase.scala 32:18:@56224.4]
  wire  x619_inr_SwitchCase_sm_io_datapathEn; // @[sm_x619_inr_SwitchCase.scala 32:18:@56224.4]
  wire  x619_inr_SwitchCase_sm_io_ctrInc; // @[sm_x619_inr_SwitchCase.scala 32:18:@56224.4]
  wire  x619_inr_SwitchCase_sm_io_parentAck; // @[sm_x619_inr_SwitchCase.scala 32:18:@56224.4]
  wire  x619_inr_SwitchCase_sm_io_break; // @[sm_x619_inr_SwitchCase.scala 32:18:@56224.4]
  wire  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_clock; // @[sm_x619_inr_SwitchCase.scala 105:24:@56302.4]
  wire  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_reset; // @[sm_x619_inr_SwitchCase.scala 105:24:@56302.4]
  wire  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x580_r_0_rPort_1_en_0; // @[sm_x619_inr_SwitchCase.scala 105:24:@56302.4]
  wire [31:0] x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x580_r_0_rPort_1_output_0; // @[sm_x619_inr_SwitchCase.scala 105:24:@56302.4]
  wire  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x595_reg_rPort_1_output_0; // @[sm_x619_inr_SwitchCase.scala 105:24:@56302.4]
  wire  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_datapathEn; // @[sm_x619_inr_SwitchCase.scala 105:24:@56302.4]
  wire  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_break; // @[sm_x619_inr_SwitchCase.scala 105:24:@56302.4]
  wire  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_rr; // @[sm_x619_inr_SwitchCase.scala 105:24:@56302.4]
  wire [31:0] x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_ret_number; // @[sm_x619_inr_SwitchCase.scala 105:24:@56302.4]
  wire  x620_inr_SwitchCase_sm_clock; // @[sm_x620_inr_SwitchCase.scala 31:18:@56508.4]
  wire  x620_inr_SwitchCase_sm_reset; // @[sm_x620_inr_SwitchCase.scala 31:18:@56508.4]
  wire  x620_inr_SwitchCase_sm_io_enable; // @[sm_x620_inr_SwitchCase.scala 31:18:@56508.4]
  wire  x620_inr_SwitchCase_sm_io_done; // @[sm_x620_inr_SwitchCase.scala 31:18:@56508.4]
  wire  x620_inr_SwitchCase_sm_io_ctrDone; // @[sm_x620_inr_SwitchCase.scala 31:18:@56508.4]
  wire  x620_inr_SwitchCase_sm_io_datapathEn; // @[sm_x620_inr_SwitchCase.scala 31:18:@56508.4]
  wire  x620_inr_SwitchCase_sm_io_ctrInc; // @[sm_x620_inr_SwitchCase.scala 31:18:@56508.4]
  wire  x620_inr_SwitchCase_sm_io_parentAck; // @[sm_x620_inr_SwitchCase.scala 31:18:@56508.4]
  wire  x620_inr_SwitchCase_sm_io_break; // @[sm_x620_inr_SwitchCase.scala 31:18:@56508.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@56662.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@56662.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@56662.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@56662.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@56662.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@56673.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@56673.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@56673.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@56673.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@56673.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@56684.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@56684.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@56684.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@56684.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@56684.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@56695.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@56695.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@56695.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@56695.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@56695.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@56706.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@56706.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@56706.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@56706.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@56706.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@56717.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@56717.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@56717.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@56717.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@56717.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@56728.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@56728.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@56728.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@56728.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@56728.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@56739.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@56739.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@56739.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@56739.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@56739.4]
  wire  _T_2361; // @[package.scala 100:49:@56253.4]
  reg  _T_2364; // @[package.scala 48:56:@56254.4]
  reg [31:0] _RAND_0;
  wire  _T_2444; // @[package.scala 100:49:@56537.4]
  reg  _T_2447; // @[package.scala 48:56:@56538.4]
  reg [31:0] _RAND_1;
  wire [31:0] x619_inr_SwitchCase_number; // @[sm_x621_inr_Switch.scala 101:37:@56265.4 sm_x621_inr_Switch.scala 104:29:@56471.4]
  wire [31:0] _T_2485; // @[Mux.scala 19:72:@56652.4]
  wire [31:0] _T_2487; // @[Mux.scala 19:72:@56653.4]
  wire  _T_2497; // @[package.scala 96:25:@56667.4 package.scala 96:25:@56668.4]
  wire  _T_2503; // @[package.scala 96:25:@56678.4 package.scala 96:25:@56679.4]
  wire  _T_2509; // @[package.scala 96:25:@56689.4 package.scala 96:25:@56690.4]
  wire  _T_2515; // @[package.scala 96:25:@56700.4 package.scala 96:25:@56701.4]
  wire  _T_2521; // @[package.scala 96:25:@56711.4 package.scala 96:25:@56712.4]
  wire  _T_2527; // @[package.scala 96:25:@56722.4 package.scala 96:25:@56723.4]
  wire  _T_2533; // @[package.scala 96:25:@56733.4 package.scala 96:25:@56734.4]
  wire  _T_2539; // @[package.scala 96:25:@56744.4 package.scala 96:25:@56745.4]
  x619_inr_SwitchCase_sm x619_inr_SwitchCase_sm ( // @[sm_x619_inr_SwitchCase.scala 32:18:@56224.4]
    .clock(x619_inr_SwitchCase_sm_clock),
    .reset(x619_inr_SwitchCase_sm_reset),
    .io_enable(x619_inr_SwitchCase_sm_io_enable),
    .io_done(x619_inr_SwitchCase_sm_io_done),
    .io_ctrDone(x619_inr_SwitchCase_sm_io_ctrDone),
    .io_datapathEn(x619_inr_SwitchCase_sm_io_datapathEn),
    .io_ctrInc(x619_inr_SwitchCase_sm_io_ctrInc),
    .io_parentAck(x619_inr_SwitchCase_sm_io_parentAck),
    .io_break(x619_inr_SwitchCase_sm_io_break)
  );
  x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1 x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1 ( // @[sm_x619_inr_SwitchCase.scala 105:24:@56302.4]
    .clock(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_clock),
    .reset(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_reset),
    .io_in_x580_r_0_rPort_1_en_0(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x580_r_0_rPort_1_en_0),
    .io_in_x580_r_0_rPort_1_output_0(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x580_r_0_rPort_1_output_0),
    .io_in_x595_reg_rPort_1_output_0(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x595_reg_rPort_1_output_0),
    .io_sigsIn_datapathEn(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_break),
    .io_rr(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_rr),
    .io_ret_number(x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_ret_number)
  );
  x619_inr_SwitchCase_sm x620_inr_SwitchCase_sm ( // @[sm_x620_inr_SwitchCase.scala 31:18:@56508.4]
    .clock(x620_inr_SwitchCase_sm_clock),
    .reset(x620_inr_SwitchCase_sm_reset),
    .io_enable(x620_inr_SwitchCase_sm_io_enable),
    .io_done(x620_inr_SwitchCase_sm_io_done),
    .io_ctrDone(x620_inr_SwitchCase_sm_io_ctrDone),
    .io_datapathEn(x620_inr_SwitchCase_sm_io_datapathEn),
    .io_ctrInc(x620_inr_SwitchCase_sm_io_ctrInc),
    .io_parentAck(x620_inr_SwitchCase_sm_io_parentAck),
    .io_break(x620_inr_SwitchCase_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@56662.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@56673.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@56684.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@56695.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@56706.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@56717.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@56728.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@56739.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign _T_2361 = x619_inr_SwitchCase_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@56253.4]
  assign _T_2444 = x620_inr_SwitchCase_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@56537.4]
  assign x619_inr_SwitchCase_number = x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_ret_number; // @[sm_x621_inr_Switch.scala 101:37:@56265.4 sm_x621_inr_Switch.scala 104:29:@56471.4]
  assign _T_2485 = io_in_x735_rd_x595 ? x619_inr_SwitchCase_number : 32'h0; // @[Mux.scala 19:72:@56652.4]
  assign _T_2487 = io_in_x736_rd_x596 ? 32'h16800000 : 32'h0; // @[Mux.scala 19:72:@56653.4]
  assign _T_2497 = RetimeWrapper_io_out; // @[package.scala 96:25:@56667.4 package.scala 96:25:@56668.4]
  assign _T_2503 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@56678.4 package.scala 96:25:@56679.4]
  assign _T_2509 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@56689.4 package.scala 96:25:@56690.4]
  assign _T_2515 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@56700.4 package.scala 96:25:@56701.4]
  assign _T_2521 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@56711.4 package.scala 96:25:@56712.4]
  assign _T_2527 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@56722.4 package.scala 96:25:@56723.4]
  assign _T_2533 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@56733.4 package.scala 96:25:@56734.4]
  assign _T_2539 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@56744.4 package.scala 96:25:@56745.4]
  assign io_in_x555_tmp_1_sEn_3 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@56681.4]
  assign io_in_x555_tmp_1_sDone_3 = io_rr ? _T_2503 : 1'h0; // @[MemInterfaceType.scala 197:17:@56682.4]
  assign io_in_x554_tmp_0_sEn_3 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@56670.4]
  assign io_in_x554_tmp_0_sDone_3 = io_rr ? _T_2497 : 1'h0; // @[MemInterfaceType.scala 197:17:@56671.4]
  assign io_in_x558_tmp_4_sEn_3 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@56714.4]
  assign io_in_x558_tmp_4_sDone_3 = io_rr ? _T_2521 : 1'h0; // @[MemInterfaceType.scala 197:17:@56715.4]
  assign io_in_x557_tmp_3_sEn_3 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@56703.4]
  assign io_in_x557_tmp_3_sDone_3 = io_rr ? _T_2515 : 1'h0; // @[MemInterfaceType.scala 197:17:@56704.4]
  assign io_in_x580_r_0_rPort_1_en_0 = x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x580_r_0_rPort_1_en_0; // @[MemInterfaceType.scala 66:44:@56420.4]
  assign io_in_x580_r_0_sEn_2 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@56725.4]
  assign io_in_x580_r_0_sDone_2 = io_rr ? _T_2527 : 1'h0; // @[MemInterfaceType.scala 197:17:@56726.4]
  assign io_in_x595_reg_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@56736.4]
  assign io_in_x595_reg_sDone_1 = io_rr ? _T_2533 : 1'h0; // @[MemInterfaceType.scala 197:17:@56737.4]
  assign io_in_x556_tmp_2_sEn_3 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@56692.4]
  assign io_in_x556_tmp_2_sDone_3 = io_rr ? _T_2509 : 1'h0; // @[MemInterfaceType.scala 197:17:@56693.4]
  assign io_in_x596_reg_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@56747.4]
  assign io_in_x596_reg_sDone_1 = io_rr ? _T_2539 : 1'h0; // @[MemInterfaceType.scala 197:17:@56748.4]
  assign io_sigsOut_smDoneIn_0 = x619_inr_SwitchCase_sm_io_done; // @[SpatialBlocks.scala 155:56:@56288.4]
  assign io_sigsOut_smDoneIn_1 = x620_inr_SwitchCase_sm_io_done; // @[SpatialBlocks.scala 155:56:@56572.4]
  assign io_ret_number = _T_2485 | _T_2487; // @[sm_x621_inr_Switch.scala 122:16:@56660.4]
  assign x619_inr_SwitchCase_sm_clock = clock; // @[:@56225.4]
  assign x619_inr_SwitchCase_sm_reset = reset; // @[:@56226.4]
  assign x619_inr_SwitchCase_sm_io_enable = io_sigsIn_smSelectsOut_0; // @[SpatialBlocks.scala 139:18:@56285.4]
  assign x619_inr_SwitchCase_sm_io_ctrDone = x619_inr_SwitchCase_sm_io_ctrInc & _T_2364; // @[sm_x621_inr_Switch.scala 96:45:@56257.4]
  assign x619_inr_SwitchCase_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@56287.4]
  assign x619_inr_SwitchCase_sm_io_break = 1'h0; // @[sm_x621_inr_Switch.scala 100:43:@56264.4]
  assign x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_clock = clock; // @[:@56303.4]
  assign x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_reset = reset; // @[:@56304.4]
  assign x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x580_r_0_rPort_1_output_0 = io_in_x580_r_0_rPort_1_output_0; // @[MemInterfaceType.scala 66:44:@56418.4]
  assign x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_in_x595_reg_rPort_1_output_0 = io_in_x595_reg_rPort_1_output_0; // @[MemInterfaceType.scala 66:44:@56439.4]
  assign x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_datapathEn = x619_inr_SwitchCase_sm_io_datapathEn; // @[sm_x619_inr_SwitchCase.scala 110:22:@56456.4]
  assign x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_sigsIn_break = x619_inr_SwitchCase_sm_io_break; // @[sm_x619_inr_SwitchCase.scala 110:22:@56454.4]
  assign x619_inr_SwitchCase_kernelx619_inr_SwitchCase_concrete1_io_rr = io_rr; // @[sm_x619_inr_SwitchCase.scala 109:18:@56444.4]
  assign x620_inr_SwitchCase_sm_clock = clock; // @[:@56509.4]
  assign x620_inr_SwitchCase_sm_reset = reset; // @[:@56510.4]
  assign x620_inr_SwitchCase_sm_io_enable = io_sigsIn_smSelectsOut_1; // @[SpatialBlocks.scala 139:18:@56569.4]
  assign x620_inr_SwitchCase_sm_io_ctrDone = x620_inr_SwitchCase_sm_io_ctrInc & _T_2447; // @[sm_x621_inr_Switch.scala 107:45:@56541.4]
  assign x620_inr_SwitchCase_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 141:21:@56571.4]
  assign x620_inr_SwitchCase_sm_io_break = 1'h0; // @[sm_x621_inr_Switch.scala 111:43:@56548.4]
  assign RetimeWrapper_clock = clock; // @[:@56663.4]
  assign RetimeWrapper_reset = reset; // @[:@56664.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@56666.4]
  assign RetimeWrapper_io_in = io_sigsIn_done; // @[package.scala 94:16:@56665.4]
  assign RetimeWrapper_1_clock = clock; // @[:@56674.4]
  assign RetimeWrapper_1_reset = reset; // @[:@56675.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@56677.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_done; // @[package.scala 94:16:@56676.4]
  assign RetimeWrapper_2_clock = clock; // @[:@56685.4]
  assign RetimeWrapper_2_reset = reset; // @[:@56686.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@56688.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_done; // @[package.scala 94:16:@56687.4]
  assign RetimeWrapper_3_clock = clock; // @[:@56696.4]
  assign RetimeWrapper_3_reset = reset; // @[:@56697.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@56699.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_done; // @[package.scala 94:16:@56698.4]
  assign RetimeWrapper_4_clock = clock; // @[:@56707.4]
  assign RetimeWrapper_4_reset = reset; // @[:@56708.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@56710.4]
  assign RetimeWrapper_4_io_in = io_sigsIn_done; // @[package.scala 94:16:@56709.4]
  assign RetimeWrapper_5_clock = clock; // @[:@56718.4]
  assign RetimeWrapper_5_reset = reset; // @[:@56719.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@56721.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_done; // @[package.scala 94:16:@56720.4]
  assign RetimeWrapper_6_clock = clock; // @[:@56729.4]
  assign RetimeWrapper_6_reset = reset; // @[:@56730.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@56732.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_done; // @[package.scala 94:16:@56731.4]
  assign RetimeWrapper_7_clock = clock; // @[:@56740.4]
  assign RetimeWrapper_7_reset = reset; // @[:@56741.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@56743.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_done; // @[package.scala 94:16:@56742.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2364 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_2447 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_2364 <= 1'h0;
    end else begin
      _T_2364 <= _T_2361;
    end
    if (reset) begin
      _T_2447 <= 1'h0;
    end else begin
      _T_2447 <= _T_2444;
    end
  end
endmodule
module x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1( // @[:@57338.2]
  input         clock, // @[:@57339.4]
  input         reset, // @[:@57340.4]
  output        io_in_x555_tmp_1_sEn_4, // @[:@57341.4]
  output        io_in_x555_tmp_1_sDone_4, // @[:@57341.4]
  output        io_in_x554_tmp_0_sEn_4, // @[:@57341.4]
  output        io_in_x554_tmp_0_sDone_4, // @[:@57341.4]
  output        io_in_x558_tmp_4_sEn_4, // @[:@57341.4]
  output        io_in_x558_tmp_4_sDone_4, // @[:@57341.4]
  output [31:0] io_in_x594_force_0_wPort_0_data_0, // @[:@57341.4]
  output        io_in_x594_force_0_wPort_0_en_0, // @[:@57341.4]
  output        io_in_x594_force_0_sEn_0, // @[:@57341.4]
  output        io_in_x594_force_0_sDone_0, // @[:@57341.4]
  input  [31:0] io_in_x621_inr_Switch_number, // @[:@57341.4]
  output        io_in_x557_tmp_3_sEn_4, // @[:@57341.4]
  output        io_in_x557_tmp_3_sDone_4, // @[:@57341.4]
  output        io_in_x556_tmp_2_sEn_4, // @[:@57341.4]
  output        io_in_x556_tmp_2_sDone_4, // @[:@57341.4]
  input         io_sigsIn_done, // @[:@57341.4]
  input         io_sigsIn_datapathEn, // @[:@57341.4]
  input         io_sigsIn_baseEn, // @[:@57341.4]
  input         io_sigsIn_break, // @[:@57341.4]
  input         io_rr // @[:@57341.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@57614.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@57614.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@57614.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@57614.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@57614.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@57625.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@57625.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@57625.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@57625.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@57625.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@57636.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@57636.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@57636.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@57636.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@57636.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@57647.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@57647.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@57647.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@57647.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@57647.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@57658.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@57658.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@57658.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@57658.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@57658.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@57669.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@57669.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@57669.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@57669.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@57669.4]
  wire  _T_1771; // @[sm_x623_inr_UnitPipe.scala 94:100:@57598.4]
  wire  _T_1777; // @[implicits.scala 56:10:@57602.4]
  wire  _T_1778; // @[sm_x623_inr_UnitPipe.scala 94:117:@57603.4]
  wire  _T_1787; // @[package.scala 96:25:@57619.4 package.scala 96:25:@57620.4]
  wire  _T_1793; // @[package.scala 96:25:@57630.4 package.scala 96:25:@57631.4]
  wire  _T_1799; // @[package.scala 96:25:@57641.4 package.scala 96:25:@57642.4]
  wire  _T_1805; // @[package.scala 96:25:@57652.4 package.scala 96:25:@57653.4]
  wire  _T_1811; // @[package.scala 96:25:@57663.4 package.scala 96:25:@57664.4]
  wire  _T_1817; // @[package.scala 96:25:@57674.4 package.scala 96:25:@57675.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@57614.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@57625.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@57636.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@57647.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@57658.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@57669.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  assign _T_1771 = ~ io_sigsIn_break; // @[sm_x623_inr_UnitPipe.scala 94:100:@57598.4]
  assign _T_1777 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 56:10:@57602.4]
  assign _T_1778 = _T_1771 & _T_1777; // @[sm_x623_inr_UnitPipe.scala 94:117:@57603.4]
  assign _T_1787 = RetimeWrapper_io_out; // @[package.scala 96:25:@57619.4 package.scala 96:25:@57620.4]
  assign _T_1793 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@57630.4 package.scala 96:25:@57631.4]
  assign _T_1799 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@57641.4 package.scala 96:25:@57642.4]
  assign _T_1805 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@57652.4 package.scala 96:25:@57653.4]
  assign _T_1811 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@57663.4 package.scala 96:25:@57664.4]
  assign _T_1817 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@57674.4 package.scala 96:25:@57675.4]
  assign io_in_x555_tmp_1_sEn_4 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@57633.4]
  assign io_in_x555_tmp_1_sDone_4 = io_rr ? _T_1793 : 1'h0; // @[MemInterfaceType.scala 197:17:@57634.4]
  assign io_in_x554_tmp_0_sEn_4 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@57622.4]
  assign io_in_x554_tmp_0_sDone_4 = io_rr ? _T_1787 : 1'h0; // @[MemInterfaceType.scala 197:17:@57623.4]
  assign io_in_x558_tmp_4_sEn_4 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@57666.4]
  assign io_in_x558_tmp_4_sDone_4 = io_rr ? _T_1811 : 1'h0; // @[MemInterfaceType.scala 197:17:@57667.4]
  assign io_in_x594_force_0_wPort_0_data_0 = io_in_x621_inr_Switch_number; // @[MemInterfaceType.scala 90:56:@57610.4]
  assign io_in_x594_force_0_wPort_0_en_0 = _T_1778 & _T_1771; // @[MemInterfaceType.scala 93:57:@57612.4]
  assign io_in_x594_force_0_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@57677.4]
  assign io_in_x594_force_0_sDone_0 = io_rr ? _T_1817 : 1'h0; // @[MemInterfaceType.scala 197:17:@57678.4]
  assign io_in_x557_tmp_3_sEn_4 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@57655.4]
  assign io_in_x557_tmp_3_sDone_4 = io_rr ? _T_1805 : 1'h0; // @[MemInterfaceType.scala 197:17:@57656.4]
  assign io_in_x556_tmp_2_sEn_4 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@57644.4]
  assign io_in_x556_tmp_2_sDone_4 = io_rr ? _T_1799 : 1'h0; // @[MemInterfaceType.scala 197:17:@57645.4]
  assign RetimeWrapper_clock = clock; // @[:@57615.4]
  assign RetimeWrapper_reset = reset; // @[:@57616.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@57618.4]
  assign RetimeWrapper_io_in = io_sigsIn_done; // @[package.scala 94:16:@57617.4]
  assign RetimeWrapper_1_clock = clock; // @[:@57626.4]
  assign RetimeWrapper_1_reset = reset; // @[:@57627.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@57629.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_done; // @[package.scala 94:16:@57628.4]
  assign RetimeWrapper_2_clock = clock; // @[:@57637.4]
  assign RetimeWrapper_2_reset = reset; // @[:@57638.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@57640.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_done; // @[package.scala 94:16:@57639.4]
  assign RetimeWrapper_3_clock = clock; // @[:@57648.4]
  assign RetimeWrapper_3_reset = reset; // @[:@57649.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@57651.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_done; // @[package.scala 94:16:@57650.4]
  assign RetimeWrapper_4_clock = clock; // @[:@57659.4]
  assign RetimeWrapper_4_reset = reset; // @[:@57660.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@57662.4]
  assign RetimeWrapper_4_io_in = io_sigsIn_done; // @[package.scala 94:16:@57661.4]
  assign RetimeWrapper_5_clock = clock; // @[:@57670.4]
  assign RetimeWrapper_5_reset = reset; // @[:@57671.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@57673.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_done; // @[package.scala 94:16:@57672.4]
endmodule
module RetimeWrapper_660( // @[:@57881.2]
  input   clock, // @[:@57882.4]
  input   reset, // @[:@57883.4]
  input   io_in, // @[:@57884.4]
  output  io_out // @[:@57884.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@57886.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@57886.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@57886.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@57886.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@57886.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@57886.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(15)) sr ( // @[RetimeShiftRegister.scala 15:20:@57886.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@57899.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@57898.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@57897.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@57896.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@57895.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@57893.4]
endmodule
module RetimeWrapper_664( // @[:@58009.2]
  input   clock, // @[:@58010.4]
  input   reset, // @[:@58011.4]
  input   io_in, // @[:@58012.4]
  output  io_out // @[:@58012.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@58014.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@58014.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@58014.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@58014.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@58014.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@58014.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(14)) sr ( // @[RetimeShiftRegister.scala 15:20:@58014.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@58027.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@58026.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@58025.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@58024.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@58023.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@58021.4]
endmodule
module x639_inr_Foreach_sm( // @[:@58029.2]
  input   clock, // @[:@58030.4]
  input   reset, // @[:@58031.4]
  input   io_enable, // @[:@58032.4]
  output  io_done, // @[:@58032.4]
  input   io_rst, // @[:@58032.4]
  input   io_ctrDone, // @[:@58032.4]
  output  io_datapathEn, // @[:@58032.4]
  output  io_ctrInc, // @[:@58032.4]
  output  io_ctrRst, // @[:@58032.4]
  input   io_parentAck, // @[:@58032.4]
  input   io_backpressure, // @[:@58032.4]
  input   io_break // @[:@58032.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@58034.4]
  wire  active_reset; // @[Controllers.scala 261:22:@58034.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@58034.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@58034.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@58034.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@58034.4]
  wire  done_clock; // @[Controllers.scala 262:20:@58037.4]
  wire  done_reset; // @[Controllers.scala 262:20:@58037.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@58037.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@58037.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@58037.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@58037.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@58071.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@58071.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@58071.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@58071.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@58093.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@58093.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@58093.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@58093.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@58105.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@58105.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@58105.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@58105.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@58105.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@58113.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@58113.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@58113.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@58113.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@58113.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@58129.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@58129.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@58129.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@58129.4]
  wire  _T_80; // @[Controllers.scala 264:48:@58042.4]
  wire  _T_81; // @[Controllers.scala 264:46:@58043.4]
  wire  _T_82; // @[Controllers.scala 264:62:@58044.4]
  wire  _T_100; // @[package.scala 100:49:@58062.4]
  reg  _T_103; // @[package.scala 48:56:@58063.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@58076.4 package.scala 96:25:@58077.4]
  wire  _T_110; // @[package.scala 100:49:@58078.4]
  reg  _T_113; // @[package.scala 48:56:@58079.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@58081.4]
  wire  _T_118; // @[Controllers.scala 283:41:@58086.4]
  wire  _T_124; // @[package.scala 96:25:@58098.4 package.scala 96:25:@58099.4]
  wire  _T_126; // @[package.scala 100:49:@58100.4]
  reg  _T_129; // @[package.scala 48:56:@58101.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@58125.4]
  reg  _T_153; // @[package.scala 48:56:@58126.4]
  reg [31:0] _RAND_3;
  SRFF active ( // @[Controllers.scala 261:22:@58034.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@58037.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_660 RetimeWrapper ( // @[package.scala 93:22:@58071.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_660 RetimeWrapper_1 ( // @[package.scala 93:22:@58093.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@58105.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@58113.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_664 RetimeWrapper_4 ( // @[package.scala 93:22:@58129.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@58042.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@58043.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@58044.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@58062.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@58076.4 package.scala 96:25:@58077.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@58078.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@58081.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@58086.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@58098.4 package.scala 96:25:@58099.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@58100.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@58125.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@58104.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@58089.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@58092.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@58084.4]
  assign active_clock = clock; // @[:@58035.4]
  assign active_reset = reset; // @[:@58036.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@58047.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@58051.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@58052.4]
  assign done_clock = clock; // @[:@58038.4]
  assign done_reset = reset; // @[:@58039.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@58067.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@58060.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@58061.4]
  assign RetimeWrapper_clock = clock; // @[:@58072.4]
  assign RetimeWrapper_reset = reset; // @[:@58073.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@58074.4]
  assign RetimeWrapper_1_clock = clock; // @[:@58094.4]
  assign RetimeWrapper_1_reset = reset; // @[:@58095.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@58096.4]
  assign RetimeWrapper_2_clock = clock; // @[:@58106.4]
  assign RetimeWrapper_2_reset = reset; // @[:@58107.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@58109.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@58108.4]
  assign RetimeWrapper_3_clock = clock; // @[:@58114.4]
  assign RetimeWrapper_3_reset = reset; // @[:@58115.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@58117.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@58116.4]
  assign RetimeWrapper_4_clock = clock; // @[:@58130.4]
  assign RetimeWrapper_4_reset = reset; // @[:@58131.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@58132.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x639_inr_Foreach_iiCtr( // @[:@58142.2]
  input   clock, // @[:@58143.4]
  input   reset, // @[:@58144.4]
  input   io_input_enable, // @[:@58145.4]
  input   io_input_reset, // @[:@58145.4]
  output  io_output_issue, // @[:@58145.4]
  output  io_output_done // @[:@58145.4]
);
  reg [5:0] _T_15; // @[Counter.scala 135:22:@58147.4]
  reg [31:0] _RAND_0;
  wire  _T_17; // @[Counter.scala 138:24:@58148.4]
  wire  _T_20; // @[Counter.scala 139:23:@58150.4]
  wire [6:0] _T_26; // @[Counter.scala 141:68:@58153.4]
  wire [5:0] _T_27; // @[Counter.scala 141:68:@58154.4]
  wire [5:0] _T_28; // @[Counter.scala 141:68:@58155.4]
  wire [5:0] _T_29; // @[Counter.scala 141:23:@58156.4]
  wire [5:0] _T_30; // @[Counter.scala 142:19:@58157.4]
  wire [5:0] _T_32; // @[Counter.scala 143:15:@58158.4]
  assign _T_17 = $signed(_T_15) == $signed(6'she); // @[Counter.scala 138:24:@58148.4]
  assign _T_20 = $signed(_T_15) == $signed(6'sh0); // @[Counter.scala 139:23:@58150.4]
  assign _T_26 = $signed(_T_15) - $signed(6'sh1); // @[Counter.scala 141:68:@58153.4]
  assign _T_27 = $signed(_T_15) - $signed(6'sh1); // @[Counter.scala 141:68:@58154.4]
  assign _T_28 = $signed(_T_27); // @[Counter.scala 141:68:@58155.4]
  assign _T_29 = _T_20 ? $signed(6'she) : $signed(_T_28); // @[Counter.scala 141:23:@58156.4]
  assign _T_30 = io_input_enable ? $signed(_T_29) : $signed(_T_15); // @[Counter.scala 142:19:@58157.4]
  assign _T_32 = io_input_reset ? $signed(6'she) : $signed(_T_30); // @[Counter.scala 143:15:@58158.4]
  assign io_output_issue = _T_17 & io_input_enable; // @[Counter.scala 146:21:@58161.4]
  assign io_output_done = _T_20 & io_input_enable; // @[Counter.scala 145:20:@58160.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 6'she;
    end else begin
      if (io_input_reset) begin
        _T_15 <= 6'she;
      end else begin
        if (io_input_enable) begin
          if (_T_20) begin
            _T_15 <= 6'she;
          end else begin
            _T_15 <= _T_28;
          end
        end
      end
    end
  end
endmodule
module RetimeWrapper_676( // @[:@58769.2]
  input         clock, // @[:@58770.4]
  input         reset, // @[:@58771.4]
  input  [31:0] io_in, // @[:@58772.4]
  output [31:0] io_out // @[:@58772.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@58774.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@58774.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@58774.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@58774.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@58774.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@58774.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(14)) sr ( // @[RetimeShiftRegister.scala 15:20:@58774.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@58787.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@58786.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@58785.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@58784.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@58783.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@58781.4]
endmodule
module x639_inr_Foreach_kernelx639_inr_Foreach_concrete1( // @[:@59205.2]
  input         clock, // @[:@59206.4]
  input         reset, // @[:@59207.4]
  output [1:0]  io_in_x555_tmp_1_wPort_1_ofs_0, // @[:@59208.4]
  output [31:0] io_in_x555_tmp_1_wPort_1_data_0, // @[:@59208.4]
  output        io_in_x555_tmp_1_wPort_1_en_0, // @[:@59208.4]
  output        io_in_x555_tmp_1_sEn_5, // @[:@59208.4]
  output        io_in_x555_tmp_1_sDone_5, // @[:@59208.4]
  output [1:0]  io_in_x554_tmp_0_wPort_1_ofs_0, // @[:@59208.4]
  output [31:0] io_in_x554_tmp_0_wPort_1_data_0, // @[:@59208.4]
  output        io_in_x554_tmp_0_wPort_1_en_0, // @[:@59208.4]
  output        io_in_x554_tmp_0_sEn_5, // @[:@59208.4]
  output        io_in_x554_tmp_0_sDone_5, // @[:@59208.4]
  output [1:0]  io_in_x558_tmp_4_wPort_1_ofs_0, // @[:@59208.4]
  output [31:0] io_in_x558_tmp_4_wPort_1_data_0, // @[:@59208.4]
  output        io_in_x558_tmp_4_wPort_1_en_0, // @[:@59208.4]
  output        io_in_x558_tmp_4_sEn_5, // @[:@59208.4]
  output        io_in_x558_tmp_4_sDone_5, // @[:@59208.4]
  input         io_in_b552, // @[:@59208.4]
  output        io_in_x594_force_0_rPort_0_en_0, // @[:@59208.4]
  input  [31:0] io_in_x594_force_0_rPort_0_output_0, // @[:@59208.4]
  output        io_in_x594_force_0_sEn_1, // @[:@59208.4]
  output        io_in_x594_force_0_sDone_1, // @[:@59208.4]
  output [1:0]  io_in_x557_tmp_3_rPort_0_ofs_0, // @[:@59208.4]
  output        io_in_x557_tmp_3_rPort_0_en_0, // @[:@59208.4]
  input  [31:0] io_in_x557_tmp_3_rPort_0_output_0, // @[:@59208.4]
  output [1:0]  io_in_x557_tmp_3_wPort_1_ofs_0, // @[:@59208.4]
  output [31:0] io_in_x557_tmp_3_wPort_1_data_0, // @[:@59208.4]
  output        io_in_x557_tmp_3_wPort_1_en_0, // @[:@59208.4]
  output        io_in_x557_tmp_3_sEn_5, // @[:@59208.4]
  output        io_in_x557_tmp_3_sDone_5, // @[:@59208.4]
  output [1:0]  io_in_x556_tmp_2_wPort_1_ofs_0, // @[:@59208.4]
  output [31:0] io_in_x556_tmp_2_wPort_1_data_0, // @[:@59208.4]
  output        io_in_x556_tmp_2_wPort_1_en_0, // @[:@59208.4]
  output        io_in_x556_tmp_2_sEn_5, // @[:@59208.4]
  output        io_in_x556_tmp_2_sDone_5, // @[:@59208.4]
  input         io_in_b543, // @[:@59208.4]
  input         io_sigsIn_done, // @[:@59208.4]
  input         io_sigsIn_iiIssue, // @[:@59208.4]
  input         io_sigsIn_datapathEn, // @[:@59208.4]
  input         io_sigsIn_baseEn, // @[:@59208.4]
  input         io_sigsIn_break, // @[:@59208.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@59208.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@59208.4]
  input         io_rr // @[:@59208.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@59465.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@59465.4]
  wire  x630_mul_1_clock; // @[Math.scala 262:24:@59499.4]
  wire  x630_mul_1_reset; // @[Math.scala 262:24:@59499.4]
  wire [31:0] x630_mul_1_io_a; // @[Math.scala 262:24:@59499.4]
  wire [31:0] x630_mul_1_io_b; // @[Math.scala 262:24:@59499.4]
  wire  x630_mul_1_io_flow; // @[Math.scala 262:24:@59499.4]
  wire [31:0] x630_mul_1_io_result; // @[Math.scala 262:24:@59499.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@59534.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@59534.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@59534.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@59534.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@59534.4]
  wire  x633_mul_1_clock; // @[Math.scala 262:24:@59543.4]
  wire  x633_mul_1_reset; // @[Math.scala 262:24:@59543.4]
  wire [31:0] x633_mul_1_io_a; // @[Math.scala 262:24:@59543.4]
  wire [31:0] x633_mul_1_io_b; // @[Math.scala 262:24:@59543.4]
  wire  x633_mul_1_io_flow; // @[Math.scala 262:24:@59543.4]
  wire [31:0] x633_mul_1_io_result; // @[Math.scala 262:24:@59543.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@59554.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@59554.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@59554.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@59554.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@59564.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@59564.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@59564.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@59564.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@59574.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@59574.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@59574.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@59574.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@59584.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@59584.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@59584.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@59584.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@59598.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@59598.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@59598.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@59598.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@59624.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@59624.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@59624.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@59624.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@59650.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@59650.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@59650.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@59650.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@59676.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@59676.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@59676.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@59676.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@59702.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@59702.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@59702.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@59702.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@59723.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@59723.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@59723.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@59723.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@59723.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@59734.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@59734.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@59734.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@59734.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@59734.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@59745.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@59745.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@59745.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@59745.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@59745.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@59756.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@59756.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@59756.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@59756.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@59756.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@59767.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@59767.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@59767.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@59767.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@59767.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@59778.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@59778.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@59778.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@59778.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@59778.4]
  wire  b627; // @[sm_x639_inr_Foreach.scala 86:18:@59473.4]
  wire  _T_1782; // @[sm_x639_inr_Foreach.scala 91:114:@59479.4]
  wire  _T_1783; // @[sm_x639_inr_Foreach.scala 91:111:@59480.4]
  wire  _T_1784; // @[sm_x639_inr_Foreach.scala 91:156:@59481.4]
  wire  _T_1788; // @[implicits.scala 56:10:@59483.4]
  wire  _T_1789; // @[sm_x639_inr_Foreach.scala 91:131:@59484.4]
  wire  _T_1790; // @[sm_x639_inr_Foreach.scala 91:228:@59485.4]
  wire  _T_1791; // @[sm_x639_inr_Foreach.scala 91:236:@59486.4]
  wire  _T_1871; // @[package.scala 96:25:@59603.4 package.scala 96:25:@59604.4]
  wire  _T_1873; // @[implicits.scala 56:10:@59605.4]
  wire  _T_1874; // @[sm_x639_inr_Foreach.scala 123:115:@59606.4]
  wire  _T_1876; // @[sm_x639_inr_Foreach.scala 123:213:@59608.4]
  wire  x787_b627_D14; // @[package.scala 96:25:@59579.4 package.scala 96:25:@59580.4]
  wire  _T_1878; // @[sm_x639_inr_Foreach.scala 123:258:@59610.4]
  wire  x785_b552_D14; // @[package.scala 96:25:@59559.4 package.scala 96:25:@59560.4]
  wire  _T_1879; // @[sm_x639_inr_Foreach.scala 123:266:@59611.4]
  wire  x788_b543_D14; // @[package.scala 96:25:@59589.4 package.scala 96:25:@59590.4]
  wire  _T_1891; // @[package.scala 96:25:@59629.4 package.scala 96:25:@59630.4]
  wire  _T_1893; // @[implicits.scala 56:10:@59631.4]
  wire  _T_1894; // @[sm_x639_inr_Foreach.scala 128:115:@59632.4]
  wire  _T_1896; // @[sm_x639_inr_Foreach.scala 128:213:@59634.4]
  wire  _T_1898; // @[sm_x639_inr_Foreach.scala 128:258:@59636.4]
  wire  _T_1899; // @[sm_x639_inr_Foreach.scala 128:266:@59637.4]
  wire  _T_1911; // @[package.scala 96:25:@59655.4 package.scala 96:25:@59656.4]
  wire  _T_1913; // @[implicits.scala 56:10:@59657.4]
  wire  _T_1914; // @[sm_x639_inr_Foreach.scala 133:115:@59658.4]
  wire  _T_1916; // @[sm_x639_inr_Foreach.scala 133:213:@59660.4]
  wire  _T_1918; // @[sm_x639_inr_Foreach.scala 133:258:@59662.4]
  wire  _T_1919; // @[sm_x639_inr_Foreach.scala 133:266:@59663.4]
  wire  _T_1931; // @[package.scala 96:25:@59681.4 package.scala 96:25:@59682.4]
  wire  _T_1933; // @[implicits.scala 56:10:@59683.4]
  wire  _T_1934; // @[sm_x639_inr_Foreach.scala 138:115:@59684.4]
  wire  _T_1936; // @[sm_x639_inr_Foreach.scala 138:213:@59686.4]
  wire  _T_1938; // @[sm_x639_inr_Foreach.scala 138:258:@59688.4]
  wire  _T_1939; // @[sm_x639_inr_Foreach.scala 138:266:@59689.4]
  wire  _T_1951; // @[package.scala 96:25:@59707.4 package.scala 96:25:@59708.4]
  wire  _T_1953; // @[implicits.scala 56:10:@59709.4]
  wire  _T_1954; // @[sm_x639_inr_Foreach.scala 143:115:@59710.4]
  wire  _T_1956; // @[sm_x639_inr_Foreach.scala 143:213:@59712.4]
  wire  _T_1958; // @[sm_x639_inr_Foreach.scala 143:258:@59714.4]
  wire  _T_1959; // @[sm_x639_inr_Foreach.scala 143:266:@59715.4]
  wire  _T_1964; // @[package.scala 96:25:@59728.4 package.scala 96:25:@59729.4]
  wire  _T_1970; // @[package.scala 96:25:@59739.4 package.scala 96:25:@59740.4]
  wire  _T_1976; // @[package.scala 96:25:@59750.4 package.scala 96:25:@59751.4]
  wire  _T_1982; // @[package.scala 96:25:@59761.4 package.scala 96:25:@59762.4]
  wire  _T_1988; // @[package.scala 96:25:@59772.4 package.scala 96:25:@59773.4]
  wire  _T_1994; // @[package.scala 96:25:@59783.4 package.scala 96:25:@59784.4]
  wire [31:0] b626_number; // @[Math.scala 723:22:@59470.4 Math.scala 724:14:@59471.4]
  wire [31:0] x786_b626_D14_number; // @[package.scala 96:25:@59569.4 package.scala 96:25:@59570.4]
  _ _ ( // @[Math.scala 720:24:@59465.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x586_mul x630_mul_1 ( // @[Math.scala 262:24:@59499.4]
    .clock(x630_mul_1_clock),
    .reset(x630_mul_1_reset),
    .io_a(x630_mul_1_io_a),
    .io_b(x630_mul_1_io_b),
    .io_flow(x630_mul_1_io_flow),
    .io_result(x630_mul_1_io_result)
  );
  RetimeWrapper_527 RetimeWrapper ( // @[package.scala 93:22:@59534.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x586_mul x633_mul_1 ( // @[Math.scala 262:24:@59543.4]
    .clock(x633_mul_1_clock),
    .reset(x633_mul_1_reset),
    .io_a(x633_mul_1_io_a),
    .io_b(x633_mul_1_io_b),
    .io_flow(x633_mul_1_io_flow),
    .io_result(x633_mul_1_io_result)
  );
  RetimeWrapper_664 RetimeWrapper_1 ( // @[package.scala 93:22:@59554.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_676 RetimeWrapper_2 ( // @[package.scala 93:22:@59564.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_664 RetimeWrapper_3 ( // @[package.scala 93:22:@59574.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_664 RetimeWrapper_4 ( // @[package.scala 93:22:@59584.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_664 RetimeWrapper_5 ( // @[package.scala 93:22:@59598.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_664 RetimeWrapper_6 ( // @[package.scala 93:22:@59624.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_664 RetimeWrapper_7 ( // @[package.scala 93:22:@59650.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_664 RetimeWrapper_8 ( // @[package.scala 93:22:@59676.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_664 RetimeWrapper_9 ( // @[package.scala 93:22:@59702.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@59723.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 ( // @[package.scala 93:22:@59734.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper RetimeWrapper_12 ( // @[package.scala 93:22:@59745.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 ( // @[package.scala 93:22:@59756.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@59767.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@59778.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  assign b627 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x639_inr_Foreach.scala 86:18:@59473.4]
  assign _T_1782 = ~ io_sigsIn_break; // @[sm_x639_inr_Foreach.scala 91:114:@59479.4]
  assign _T_1783 = io_rr & _T_1782; // @[sm_x639_inr_Foreach.scala 91:111:@59480.4]
  assign _T_1784 = io_sigsIn_datapathEn & io_sigsIn_iiIssue; // @[sm_x639_inr_Foreach.scala 91:156:@59481.4]
  assign _T_1788 = io_rr ? _T_1784 : 1'h0; // @[implicits.scala 56:10:@59483.4]
  assign _T_1789 = _T_1783 & _T_1788; // @[sm_x639_inr_Foreach.scala 91:131:@59484.4]
  assign _T_1790 = _T_1789 & b627; // @[sm_x639_inr_Foreach.scala 91:228:@59485.4]
  assign _T_1791 = _T_1790 & io_in_b552; // @[sm_x639_inr_Foreach.scala 91:236:@59486.4]
  assign _T_1871 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@59603.4 package.scala 96:25:@59604.4]
  assign _T_1873 = io_rr ? _T_1871 : 1'h0; // @[implicits.scala 56:10:@59605.4]
  assign _T_1874 = _T_1782 & _T_1873; // @[sm_x639_inr_Foreach.scala 123:115:@59606.4]
  assign _T_1876 = _T_1874 & _T_1782; // @[sm_x639_inr_Foreach.scala 123:213:@59608.4]
  assign x787_b627_D14 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@59579.4 package.scala 96:25:@59580.4]
  assign _T_1878 = _T_1876 & x787_b627_D14; // @[sm_x639_inr_Foreach.scala 123:258:@59610.4]
  assign x785_b552_D14 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@59559.4 package.scala 96:25:@59560.4]
  assign _T_1879 = _T_1878 & x785_b552_D14; // @[sm_x639_inr_Foreach.scala 123:266:@59611.4]
  assign x788_b543_D14 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@59589.4 package.scala 96:25:@59590.4]
  assign _T_1891 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@59629.4 package.scala 96:25:@59630.4]
  assign _T_1893 = io_rr ? _T_1891 : 1'h0; // @[implicits.scala 56:10:@59631.4]
  assign _T_1894 = _T_1782 & _T_1893; // @[sm_x639_inr_Foreach.scala 128:115:@59632.4]
  assign _T_1896 = _T_1894 & _T_1782; // @[sm_x639_inr_Foreach.scala 128:213:@59634.4]
  assign _T_1898 = _T_1896 & x787_b627_D14; // @[sm_x639_inr_Foreach.scala 128:258:@59636.4]
  assign _T_1899 = _T_1898 & x785_b552_D14; // @[sm_x639_inr_Foreach.scala 128:266:@59637.4]
  assign _T_1911 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@59655.4 package.scala 96:25:@59656.4]
  assign _T_1913 = io_rr ? _T_1911 : 1'h0; // @[implicits.scala 56:10:@59657.4]
  assign _T_1914 = _T_1782 & _T_1913; // @[sm_x639_inr_Foreach.scala 133:115:@59658.4]
  assign _T_1916 = _T_1914 & _T_1782; // @[sm_x639_inr_Foreach.scala 133:213:@59660.4]
  assign _T_1918 = _T_1916 & x787_b627_D14; // @[sm_x639_inr_Foreach.scala 133:258:@59662.4]
  assign _T_1919 = _T_1918 & x785_b552_D14; // @[sm_x639_inr_Foreach.scala 133:266:@59663.4]
  assign _T_1931 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@59681.4 package.scala 96:25:@59682.4]
  assign _T_1933 = io_rr ? _T_1931 : 1'h0; // @[implicits.scala 56:10:@59683.4]
  assign _T_1934 = _T_1782 & _T_1933; // @[sm_x639_inr_Foreach.scala 138:115:@59684.4]
  assign _T_1936 = _T_1934 & _T_1782; // @[sm_x639_inr_Foreach.scala 138:213:@59686.4]
  assign _T_1938 = _T_1936 & x787_b627_D14; // @[sm_x639_inr_Foreach.scala 138:258:@59688.4]
  assign _T_1939 = _T_1938 & x785_b552_D14; // @[sm_x639_inr_Foreach.scala 138:266:@59689.4]
  assign _T_1951 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@59707.4 package.scala 96:25:@59708.4]
  assign _T_1953 = io_rr ? _T_1951 : 1'h0; // @[implicits.scala 56:10:@59709.4]
  assign _T_1954 = _T_1782 & _T_1953; // @[sm_x639_inr_Foreach.scala 143:115:@59710.4]
  assign _T_1956 = _T_1954 & _T_1782; // @[sm_x639_inr_Foreach.scala 143:213:@59712.4]
  assign _T_1958 = _T_1956 & x787_b627_D14; // @[sm_x639_inr_Foreach.scala 143:258:@59714.4]
  assign _T_1959 = _T_1958 & x785_b552_D14; // @[sm_x639_inr_Foreach.scala 143:266:@59715.4]
  assign _T_1964 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@59728.4 package.scala 96:25:@59729.4]
  assign _T_1970 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@59739.4 package.scala 96:25:@59740.4]
  assign _T_1976 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@59750.4 package.scala 96:25:@59751.4]
  assign _T_1982 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@59761.4 package.scala 96:25:@59762.4]
  assign _T_1988 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@59772.4 package.scala 96:25:@59773.4]
  assign _T_1994 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@59783.4 package.scala 96:25:@59784.4]
  assign b626_number = __io_result; // @[Math.scala 723:22:@59470.4 Math.scala 724:14:@59471.4]
  assign x786_b626_D14_number = RetimeWrapper_2_io_out; // @[package.scala 96:25:@59569.4 package.scala 96:25:@59570.4]
  assign io_in_x555_tmp_1_wPort_1_ofs_0 = x786_b626_D14_number[1:0]; // @[MemInterfaceType.scala 89:54:@59614.4]
  assign io_in_x555_tmp_1_wPort_1_data_0 = x633_mul_1_io_result; // @[MemInterfaceType.scala 90:56:@59615.4]
  assign io_in_x555_tmp_1_wPort_1_en_0 = _T_1879 & x788_b543_D14; // @[MemInterfaceType.scala 93:57:@59617.4]
  assign io_in_x555_tmp_1_sEn_5 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@59742.4]
  assign io_in_x555_tmp_1_sDone_5 = io_rr ? _T_1970 : 1'h0; // @[MemInterfaceType.scala 197:17:@59743.4]
  assign io_in_x554_tmp_0_wPort_1_ofs_0 = x786_b626_D14_number[1:0]; // @[MemInterfaceType.scala 89:54:@59640.4]
  assign io_in_x554_tmp_0_wPort_1_data_0 = x633_mul_1_io_result; // @[MemInterfaceType.scala 90:56:@59641.4]
  assign io_in_x554_tmp_0_wPort_1_en_0 = _T_1899 & x788_b543_D14; // @[MemInterfaceType.scala 93:57:@59643.4]
  assign io_in_x554_tmp_0_sEn_5 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@59731.4]
  assign io_in_x554_tmp_0_sDone_5 = io_rr ? _T_1964 : 1'h0; // @[MemInterfaceType.scala 197:17:@59732.4]
  assign io_in_x558_tmp_4_wPort_1_ofs_0 = x786_b626_D14_number[1:0]; // @[MemInterfaceType.scala 89:54:@59666.4]
  assign io_in_x558_tmp_4_wPort_1_data_0 = x633_mul_1_io_result; // @[MemInterfaceType.scala 90:56:@59667.4]
  assign io_in_x558_tmp_4_wPort_1_en_0 = _T_1919 & x788_b543_D14; // @[MemInterfaceType.scala 93:57:@59669.4]
  assign io_in_x558_tmp_4_sEn_5 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@59775.4]
  assign io_in_x558_tmp_4_sDone_5 = io_rr ? _T_1988 : 1'h0; // @[MemInterfaceType.scala 197:17:@59776.4]
  assign io_in_x594_force_0_rPort_0_en_0 = _T_1791 & io_in_b543; // @[MemInterfaceType.scala 110:79:@59528.4]
  assign io_in_x594_force_0_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@59786.4]
  assign io_in_x594_force_0_sDone_1 = io_rr ? _T_1994 : 1'h0; // @[MemInterfaceType.scala 197:17:@59787.4]
  assign io_in_x557_tmp_3_rPort_0_ofs_0 = b626_number[1:0]; // @[MemInterfaceType.scala 107:54:@59490.4]
  assign io_in_x557_tmp_3_rPort_0_en_0 = _T_1791 & io_in_b543; // @[MemInterfaceType.scala 110:79:@59492.4]
  assign io_in_x557_tmp_3_wPort_1_ofs_0 = x786_b626_D14_number[1:0]; // @[MemInterfaceType.scala 89:54:@59692.4]
  assign io_in_x557_tmp_3_wPort_1_data_0 = x633_mul_1_io_result; // @[MemInterfaceType.scala 90:56:@59693.4]
  assign io_in_x557_tmp_3_wPort_1_en_0 = _T_1939 & x788_b543_D14; // @[MemInterfaceType.scala 93:57:@59695.4]
  assign io_in_x557_tmp_3_sEn_5 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@59764.4]
  assign io_in_x557_tmp_3_sDone_5 = io_rr ? _T_1982 : 1'h0; // @[MemInterfaceType.scala 197:17:@59765.4]
  assign io_in_x556_tmp_2_wPort_1_ofs_0 = x786_b626_D14_number[1:0]; // @[MemInterfaceType.scala 89:54:@59718.4]
  assign io_in_x556_tmp_2_wPort_1_data_0 = x633_mul_1_io_result; // @[MemInterfaceType.scala 90:56:@59719.4]
  assign io_in_x556_tmp_2_wPort_1_en_0 = _T_1959 & x788_b543_D14; // @[MemInterfaceType.scala 93:57:@59721.4]
  assign io_in_x556_tmp_2_sEn_5 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@59753.4]
  assign io_in_x556_tmp_2_sDone_5 = io_rr ? _T_1976 : 1'h0; // @[MemInterfaceType.scala 197:17:@59754.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@59468.4]
  assign x630_mul_1_clock = clock; // @[:@59500.4]
  assign x630_mul_1_reset = reset; // @[:@59501.4]
  assign x630_mul_1_io_a = io_in_x557_tmp_3_rPort_0_output_0; // @[Math.scala 263:17:@59502.4]
  assign x630_mul_1_io_b = 32'h66666; // @[Math.scala 264:17:@59503.4]
  assign x630_mul_1_io_flow = 1'h1; // @[Math.scala 265:20:@59504.4]
  assign RetimeWrapper_clock = clock; // @[:@59535.4]
  assign RetimeWrapper_reset = reset; // @[:@59536.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@59538.4]
  assign RetimeWrapper_io_in = io_in_x594_force_0_rPort_0_output_0; // @[package.scala 94:16:@59537.4]
  assign x633_mul_1_clock = clock; // @[:@59544.4]
  assign x633_mul_1_reset = reset; // @[:@59545.4]
  assign x633_mul_1_io_a = x630_mul_1_io_result; // @[Math.scala 263:17:@59546.4]
  assign x633_mul_1_io_b = RetimeWrapper_io_out; // @[Math.scala 264:17:@59547.4]
  assign x633_mul_1_io_flow = 1'h1; // @[Math.scala 265:20:@59548.4]
  assign RetimeWrapper_1_clock = clock; // @[:@59555.4]
  assign RetimeWrapper_1_reset = reset; // @[:@59556.4]
  assign RetimeWrapper_1_io_in = io_in_b552; // @[package.scala 94:16:@59557.4]
  assign RetimeWrapper_2_clock = clock; // @[:@59565.4]
  assign RetimeWrapper_2_reset = reset; // @[:@59566.4]
  assign RetimeWrapper_2_io_in = __io_result; // @[package.scala 94:16:@59567.4]
  assign RetimeWrapper_3_clock = clock; // @[:@59575.4]
  assign RetimeWrapper_3_reset = reset; // @[:@59576.4]
  assign RetimeWrapper_3_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@59577.4]
  assign RetimeWrapper_4_clock = clock; // @[:@59585.4]
  assign RetimeWrapper_4_reset = reset; // @[:@59586.4]
  assign RetimeWrapper_4_io_in = io_in_b543; // @[package.scala 94:16:@59587.4]
  assign RetimeWrapper_5_clock = clock; // @[:@59599.4]
  assign RetimeWrapper_5_reset = reset; // @[:@59600.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_datapathEn & io_sigsIn_iiIssue; // @[package.scala 94:16:@59601.4]
  assign RetimeWrapper_6_clock = clock; // @[:@59625.4]
  assign RetimeWrapper_6_reset = reset; // @[:@59626.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn & io_sigsIn_iiIssue; // @[package.scala 94:16:@59627.4]
  assign RetimeWrapper_7_clock = clock; // @[:@59651.4]
  assign RetimeWrapper_7_reset = reset; // @[:@59652.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_datapathEn & io_sigsIn_iiIssue; // @[package.scala 94:16:@59653.4]
  assign RetimeWrapper_8_clock = clock; // @[:@59677.4]
  assign RetimeWrapper_8_reset = reset; // @[:@59678.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_datapathEn & io_sigsIn_iiIssue; // @[package.scala 94:16:@59679.4]
  assign RetimeWrapper_9_clock = clock; // @[:@59703.4]
  assign RetimeWrapper_9_reset = reset; // @[:@59704.4]
  assign RetimeWrapper_9_io_in = io_sigsIn_datapathEn & io_sigsIn_iiIssue; // @[package.scala 94:16:@59705.4]
  assign RetimeWrapper_10_clock = clock; // @[:@59724.4]
  assign RetimeWrapper_10_reset = reset; // @[:@59725.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@59727.4]
  assign RetimeWrapper_10_io_in = io_sigsIn_done; // @[package.scala 94:16:@59726.4]
  assign RetimeWrapper_11_clock = clock; // @[:@59735.4]
  assign RetimeWrapper_11_reset = reset; // @[:@59736.4]
  assign RetimeWrapper_11_io_flow = 1'h1; // @[package.scala 95:18:@59738.4]
  assign RetimeWrapper_11_io_in = io_sigsIn_done; // @[package.scala 94:16:@59737.4]
  assign RetimeWrapper_12_clock = clock; // @[:@59746.4]
  assign RetimeWrapper_12_reset = reset; // @[:@59747.4]
  assign RetimeWrapper_12_io_flow = 1'h1; // @[package.scala 95:18:@59749.4]
  assign RetimeWrapper_12_io_in = io_sigsIn_done; // @[package.scala 94:16:@59748.4]
  assign RetimeWrapper_13_clock = clock; // @[:@59757.4]
  assign RetimeWrapper_13_reset = reset; // @[:@59758.4]
  assign RetimeWrapper_13_io_flow = 1'h1; // @[package.scala 95:18:@59760.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_done; // @[package.scala 94:16:@59759.4]
  assign RetimeWrapper_14_clock = clock; // @[:@59768.4]
  assign RetimeWrapper_14_reset = reset; // @[:@59769.4]
  assign RetimeWrapper_14_io_flow = 1'h1; // @[package.scala 95:18:@59771.4]
  assign RetimeWrapper_14_io_in = io_sigsIn_done; // @[package.scala 94:16:@59770.4]
  assign RetimeWrapper_15_clock = clock; // @[:@59779.4]
  assign RetimeWrapper_15_reset = reset; // @[:@59780.4]
  assign RetimeWrapper_15_io_flow = 1'h1; // @[package.scala 95:18:@59782.4]
  assign RetimeWrapper_15_io_in = io_sigsIn_done; // @[package.scala 94:16:@59781.4]
endmodule
module x652_inr_Foreach_sm( // @[:@59975.2]
  input   clock, // @[:@59976.4]
  input   reset, // @[:@59977.4]
  input   io_enable, // @[:@59978.4]
  output  io_done, // @[:@59978.4]
  output  io_doneLatch, // @[:@59978.4]
  input   io_ctrDone, // @[:@59978.4]
  output  io_datapathEn, // @[:@59978.4]
  output  io_ctrInc, // @[:@59978.4]
  output  io_ctrRst, // @[:@59978.4]
  input   io_parentAck, // @[:@59978.4]
  input   io_backpressure, // @[:@59978.4]
  input   io_break // @[:@59978.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@59980.4]
  wire  active_reset; // @[Controllers.scala 261:22:@59980.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@59980.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@59980.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@59980.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@59980.4]
  wire  done_clock; // @[Controllers.scala 262:20:@59983.4]
  wire  done_reset; // @[Controllers.scala 262:20:@59983.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@59983.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@59983.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@59983.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@59983.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@60017.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@60017.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@60017.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@60017.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@60017.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@60039.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@60039.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@60039.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@60039.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@60039.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@60051.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@60051.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@60051.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@60051.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@60051.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@60059.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@60059.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@60059.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@60059.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@60059.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@60075.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@60075.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@60075.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@60075.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@60075.4]
  wire  _T_80; // @[Controllers.scala 264:48:@59988.4]
  wire  _T_81; // @[Controllers.scala 264:46:@59989.4]
  wire  _T_82; // @[Controllers.scala 264:62:@59990.4]
  wire  _T_83; // @[Controllers.scala 264:60:@59991.4]
  wire  _T_100; // @[package.scala 100:49:@60008.4]
  reg  _T_103; // @[package.scala 48:56:@60009.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@60022.4 package.scala 96:25:@60023.4]
  wire  _T_110; // @[package.scala 100:49:@60024.4]
  reg  _T_113; // @[package.scala 48:56:@60025.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@60027.4]
  wire  _T_118; // @[Controllers.scala 283:41:@60032.4]
  wire  _T_119; // @[Controllers.scala 283:59:@60033.4]
  wire  _T_121; // @[Controllers.scala 284:37:@60036.4]
  wire  _T_124; // @[package.scala 96:25:@60044.4 package.scala 96:25:@60045.4]
  wire  _T_126; // @[package.scala 100:49:@60046.4]
  reg  _T_129; // @[package.scala 48:56:@60047.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@60069.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@60071.4]
  reg  _T_153; // @[package.scala 48:56:@60072.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@60080.4 package.scala 96:25:@60081.4]
  wire  _T_158; // @[Controllers.scala 292:61:@60082.4]
  wire  _T_159; // @[Controllers.scala 292:24:@60083.4]
  SRFF active ( // @[Controllers.scala 261:22:@59980.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@59983.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_25 RetimeWrapper ( // @[package.scala 93:22:@60017.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@60039.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@60051.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@60059.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_58 RetimeWrapper_4 ( // @[package.scala 93:22:@60075.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@59988.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@59989.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@59990.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@59991.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@60008.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@60022.4 package.scala 96:25:@60023.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@60024.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@60027.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@60032.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@60033.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@60036.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@60044.4 package.scala 96:25:@60045.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@60046.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@60071.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@60080.4 package.scala 96:25:@60081.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@60082.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@60083.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@60050.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@60085.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@60035.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@60038.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@60030.4]
  assign active_clock = clock; // @[:@59981.4]
  assign active_reset = reset; // @[:@59982.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@59993.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@59997.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@59998.4]
  assign done_clock = clock; // @[:@59984.4]
  assign done_reset = reset; // @[:@59985.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@60013.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@60006.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@60007.4]
  assign RetimeWrapper_clock = clock; // @[:@60018.4]
  assign RetimeWrapper_reset = reset; // @[:@60019.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@60021.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@60020.4]
  assign RetimeWrapper_1_clock = clock; // @[:@60040.4]
  assign RetimeWrapper_1_reset = reset; // @[:@60041.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@60043.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@60042.4]
  assign RetimeWrapper_2_clock = clock; // @[:@60052.4]
  assign RetimeWrapper_2_reset = reset; // @[:@60053.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@60055.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@60054.4]
  assign RetimeWrapper_3_clock = clock; // @[:@60060.4]
  assign RetimeWrapper_3_reset = reset; // @[:@60061.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@60063.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@60062.4]
  assign RetimeWrapper_4_clock = clock; // @[:@60076.4]
  assign RetimeWrapper_4_reset = reset; // @[:@60077.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@60079.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@60078.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x648_sum( // @[:@60428.2]
  input         clock, // @[:@60429.4]
  input         reset, // @[:@60430.4]
  input  [31:0] io_a, // @[:@60431.4]
  input  [31:0] io_b, // @[:@60431.4]
  output [31:0] io_result // @[:@60431.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@60439.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@60439.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@60446.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@60446.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@60464.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@60464.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@60464.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@60464.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@60464.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@60444.4 Math.scala 724:14:@60445.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@60451.4 Math.scala 724:14:@60452.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@60453.4]
  __37 _ ( // @[Math.scala 720:24:@60439.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __37 __1 ( // @[Math.scala 720:24:@60446.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_52 fix2fixBox ( // @[Math.scala 141:30:@60464.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@60444.4 Math.scala 724:14:@60445.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@60451.4 Math.scala 724:14:@60452.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@60453.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@60472.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@60442.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@60449.4]
  assign fix2fixBox_clock = clock; // @[:@60465.4]
  assign fix2fixBox_reset = reset; // @[:@60466.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@60467.4]
  assign fix2fixBox_io_flow = 1'h1; // @[Math.scala 145:26:@60470.4]
endmodule
module RetimeWrapper_705( // @[:@60614.2]
  input         clock, // @[:@60615.4]
  input         reset, // @[:@60616.4]
  input  [31:0] io_in, // @[:@60617.4]
  output [31:0] io_out // @[:@60617.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@60619.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@60619.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@60619.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@60619.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@60619.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@60619.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@60619.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@60632.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@60631.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@60630.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@60629.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@60628.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@60626.4]
endmodule
module x652_inr_Foreach_kernelx652_inr_Foreach_concrete1( // @[:@60730.2]
  input         clock, // @[:@60731.4]
  input         reset, // @[:@60732.4]
  input  [31:0] io_in_b550_number, // @[:@60733.4]
  output [1:0]  io_in_x558_tmp_4_rPort_0_ofs_0, // @[:@60733.4]
  output        io_in_x558_tmp_4_rPort_0_en_0, // @[:@60733.4]
  input  [31:0] io_in_x558_tmp_4_rPort_0_output_0, // @[:@60733.4]
  output        io_in_x558_tmp_4_sEn_6, // @[:@60733.4]
  output        io_in_x558_tmp_4_sDone_6, // @[:@60733.4]
  output [1:0]  io_in_x545_accum_1_wPort_0_ofs_0, // @[:@60733.4]
  output [31:0] io_in_x545_accum_1_wPort_0_data_0, // @[:@60733.4]
  output        io_in_x545_accum_1_wPort_0_en_0, // @[:@60733.4]
  output [1:0]  io_in_x544_accum_0_rPort_0_ofs_0, // @[:@60733.4]
  output        io_in_x544_accum_0_rPort_0_en_0, // @[:@60733.4]
  input  [31:0] io_in_x544_accum_0_rPort_0_output_0, // @[:@60733.4]
  output [1:0]  io_in_x544_accum_0_wPort_0_ofs_0, // @[:@60733.4]
  output [31:0] io_in_x544_accum_0_wPort_0_data_0, // @[:@60733.4]
  output        io_in_x544_accum_0_wPort_0_en_0, // @[:@60733.4]
  input         io_in_b543, // @[:@60733.4]
  input         io_sigsIn_done, // @[:@60733.4]
  input         io_sigsIn_datapathEn, // @[:@60733.4]
  input         io_sigsIn_baseEn, // @[:@60733.4]
  input         io_sigsIn_break, // @[:@60733.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@60733.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@60733.4]
  input         io_rr // @[:@60733.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@60831.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@60831.4]
  wire  x648_sum_1_clock; // @[Math.scala 150:24:@60890.4]
  wire  x648_sum_1_reset; // @[Math.scala 150:24:@60890.4]
  wire [31:0] x648_sum_1_io_a; // @[Math.scala 150:24:@60890.4]
  wire [31:0] x648_sum_1_io_b; // @[Math.scala 150:24:@60890.4]
  wire [31:0] x648_sum_1_io_result; // @[Math.scala 150:24:@60890.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@60901.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@60901.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@60901.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@60901.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@60901.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@60911.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@60911.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@60911.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@60911.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@60911.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@60924.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@60924.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@60924.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@60924.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@60924.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@60934.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@60934.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@60934.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@60934.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@60934.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@60944.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@60944.4]
  wire [31:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@60944.4]
  wire [31:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@60944.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@60958.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@60958.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@60958.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@60958.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@60958.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@60983.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@60983.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@60983.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@60983.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@60983.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@61003.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@61003.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@61003.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@61003.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@61003.4]
  wire  b553; // @[sm_x652_inr_Foreach.scala 76:18:@60839.4]
  wire  _T_764; // @[sm_x652_inr_Foreach.scala 81:114:@60845.4]
  wire  _T_765; // @[sm_x652_inr_Foreach.scala 81:111:@60846.4]
  wire  _T_770; // @[implicits.scala 56:10:@60849.4]
  wire  _T_771; // @[sm_x652_inr_Foreach.scala 81:131:@60850.4]
  wire  _T_772; // @[sm_x652_inr_Foreach.scala 81:228:@60851.4]
  wire [31:0] _T_806; // @[Math.scala 510:37:@60885.4]
  wire  x790_x647_D3; // @[package.scala 96:25:@60916.4 package.scala 96:25:@60917.4]
  wire [31:0] x789_x641_elem_0_D1_number; // @[package.scala 96:25:@60906.4 package.scala 96:25:@60907.4]
  wire [31:0] x648_sum_number; // @[Math.scala 154:22:@60896.4 Math.scala 155:14:@60897.4]
  wire  _T_850; // @[package.scala 96:25:@60963.4 package.scala 96:25:@60964.4]
  wire  _T_852; // @[implicits.scala 56:10:@60965.4]
  wire  _T_853; // @[sm_x652_inr_Foreach.scala 115:117:@60966.4]
  wire  _T_855; // @[sm_x652_inr_Foreach.scala 115:214:@60968.4]
  wire  x792_b553_D3; // @[package.scala 96:25:@60939.4 package.scala 96:25:@60940.4]
  wire  _T_857; // @[sm_x652_inr_Foreach.scala 115:259:@60970.4]
  wire  x791_b543_D3; // @[package.scala 96:25:@60929.4 package.scala 96:25:@60930.4]
  wire  _T_869; // @[package.scala 96:25:@60988.4 package.scala 96:25:@60989.4]
  wire  _T_871; // @[implicits.scala 56:10:@60990.4]
  wire  _T_872; // @[sm_x652_inr_Foreach.scala 120:117:@60991.4]
  wire  _T_874; // @[sm_x652_inr_Foreach.scala 120:214:@60993.4]
  wire  _T_876; // @[sm_x652_inr_Foreach.scala 120:259:@60995.4]
  wire  _T_881; // @[package.scala 96:25:@61008.4 package.scala 96:25:@61009.4]
  wire [31:0] b551_number; // @[Math.scala 723:22:@60836.4 Math.scala 724:14:@60837.4]
  wire [31:0] x793_b551_D3_number; // @[package.scala 96:25:@60949.4 package.scala 96:25:@60950.4]
  _ _ ( // @[Math.scala 720:24:@60831.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x648_sum x648_sum_1 ( // @[Math.scala 150:24:@60890.4]
    .clock(x648_sum_1_clock),
    .reset(x648_sum_1_reset),
    .io_a(x648_sum_1_io_a),
    .io_b(x648_sum_1_io_b),
    .io_result(x648_sum_1_io_result)
  );
  RetimeWrapper_31 RetimeWrapper ( // @[package.scala 93:22:@60901.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_58 RetimeWrapper_1 ( // @[package.scala 93:22:@60911.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_58 RetimeWrapper_2 ( // @[package.scala 93:22:@60924.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_58 RetimeWrapper_3 ( // @[package.scala 93:22:@60934.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_705 RetimeWrapper_4 ( // @[package.scala 93:22:@60944.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_58 RetimeWrapper_5 ( // @[package.scala 93:22:@60958.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_58 RetimeWrapper_6 ( // @[package.scala 93:22:@60983.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@61003.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign b553 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x652_inr_Foreach.scala 76:18:@60839.4]
  assign _T_764 = ~ io_sigsIn_break; // @[sm_x652_inr_Foreach.scala 81:114:@60845.4]
  assign _T_765 = io_rr & _T_764; // @[sm_x652_inr_Foreach.scala 81:111:@60846.4]
  assign _T_770 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 56:10:@60849.4]
  assign _T_771 = _T_765 & _T_770; // @[sm_x652_inr_Foreach.scala 81:131:@60850.4]
  assign _T_772 = _T_771 & b553; // @[sm_x652_inr_Foreach.scala 81:228:@60851.4]
  assign _T_806 = $signed(io_in_b550_number); // @[Math.scala 510:37:@60885.4]
  assign x790_x647_D3 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@60916.4 package.scala 96:25:@60917.4]
  assign x789_x641_elem_0_D1_number = RetimeWrapper_io_out; // @[package.scala 96:25:@60906.4 package.scala 96:25:@60907.4]
  assign x648_sum_number = x648_sum_1_io_result; // @[Math.scala 154:22:@60896.4 Math.scala 155:14:@60897.4]
  assign _T_850 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@60963.4 package.scala 96:25:@60964.4]
  assign _T_852 = io_rr ? _T_850 : 1'h0; // @[implicits.scala 56:10:@60965.4]
  assign _T_853 = _T_764 & _T_852; // @[sm_x652_inr_Foreach.scala 115:117:@60966.4]
  assign _T_855 = _T_853 & _T_764; // @[sm_x652_inr_Foreach.scala 115:214:@60968.4]
  assign x792_b553_D3 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@60939.4 package.scala 96:25:@60940.4]
  assign _T_857 = _T_855 & x792_b553_D3; // @[sm_x652_inr_Foreach.scala 115:259:@60970.4]
  assign x791_b543_D3 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@60929.4 package.scala 96:25:@60930.4]
  assign _T_869 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@60988.4 package.scala 96:25:@60989.4]
  assign _T_871 = io_rr ? _T_869 : 1'h0; // @[implicits.scala 56:10:@60990.4]
  assign _T_872 = _T_764 & _T_871; // @[sm_x652_inr_Foreach.scala 120:117:@60991.4]
  assign _T_874 = _T_872 & _T_764; // @[sm_x652_inr_Foreach.scala 120:214:@60993.4]
  assign _T_876 = _T_874 & x792_b553_D3; // @[sm_x652_inr_Foreach.scala 120:259:@60995.4]
  assign _T_881 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@61008.4 package.scala 96:25:@61009.4]
  assign b551_number = __io_result; // @[Math.scala 723:22:@60836.4 Math.scala 724:14:@60837.4]
  assign x793_b551_D3_number = RetimeWrapper_4_io_out; // @[package.scala 96:25:@60949.4 package.scala 96:25:@60950.4]
  assign io_in_x558_tmp_4_rPort_0_ofs_0 = b551_number[1:0]; // @[MemInterfaceType.scala 107:54:@60855.4]
  assign io_in_x558_tmp_4_rPort_0_en_0 = _T_772 & io_in_b543; // @[MemInterfaceType.scala 110:79:@60857.4]
  assign io_in_x558_tmp_4_sEn_6 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@61011.4]
  assign io_in_x558_tmp_4_sDone_6 = io_rr ? _T_881 : 1'h0; // @[MemInterfaceType.scala 197:17:@61012.4]
  assign io_in_x545_accum_1_wPort_0_ofs_0 = x793_b551_D3_number[1:0]; // @[MemInterfaceType.scala 89:54:@60973.4]
  assign io_in_x545_accum_1_wPort_0_data_0 = x790_x647_D3 ? x789_x641_elem_0_D1_number : x648_sum_number; // @[MemInterfaceType.scala 90:56:@60974.4]
  assign io_in_x545_accum_1_wPort_0_en_0 = _T_857 & x791_b543_D3; // @[MemInterfaceType.scala 93:57:@60976.4]
  assign io_in_x544_accum_0_rPort_0_ofs_0 = b551_number[1:0]; // @[MemInterfaceType.scala 107:54:@60876.4]
  assign io_in_x544_accum_0_rPort_0_en_0 = _T_772 & io_in_b543; // @[MemInterfaceType.scala 110:79:@60878.4]
  assign io_in_x544_accum_0_wPort_0_ofs_0 = x793_b551_D3_number[1:0]; // @[MemInterfaceType.scala 89:54:@60998.4]
  assign io_in_x544_accum_0_wPort_0_data_0 = x790_x647_D3 ? x789_x641_elem_0_D1_number : x648_sum_number; // @[MemInterfaceType.scala 90:56:@60999.4]
  assign io_in_x544_accum_0_wPort_0_en_0 = _T_876 & x791_b543_D3; // @[MemInterfaceType.scala 93:57:@61001.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@60834.4]
  assign x648_sum_1_clock = clock; // @[:@60891.4]
  assign x648_sum_1_reset = reset; // @[:@60892.4]
  assign x648_sum_1_io_a = io_in_x558_tmp_4_rPort_0_output_0; // @[Math.scala 151:17:@60893.4]
  assign x648_sum_1_io_b = io_in_x544_accum_0_rPort_0_output_0; // @[Math.scala 152:17:@60894.4]
  assign RetimeWrapper_clock = clock; // @[:@60902.4]
  assign RetimeWrapper_reset = reset; // @[:@60903.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@60905.4]
  assign RetimeWrapper_io_in = io_in_x558_tmp_4_rPort_0_output_0; // @[package.scala 94:16:@60904.4]
  assign RetimeWrapper_1_clock = clock; // @[:@60912.4]
  assign RetimeWrapper_1_reset = reset; // @[:@60913.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@60915.4]
  assign RetimeWrapper_1_io_in = $signed(_T_806) == $signed(32'sh0); // @[package.scala 94:16:@60914.4]
  assign RetimeWrapper_2_clock = clock; // @[:@60925.4]
  assign RetimeWrapper_2_reset = reset; // @[:@60926.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@60928.4]
  assign RetimeWrapper_2_io_in = io_in_b543; // @[package.scala 94:16:@60927.4]
  assign RetimeWrapper_3_clock = clock; // @[:@60935.4]
  assign RetimeWrapper_3_reset = reset; // @[:@60936.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@60938.4]
  assign RetimeWrapper_3_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@60937.4]
  assign RetimeWrapper_4_clock = clock; // @[:@60945.4]
  assign RetimeWrapper_4_reset = reset; // @[:@60946.4]
  assign RetimeWrapper_4_io_in = __io_result; // @[package.scala 94:16:@60947.4]
  assign RetimeWrapper_5_clock = clock; // @[:@60959.4]
  assign RetimeWrapper_5_reset = reset; // @[:@60960.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@60962.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@60961.4]
  assign RetimeWrapper_6_clock = clock; // @[:@60984.4]
  assign RetimeWrapper_6_reset = reset; // @[:@60985.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@60987.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@60986.4]
  assign RetimeWrapper_7_clock = clock; // @[:@61004.4]
  assign RetimeWrapper_7_reset = reset; // @[:@61005.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@61007.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_done; // @[package.scala 94:16:@61006.4]
endmodule
module x653_outr_Reduce_kernelx653_outr_Reduce_concrete1( // @[:@61046.2]
  input         clock, // @[:@61047.4]
  input         reset, // @[:@61048.4]
  output [8:0]  io_in_x472_A_sram_1_rPort_0_ofs_0, // @[:@61049.4]
  output        io_in_x472_A_sram_1_rPort_0_en_0, // @[:@61049.4]
  input  [31:0] io_in_x472_A_sram_1_rPort_0_output_0, // @[:@61049.4]
  input  [31:0] io_in_b542_number, // @[:@61049.4]
  output [8:0]  io_in_x471_A_sram_0_rPort_0_ofs_0, // @[:@61049.4]
  output        io_in_x471_A_sram_0_rPort_0_en_0, // @[:@61049.4]
  input  [31:0] io_in_x471_A_sram_0_rPort_0_output_0, // @[:@61049.4]
  output [1:0]  io_in_x545_accum_1_wPort_0_ofs_0, // @[:@61049.4]
  output [31:0] io_in_x545_accum_1_wPort_0_data_0, // @[:@61049.4]
  output        io_in_x545_accum_1_wPort_0_en_0, // @[:@61049.4]
  output        io_in_x545_accum_1_sEn_0, // @[:@61049.4]
  output        io_in_x545_accum_1_sDone_0, // @[:@61049.4]
  output [1:0]  io_in_x544_accum_0_rPort_0_ofs_0, // @[:@61049.4]
  output        io_in_x544_accum_0_rPort_0_en_0, // @[:@61049.4]
  input  [31:0] io_in_x544_accum_0_rPort_0_output_0, // @[:@61049.4]
  output [1:0]  io_in_x544_accum_0_wPort_0_ofs_0, // @[:@61049.4]
  output [31:0] io_in_x544_accum_0_wPort_0_data_0, // @[:@61049.4]
  output        io_in_x544_accum_0_wPort_0_en_0, // @[:@61049.4]
  output        io_in_x549_ctrchain_input_reset, // @[:@61049.4]
  output        io_in_x549_ctrchain_input_enable, // @[:@61049.4]
  input  [3:0]  io_in_x549_ctrchain_output_counts_0, // @[:@61049.4]
  input         io_in_x549_ctrchain_output_oobs_0, // @[:@61049.4]
  input         io_in_x549_ctrchain_output_done, // @[:@61049.4]
  input         io_in_b543, // @[:@61049.4]
  input         io_sigsIn_done, // @[:@61049.4]
  input         io_sigsIn_baseEn, // @[:@61049.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@61049.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@61049.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@61049.4]
  input         io_sigsIn_smEnableOuts_3, // @[:@61049.4]
  input         io_sigsIn_smEnableOuts_4, // @[:@61049.4]
  input         io_sigsIn_smEnableOuts_5, // @[:@61049.4]
  input         io_sigsIn_smEnableOuts_6, // @[:@61049.4]
  input         io_sigsIn_smChildAcks_0, // @[:@61049.4]
  input         io_sigsIn_smChildAcks_1, // @[:@61049.4]
  input         io_sigsIn_smChildAcks_2, // @[:@61049.4]
  input         io_sigsIn_smChildAcks_3, // @[:@61049.4]
  input         io_sigsIn_smChildAcks_4, // @[:@61049.4]
  input         io_sigsIn_smChildAcks_5, // @[:@61049.4]
  input         io_sigsIn_smChildAcks_6, // @[:@61049.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@61049.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@61049.4]
  output        io_sigsOut_smDoneIn_0, // @[:@61049.4]
  output        io_sigsOut_smDoneIn_1, // @[:@61049.4]
  output        io_sigsOut_smDoneIn_2, // @[:@61049.4]
  output        io_sigsOut_smDoneIn_3, // @[:@61049.4]
  output        io_sigsOut_smDoneIn_4, // @[:@61049.4]
  output        io_sigsOut_smDoneIn_5, // @[:@61049.4]
  output        io_sigsOut_smDoneIn_6, // @[:@61049.4]
  output        io_sigsOut_smMaskIn_0, // @[:@61049.4]
  output        io_sigsOut_smMaskIn_1, // @[:@61049.4]
  output        io_sigsOut_smMaskIn_2, // @[:@61049.4]
  output        io_sigsOut_smMaskIn_4, // @[:@61049.4]
  output        io_sigsOut_smMaskIn_5, // @[:@61049.4]
  input         io_rr // @[:@61049.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@61152.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@61152.4]
  wire  b550_chain_clock; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_reset; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire [31:0] b550_chain_io_rPort_5_output_0; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire [31:0] b550_chain_io_rPort_4_output_0; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire [31:0] b550_chain_io_rPort_3_output_0; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire [31:0] b550_chain_io_rPort_2_output_0; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire [31:0] b550_chain_io_rPort_1_output_0; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire [31:0] b550_chain_io_rPort_0_output_0; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire [31:0] b550_chain_io_wPort_0_data_0; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_io_wPort_0_reset; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_io_wPort_0_en_0; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_io_sEn_0; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_io_sEn_1; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_io_sEn_2; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_io_sEn_3; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_io_sEn_4; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_io_sEn_5; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_io_sEn_6; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_io_sDone_0; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_io_sDone_1; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_io_sDone_2; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_io_sDone_3; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_io_sDone_4; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_io_sDone_5; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  b550_chain_io_sDone_6; // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@61224.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@61224.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@61224.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@61224.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@61224.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@61236.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@61236.4]
  wire [31:0] __2_io_b; // @[Math.scala 720:24:@61247.4]
  wire [31:0] __2_io_result; // @[Math.scala 720:24:@61247.4]
  wire [31:0] __3_io_b; // @[Math.scala 720:24:@61258.4]
  wire [31:0] __3_io_result; // @[Math.scala 720:24:@61258.4]
  wire [31:0] __4_io_b; // @[Math.scala 720:24:@61269.4]
  wire [31:0] __4_io_result; // @[Math.scala 720:24:@61269.4]
  wire [31:0] __5_io_b; // @[Math.scala 720:24:@61280.4]
  wire [31:0] __5_io_result; // @[Math.scala 720:24:@61280.4]
  wire [31:0] __6_io_b; // @[Math.scala 720:24:@61291.4]
  wire [31:0] __6_io_result; // @[Math.scala 720:24:@61291.4]
  wire  b552_chain_clock; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_reset; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_rPort_4_output_0; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_rPort_3_output_0; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_rPort_1_output_0; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_rPort_0_output_0; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_wPort_0_data_0; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_wPort_0_reset; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_wPort_0_en_0; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_sEn_0; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_sEn_1; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_sEn_2; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_sEn_3; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_sEn_4; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_sEn_5; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_sEn_6; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_sDone_0; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_sDone_1; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_sDone_2; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_sDone_3; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_sDone_4; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_sDone_5; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  b552_chain_io_sDone_6; // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@61364.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@61364.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@61364.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@61364.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@61364.4]
  wire  x554_tmp_0_clock; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x554_tmp_0_reset; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire [1:0] x554_tmp_0_io_rPort_0_ofs_0; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x554_tmp_0_io_rPort_0_en_0; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire [31:0] x554_tmp_0_io_rPort_0_output_0; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire [1:0] x554_tmp_0_io_wPort_1_ofs_0; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire [31:0] x554_tmp_0_io_wPort_1_data_0; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x554_tmp_0_io_wPort_1_en_0; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire [1:0] x554_tmp_0_io_wPort_0_ofs_0; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire [31:0] x554_tmp_0_io_wPort_0_data_0; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x554_tmp_0_io_wPort_0_en_0; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x554_tmp_0_io_sEn_0; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x554_tmp_0_io_sEn_1; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x554_tmp_0_io_sEn_2; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x554_tmp_0_io_sEn_3; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x554_tmp_0_io_sEn_4; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x554_tmp_0_io_sEn_5; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x554_tmp_0_io_sDone_0; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x554_tmp_0_io_sDone_1; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x554_tmp_0_io_sDone_2; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x554_tmp_0_io_sDone_3; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x554_tmp_0_io_sDone_4; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x554_tmp_0_io_sDone_5; // @[m_x554_tmp_0.scala 28:22:@61379.4]
  wire  x555_tmp_1_clock; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x555_tmp_1_reset; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire [1:0] x555_tmp_1_io_rPort_0_ofs_0; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x555_tmp_1_io_rPort_0_en_0; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire [31:0] x555_tmp_1_io_rPort_0_output_0; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire [1:0] x555_tmp_1_io_wPort_1_ofs_0; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire [31:0] x555_tmp_1_io_wPort_1_data_0; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x555_tmp_1_io_wPort_1_en_0; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire [1:0] x555_tmp_1_io_wPort_0_ofs_0; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire [31:0] x555_tmp_1_io_wPort_0_data_0; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x555_tmp_1_io_wPort_0_en_0; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x555_tmp_1_io_sEn_0; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x555_tmp_1_io_sEn_1; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x555_tmp_1_io_sEn_2; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x555_tmp_1_io_sEn_3; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x555_tmp_1_io_sEn_4; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x555_tmp_1_io_sEn_5; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x555_tmp_1_io_sDone_0; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x555_tmp_1_io_sDone_1; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x555_tmp_1_io_sDone_2; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x555_tmp_1_io_sDone_3; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x555_tmp_1_io_sDone_4; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x555_tmp_1_io_sDone_5; // @[m_x555_tmp_1.scala 28:22:@61426.4]
  wire  x556_tmp_2_clock; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x556_tmp_2_reset; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire [1:0] x556_tmp_2_io_rPort_0_ofs_0; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x556_tmp_2_io_rPort_0_en_0; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire [31:0] x556_tmp_2_io_rPort_0_output_0; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire [1:0] x556_tmp_2_io_wPort_1_ofs_0; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire [31:0] x556_tmp_2_io_wPort_1_data_0; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x556_tmp_2_io_wPort_1_en_0; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire [1:0] x556_tmp_2_io_wPort_0_ofs_0; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire [31:0] x556_tmp_2_io_wPort_0_data_0; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x556_tmp_2_io_wPort_0_en_0; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x556_tmp_2_io_sEn_0; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x556_tmp_2_io_sEn_1; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x556_tmp_2_io_sEn_2; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x556_tmp_2_io_sEn_3; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x556_tmp_2_io_sEn_4; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x556_tmp_2_io_sEn_5; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x556_tmp_2_io_sDone_0; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x556_tmp_2_io_sDone_1; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x556_tmp_2_io_sDone_2; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x556_tmp_2_io_sDone_3; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x556_tmp_2_io_sDone_4; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x556_tmp_2_io_sDone_5; // @[m_x556_tmp_2.scala 28:22:@61473.4]
  wire  x557_tmp_3_clock; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x557_tmp_3_reset; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire [1:0] x557_tmp_3_io_rPort_0_ofs_0; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x557_tmp_3_io_rPort_0_en_0; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire [31:0] x557_tmp_3_io_rPort_0_output_0; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire [1:0] x557_tmp_3_io_wPort_1_ofs_0; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire [31:0] x557_tmp_3_io_wPort_1_data_0; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x557_tmp_3_io_wPort_1_en_0; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire [1:0] x557_tmp_3_io_wPort_0_ofs_0; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire [31:0] x557_tmp_3_io_wPort_0_data_0; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x557_tmp_3_io_wPort_0_en_0; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x557_tmp_3_io_sEn_0; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x557_tmp_3_io_sEn_1; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x557_tmp_3_io_sEn_2; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x557_tmp_3_io_sEn_3; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x557_tmp_3_io_sEn_4; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x557_tmp_3_io_sEn_5; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x557_tmp_3_io_sDone_0; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x557_tmp_3_io_sDone_1; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x557_tmp_3_io_sDone_2; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x557_tmp_3_io_sDone_3; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x557_tmp_3_io_sDone_4; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x557_tmp_3_io_sDone_5; // @[m_x557_tmp_3.scala 28:22:@61520.4]
  wire  x558_tmp_4_clock; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_reset; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire [1:0] x558_tmp_4_io_rPort_0_ofs_0; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_rPort_0_en_0; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire [31:0] x558_tmp_4_io_rPort_0_output_0; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire [1:0] x558_tmp_4_io_wPort_1_ofs_0; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire [31:0] x558_tmp_4_io_wPort_1_data_0; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_wPort_1_en_0; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire [1:0] x558_tmp_4_io_wPort_0_ofs_0; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire [31:0] x558_tmp_4_io_wPort_0_data_0; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_wPort_0_en_0; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_sEn_0; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_sEn_1; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_sEn_2; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_sEn_3; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_sEn_4; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_sEn_5; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_sEn_6; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_sDone_0; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_sDone_1; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_sDone_2; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_sDone_3; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_sDone_4; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_sDone_5; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x558_tmp_4_io_sDone_6; // @[m_x558_tmp_4.scala 28:22:@61567.4]
  wire  x560_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@61616.4]
  wire  x560_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@61616.4]
  wire  x560_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@61616.4]
  wire  x560_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@61616.4]
  wire [3:0] x560_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@61616.4]
  wire  x560_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@61616.4]
  wire  x560_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@61616.4]
  wire  x579_inr_Foreach_sm_clock; // @[sm_x579_inr_Foreach.scala 35:18:@61669.4]
  wire  x579_inr_Foreach_sm_reset; // @[sm_x579_inr_Foreach.scala 35:18:@61669.4]
  wire  x579_inr_Foreach_sm_io_enable; // @[sm_x579_inr_Foreach.scala 35:18:@61669.4]
  wire  x579_inr_Foreach_sm_io_done; // @[sm_x579_inr_Foreach.scala 35:18:@61669.4]
  wire  x579_inr_Foreach_sm_io_ctrDone; // @[sm_x579_inr_Foreach.scala 35:18:@61669.4]
  wire  x579_inr_Foreach_sm_io_datapathEn; // @[sm_x579_inr_Foreach.scala 35:18:@61669.4]
  wire  x579_inr_Foreach_sm_io_ctrInc; // @[sm_x579_inr_Foreach.scala 35:18:@61669.4]
  wire  x579_inr_Foreach_sm_io_ctrRst; // @[sm_x579_inr_Foreach.scala 35:18:@61669.4]
  wire  x579_inr_Foreach_sm_io_parentAck; // @[sm_x579_inr_Foreach.scala 35:18:@61669.4]
  wire  x579_inr_Foreach_sm_io_backpressure; // @[sm_x579_inr_Foreach.scala 35:18:@61669.4]
  wire  x579_inr_Foreach_sm_io_break; // @[sm_x579_inr_Foreach.scala 35:18:@61669.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@61698.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@61698.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@61698.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@61698.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@61698.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@61707.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@61707.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@61707.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@61707.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@61707.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@61717.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@61717.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@61717.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@61717.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@61717.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@61759.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@61759.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@61759.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@61759.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@61759.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@61767.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@61767.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@61767.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@61767.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@61767.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_clock; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_reset; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [1:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_ofs_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_data_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_en_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_sEn_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_sDone_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b550_number; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [8:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_en_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_output_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b542_number; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [8:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_en_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_output_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [1:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_ofs_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_data_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_en_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_sEn_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_sDone_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [1:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_ofs_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_data_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_en_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b552; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [1:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_ofs_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_data_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_en_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_sEn_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_sDone_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [1:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_ofs_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_data_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_en_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_sEn_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_sDone_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b543; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_done; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire [31:0] x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_rr; // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
  wire  x580_r_0_clock; // @[m_x580_r_0.scala 28:22:@62245.4]
  wire  x580_r_0_reset; // @[m_x580_r_0.scala 28:22:@62245.4]
  wire  x580_r_0_io_rPort_1_en_0; // @[m_x580_r_0.scala 28:22:@62245.4]
  wire [31:0] x580_r_0_io_rPort_1_output_0; // @[m_x580_r_0.scala 28:22:@62245.4]
  wire  x580_r_0_io_rPort_0_en_0; // @[m_x580_r_0.scala 28:22:@62245.4]
  wire [31:0] x580_r_0_io_rPort_0_output_0; // @[m_x580_r_0.scala 28:22:@62245.4]
  wire [31:0] x580_r_0_io_wPort_0_data_0; // @[m_x580_r_0.scala 28:22:@62245.4]
  wire  x580_r_0_io_wPort_0_en_0; // @[m_x580_r_0.scala 28:22:@62245.4]
  wire  x580_r_0_io_sEn_0; // @[m_x580_r_0.scala 28:22:@62245.4]
  wire  x580_r_0_io_sEn_1; // @[m_x580_r_0.scala 28:22:@62245.4]
  wire  x580_r_0_io_sEn_2; // @[m_x580_r_0.scala 28:22:@62245.4]
  wire  x580_r_0_io_sDone_0; // @[m_x580_r_0.scala 28:22:@62245.4]
  wire  x580_r_0_io_sDone_1; // @[m_x580_r_0.scala 28:22:@62245.4]
  wire  x580_r_0_io_sDone_2; // @[m_x580_r_0.scala 28:22:@62245.4]
  wire  x593_inr_UnitPipe_sm_clock; // @[sm_x593_inr_UnitPipe.scala 33:18:@62320.4]
  wire  x593_inr_UnitPipe_sm_reset; // @[sm_x593_inr_UnitPipe.scala 33:18:@62320.4]
  wire  x593_inr_UnitPipe_sm_io_enable; // @[sm_x593_inr_UnitPipe.scala 33:18:@62320.4]
  wire  x593_inr_UnitPipe_sm_io_done; // @[sm_x593_inr_UnitPipe.scala 33:18:@62320.4]
  wire  x593_inr_UnitPipe_sm_io_ctrDone; // @[sm_x593_inr_UnitPipe.scala 33:18:@62320.4]
  wire  x593_inr_UnitPipe_sm_io_datapathEn; // @[sm_x593_inr_UnitPipe.scala 33:18:@62320.4]
  wire  x593_inr_UnitPipe_sm_io_ctrInc; // @[sm_x593_inr_UnitPipe.scala 33:18:@62320.4]
  wire  x593_inr_UnitPipe_sm_io_parentAck; // @[sm_x593_inr_UnitPipe.scala 33:18:@62320.4]
  wire  x593_inr_UnitPipe_sm_io_backpressure; // @[sm_x593_inr_UnitPipe.scala 33:18:@62320.4]
  wire  x593_inr_UnitPipe_sm_io_break; // @[sm_x593_inr_UnitPipe.scala 33:18:@62320.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@62353.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@62353.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@62353.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@62353.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@62353.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@62363.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@62363.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@62363.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@62363.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@62363.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@62399.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@62399.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@62399.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@62399.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@62399.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@62407.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@62407.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@62407.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@62407.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@62407.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_clock; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_reset; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_rPort_0_en_0; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire [31:0] x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_rPort_0_output_0; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_1; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_1; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_rPort_0_en_0; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire [31:0] x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_rPort_0_output_0; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_1; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_1; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_1; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_1; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_1; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_1; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire [31:0] x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_wPort_0_data_0; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_wPort_0_en_0; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_sEn_0; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_sDone_0; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_rPort_0_en_0; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire [31:0] x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_rPort_0_output_0; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_1; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_1; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_done; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_baseEn; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_break; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_rr; // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
  wire  x594_force_0_clock; // @[m_x594_force_0.scala 27:22:@62880.4]
  wire  x594_force_0_reset; // @[m_x594_force_0.scala 27:22:@62880.4]
  wire  x594_force_0_io_rPort_0_en_0; // @[m_x594_force_0.scala 27:22:@62880.4]
  wire [31:0] x594_force_0_io_rPort_0_output_0; // @[m_x594_force_0.scala 27:22:@62880.4]
  wire [31:0] x594_force_0_io_wPort_0_data_0; // @[m_x594_force_0.scala 27:22:@62880.4]
  wire  x594_force_0_io_wPort_0_en_0; // @[m_x594_force_0.scala 27:22:@62880.4]
  wire  x594_force_0_io_sEn_0; // @[m_x594_force_0.scala 27:22:@62880.4]
  wire  x594_force_0_io_sEn_1; // @[m_x594_force_0.scala 27:22:@62880.4]
  wire  x594_force_0_io_sDone_0; // @[m_x594_force_0.scala 27:22:@62880.4]
  wire  x594_force_0_io_sDone_1; // @[m_x594_force_0.scala 27:22:@62880.4]
  wire  x595_reg_clock; // @[m_x595_reg.scala 28:22:@62910.4]
  wire  x595_reg_reset; // @[m_x595_reg.scala 28:22:@62910.4]
  wire  x595_reg_io_rPort_1_output_0; // @[m_x595_reg.scala 28:22:@62910.4]
  wire  x595_reg_io_rPort_0_output_0; // @[m_x595_reg.scala 28:22:@62910.4]
  wire  x595_reg_io_wPort_0_data_0; // @[m_x595_reg.scala 28:22:@62910.4]
  wire  x595_reg_io_wPort_0_reset; // @[m_x595_reg.scala 28:22:@62910.4]
  wire  x595_reg_io_wPort_0_en_0; // @[m_x595_reg.scala 28:22:@62910.4]
  wire  x595_reg_io_sEn_0; // @[m_x595_reg.scala 28:22:@62910.4]
  wire  x595_reg_io_sEn_1; // @[m_x595_reg.scala 28:22:@62910.4]
  wire  x595_reg_io_sDone_0; // @[m_x595_reg.scala 28:22:@62910.4]
  wire  x595_reg_io_sDone_1; // @[m_x595_reg.scala 28:22:@62910.4]
  wire  x596_reg_clock; // @[m_x596_reg.scala 27:22:@62947.4]
  wire  x596_reg_reset; // @[m_x596_reg.scala 27:22:@62947.4]
  wire  x596_reg_io_rPort_0_output_0; // @[m_x596_reg.scala 27:22:@62947.4]
  wire  x596_reg_io_wPort_0_data_0; // @[m_x596_reg.scala 27:22:@62947.4]
  wire  x596_reg_io_wPort_0_reset; // @[m_x596_reg.scala 27:22:@62947.4]
  wire  x596_reg_io_wPort_0_en_0; // @[m_x596_reg.scala 27:22:@62947.4]
  wire  x596_reg_io_sEn_0; // @[m_x596_reg.scala 27:22:@62947.4]
  wire  x596_reg_io_sEn_1; // @[m_x596_reg.scala 27:22:@62947.4]
  wire  x596_reg_io_sDone_0; // @[m_x596_reg.scala 27:22:@62947.4]
  wire  x596_reg_io_sDone_1; // @[m_x596_reg.scala 27:22:@62947.4]
  wire  x605_inr_UnitPipe_sm_clock; // @[sm_x605_inr_UnitPipe.scala 33:18:@63013.4]
  wire  x605_inr_UnitPipe_sm_reset; // @[sm_x605_inr_UnitPipe.scala 33:18:@63013.4]
  wire  x605_inr_UnitPipe_sm_io_enable; // @[sm_x605_inr_UnitPipe.scala 33:18:@63013.4]
  wire  x605_inr_UnitPipe_sm_io_done; // @[sm_x605_inr_UnitPipe.scala 33:18:@63013.4]
  wire  x605_inr_UnitPipe_sm_io_doneLatch; // @[sm_x605_inr_UnitPipe.scala 33:18:@63013.4]
  wire  x605_inr_UnitPipe_sm_io_ctrDone; // @[sm_x605_inr_UnitPipe.scala 33:18:@63013.4]
  wire  x605_inr_UnitPipe_sm_io_datapathEn; // @[sm_x605_inr_UnitPipe.scala 33:18:@63013.4]
  wire  x605_inr_UnitPipe_sm_io_ctrInc; // @[sm_x605_inr_UnitPipe.scala 33:18:@63013.4]
  wire  x605_inr_UnitPipe_sm_io_ctrRst; // @[sm_x605_inr_UnitPipe.scala 33:18:@63013.4]
  wire  x605_inr_UnitPipe_sm_io_parentAck; // @[sm_x605_inr_UnitPipe.scala 33:18:@63013.4]
  wire  x605_inr_UnitPipe_sm_io_backpressure; // @[sm_x605_inr_UnitPipe.scala 33:18:@63013.4]
  wire  x605_inr_UnitPipe_sm_io_break; // @[sm_x605_inr_UnitPipe.scala 33:18:@63013.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@63046.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@63046.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@63046.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@63046.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@63046.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@63056.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@63056.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@63056.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@63056.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@63056.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@63092.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@63092.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@63092.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@63092.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@63092.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@63100.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@63100.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@63100.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@63100.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@63100.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_clock; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_reset; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_2; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_2; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_2; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_2; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_2; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_2; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_2; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_2; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_rPort_0_en_0; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire [31:0] x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_rPort_0_output_0; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_sEn_1; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_sDone_1; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_data_0; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_reset; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_en_0; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_reset; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_sEn_0; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_sDone_0; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_2; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_2; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_data_0; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_reset; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_en_0; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_reset; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_sEn_0; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_sDone_0; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_done; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_baseEn; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_break; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_rr; // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
  wire  x621_inr_Switch_sm_clock; // @[sm_x621_inr_Switch.scala 33:18:@63732.4]
  wire  x621_inr_Switch_sm_reset; // @[sm_x621_inr_Switch.scala 33:18:@63732.4]
  wire  x621_inr_Switch_sm_io_enable; // @[sm_x621_inr_Switch.scala 33:18:@63732.4]
  wire  x621_inr_Switch_sm_io_done; // @[sm_x621_inr_Switch.scala 33:18:@63732.4]
  wire  x621_inr_Switch_sm_io_parentAck; // @[sm_x621_inr_Switch.scala 33:18:@63732.4]
  wire  x621_inr_Switch_sm_io_backpressure; // @[sm_x621_inr_Switch.scala 33:18:@63732.4]
  wire  x621_inr_Switch_sm_io_doneIn_0; // @[sm_x621_inr_Switch.scala 33:18:@63732.4]
  wire  x621_inr_Switch_sm_io_doneIn_1; // @[sm_x621_inr_Switch.scala 33:18:@63732.4]
  wire  x621_inr_Switch_sm_io_childAck_0; // @[sm_x621_inr_Switch.scala 33:18:@63732.4]
  wire  x621_inr_Switch_sm_io_childAck_1; // @[sm_x621_inr_Switch.scala 33:18:@63732.4]
  wire  x621_inr_Switch_sm_io_selectsIn_0; // @[sm_x621_inr_Switch.scala 33:18:@63732.4]
  wire  x621_inr_Switch_sm_io_selectsIn_1; // @[sm_x621_inr_Switch.scala 33:18:@63732.4]
  wire  x621_inr_Switch_sm_io_selectsOut_0; // @[sm_x621_inr_Switch.scala 33:18:@63732.4]
  wire  x621_inr_Switch_sm_io_selectsOut_1; // @[sm_x621_inr_Switch.scala 33:18:@63732.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@63769.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@63769.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@63769.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@63769.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@63769.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@63779.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@63779.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@63779.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@63779.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@63779.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@63821.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@63821.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@63821.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@63821.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@63821.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@63829.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@63829.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@63829.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@63829.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@63829.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_clock; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_reset; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x555_tmp_1_sEn_3; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x555_tmp_1_sDone_3; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x554_tmp_0_sEn_3; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x554_tmp_0_sDone_3; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x558_tmp_4_sEn_3; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x558_tmp_4_sDone_3; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x736_rd_x596; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x557_tmp_3_sEn_3; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x557_tmp_3_sDone_3; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_rPort_1_en_0; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire [31:0] x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_rPort_1_output_0; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_sEn_2; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_sDone_2; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_rPort_1_output_0; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_sEn_1; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_sDone_1; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x556_tmp_2_sEn_3; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x556_tmp_2_sDone_3; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x735_rd_x595; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x596_reg_sEn_1; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x596_reg_sDone_1; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_done; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_baseEn; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smSelectsOut_0; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smSelectsOut_1; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_rr; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire [31:0] x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_ret_number; // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
  wire  x623_inr_UnitPipe_sm_clock; // @[sm_x623_inr_UnitPipe.scala 34:18:@64431.4]
  wire  x623_inr_UnitPipe_sm_reset; // @[sm_x623_inr_UnitPipe.scala 34:18:@64431.4]
  wire  x623_inr_UnitPipe_sm_io_enable; // @[sm_x623_inr_UnitPipe.scala 34:18:@64431.4]
  wire  x623_inr_UnitPipe_sm_io_done; // @[sm_x623_inr_UnitPipe.scala 34:18:@64431.4]
  wire  x623_inr_UnitPipe_sm_io_doneLatch; // @[sm_x623_inr_UnitPipe.scala 34:18:@64431.4]
  wire  x623_inr_UnitPipe_sm_io_ctrDone; // @[sm_x623_inr_UnitPipe.scala 34:18:@64431.4]
  wire  x623_inr_UnitPipe_sm_io_datapathEn; // @[sm_x623_inr_UnitPipe.scala 34:18:@64431.4]
  wire  x623_inr_UnitPipe_sm_io_ctrInc; // @[sm_x623_inr_UnitPipe.scala 34:18:@64431.4]
  wire  x623_inr_UnitPipe_sm_io_parentAck; // @[sm_x623_inr_UnitPipe.scala 34:18:@64431.4]
  wire  x623_inr_UnitPipe_sm_io_backpressure; // @[sm_x623_inr_UnitPipe.scala 34:18:@64431.4]
  wire  x623_inr_UnitPipe_sm_io_break; // @[sm_x623_inr_UnitPipe.scala 34:18:@64431.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@64464.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@64464.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@64464.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@64464.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@64464.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@64474.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@64474.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@64474.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@64474.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@64474.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@64510.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@64510.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@64510.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@64510.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@64510.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@64518.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@64518.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@64518.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@64518.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@64518.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_clock; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_reset; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_4; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_4; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_4; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_4; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_4; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_4; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire [31:0] x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_wPort_0_data_0; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_wPort_0_en_0; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_sEn_0; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_sDone_0; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire [31:0] x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x621_inr_Switch_number; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_4; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_4; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_4; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_4; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_done; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_baseEn; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_break; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_rr; // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
  wire  x625_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@64967.4]
  wire  x625_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@64967.4]
  wire  x625_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@64967.4]
  wire  x625_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@64967.4]
  wire [3:0] x625_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@64967.4]
  wire  x625_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@64967.4]
  wire  x625_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@64967.4]
  wire  x639_inr_Foreach_sm_clock; // @[sm_x639_inr_Foreach.scala 33:18:@65020.4]
  wire  x639_inr_Foreach_sm_reset; // @[sm_x639_inr_Foreach.scala 33:18:@65020.4]
  wire  x639_inr_Foreach_sm_io_enable; // @[sm_x639_inr_Foreach.scala 33:18:@65020.4]
  wire  x639_inr_Foreach_sm_io_done; // @[sm_x639_inr_Foreach.scala 33:18:@65020.4]
  wire  x639_inr_Foreach_sm_io_rst; // @[sm_x639_inr_Foreach.scala 33:18:@65020.4]
  wire  x639_inr_Foreach_sm_io_ctrDone; // @[sm_x639_inr_Foreach.scala 33:18:@65020.4]
  wire  x639_inr_Foreach_sm_io_datapathEn; // @[sm_x639_inr_Foreach.scala 33:18:@65020.4]
  wire  x639_inr_Foreach_sm_io_ctrInc; // @[sm_x639_inr_Foreach.scala 33:18:@65020.4]
  wire  x639_inr_Foreach_sm_io_ctrRst; // @[sm_x639_inr_Foreach.scala 33:18:@65020.4]
  wire  x639_inr_Foreach_sm_io_parentAck; // @[sm_x639_inr_Foreach.scala 33:18:@65020.4]
  wire  x639_inr_Foreach_sm_io_backpressure; // @[sm_x639_inr_Foreach.scala 33:18:@65020.4]
  wire  x639_inr_Foreach_sm_io_break; // @[sm_x639_inr_Foreach.scala 33:18:@65020.4]
  wire  x639_inr_Foreach_iiCtr_clock; // @[sm_x639_inr_Foreach.scala 34:21:@65045.4]
  wire  x639_inr_Foreach_iiCtr_reset; // @[sm_x639_inr_Foreach.scala 34:21:@65045.4]
  wire  x639_inr_Foreach_iiCtr_io_input_enable; // @[sm_x639_inr_Foreach.scala 34:21:@65045.4]
  wire  x639_inr_Foreach_iiCtr_io_input_reset; // @[sm_x639_inr_Foreach.scala 34:21:@65045.4]
  wire  x639_inr_Foreach_iiCtr_io_output_issue; // @[sm_x639_inr_Foreach.scala 34:21:@65045.4]
  wire  x639_inr_Foreach_iiCtr_io_output_done; // @[sm_x639_inr_Foreach.scala 34:21:@65045.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@65049.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@65049.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@65049.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@65049.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@65049.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@65058.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@65058.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@65058.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@65058.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@65058.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@65068.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@65068.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@65068.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@65068.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@65068.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@65110.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@65110.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@65110.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@65110.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@65110.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@65118.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@65118.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@65118.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@65118.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@65118.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_clock; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_reset; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire [1:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_ofs_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire [31:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_data_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_en_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_sEn_5; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_sDone_5; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire [1:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_ofs_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire [31:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_data_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_en_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_sEn_5; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_sDone_5; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire [1:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_ofs_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire [31:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_data_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_en_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_5; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_5; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_b552; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_rPort_0_en_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire [31:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_rPort_0_output_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_sEn_1; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_sDone_1; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire [1:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_ofs_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_en_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire [31:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_output_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire [1:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_ofs_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire [31:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_data_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_en_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_sEn_5; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_sDone_5; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire [1:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_ofs_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire [31:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_data_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_en_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_sEn_5; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_sDone_5; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_b543; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_done; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_iiIssue; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire [31:0] x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_rr; // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
  wire  x652_inr_Foreach_sm_clock; // @[sm_x652_inr_Foreach.scala 35:18:@65644.4]
  wire  x652_inr_Foreach_sm_reset; // @[sm_x652_inr_Foreach.scala 35:18:@65644.4]
  wire  x652_inr_Foreach_sm_io_enable; // @[sm_x652_inr_Foreach.scala 35:18:@65644.4]
  wire  x652_inr_Foreach_sm_io_done; // @[sm_x652_inr_Foreach.scala 35:18:@65644.4]
  wire  x652_inr_Foreach_sm_io_doneLatch; // @[sm_x652_inr_Foreach.scala 35:18:@65644.4]
  wire  x652_inr_Foreach_sm_io_ctrDone; // @[sm_x652_inr_Foreach.scala 35:18:@65644.4]
  wire  x652_inr_Foreach_sm_io_datapathEn; // @[sm_x652_inr_Foreach.scala 35:18:@65644.4]
  wire  x652_inr_Foreach_sm_io_ctrInc; // @[sm_x652_inr_Foreach.scala 35:18:@65644.4]
  wire  x652_inr_Foreach_sm_io_ctrRst; // @[sm_x652_inr_Foreach.scala 35:18:@65644.4]
  wire  x652_inr_Foreach_sm_io_parentAck; // @[sm_x652_inr_Foreach.scala 35:18:@65644.4]
  wire  x652_inr_Foreach_sm_io_backpressure; // @[sm_x652_inr_Foreach.scala 35:18:@65644.4]
  wire  x652_inr_Foreach_sm_io_break; // @[sm_x652_inr_Foreach.scala 35:18:@65644.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@65673.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@65673.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@65673.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@65673.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@65673.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@65682.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@65682.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@65682.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@65682.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@65682.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@65692.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@65692.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@65692.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@65692.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@65692.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@65733.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@65733.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@65733.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@65733.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@65733.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@65741.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@65741.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@65741.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@65741.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@65741.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_clock; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_reset; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire [31:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_b550_number; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire [1:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_ofs_0; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_en_0; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire [31:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_output_0; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_6; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_6; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire [1:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_ofs_0; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire [31:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_data_0; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_en_0; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire [1:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_ofs_0; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_en_0; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire [31:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_output_0; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire [1:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_ofs_0; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire [31:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_data_0; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_en_0; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_b543; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_done; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire [31:0] x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_rr; // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@65978.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@65978.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@65978.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@65978.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@65978.4]
  wire  b552; // @[sm_x653_outr_Reduce.scala 93:18:@61299.4]
  wire  b552_chain_read_1; // @[sm_x653_outr_Reduce.scala 96:61:@61373.4]
  wire  b552_chain_read_2; // @[sm_x653_outr_Reduce.scala 97:61:@61374.4]
  wire  b552_chain_read_4; // @[sm_x653_outr_Reduce.scala 99:61:@61376.4]
  wire  b552_chain_read_5; // @[sm_x653_outr_Reduce.scala 100:61:@61377.4]
  wire  _T_897; // @[package.scala 96:25:@61703.4 package.scala 96:25:@61704.4]
  wire  _T_901; // @[package.scala 96:25:@61712.4 package.scala 96:25:@61713.4]
  wire  _T_905; // @[package.scala 96:25:@61722.4 package.scala 96:25:@61723.4]
  wire  x579_inr_Foreach_mySignalsIn_mask; // @[sm_x653_outr_Reduce.scala 119:81:@61736.4]
  wire  _T_922; // @[package.scala 96:25:@61764.4 package.scala 96:25:@61765.4]
  wire  _T_928; // @[package.scala 96:25:@61772.4 package.scala 96:25:@61773.4]
  wire  _T_931; // @[SpatialBlocks.scala 137:99:@61775.4]
  wire  _T_933; // @[SpatialBlocks.scala 156:36:@61784.4]
  wire  _T_934; // @[SpatialBlocks.scala 156:78:@61785.4]
  wire  _T_1002; // @[package.scala 100:49:@62348.4]
  reg  _T_1005; // @[package.scala 48:56:@62349.4]
  reg [31:0] _RAND_0;
  wire  _T_1008; // @[package.scala 96:25:@62358.4 package.scala 96:25:@62359.4]
  wire  _T_1012; // @[package.scala 96:25:@62368.4 package.scala 96:25:@62369.4]
  wire  x593_inr_UnitPipe_mySignalsIn_mask; // @[sm_x653_outr_Reduce.scala 131:60:@62381.4]
  wire  _T_1029; // @[package.scala 96:25:@62404.4 package.scala 96:25:@62405.4]
  wire  _T_1035; // @[package.scala 96:25:@62412.4 package.scala 96:25:@62413.4]
  wire  _T_1038; // @[SpatialBlocks.scala 137:99:@62415.4]
  wire  _T_1109; // @[package.scala 100:49:@63041.4]
  reg  _T_1112; // @[package.scala 48:56:@63042.4]
  reg [31:0] _RAND_1;
  wire  _T_1115; // @[package.scala 96:25:@63051.4 package.scala 96:25:@63052.4]
  wire  _T_1119; // @[package.scala 96:25:@63061.4 package.scala 96:25:@63062.4]
  wire  x605_inr_UnitPipe_mySignalsIn_mask; // @[sm_x653_outr_Reduce.scala 145:60:@63074.4]
  wire  _T_1136; // @[package.scala 96:25:@63097.4 package.scala 96:25:@63098.4]
  wire  _T_1142; // @[package.scala 96:25:@63105.4 package.scala 96:25:@63106.4]
  wire  _T_1145; // @[SpatialBlocks.scala 137:99:@63108.4]
  wire  _T_1243; // @[package.scala 96:25:@63774.4 package.scala 96:25:@63775.4]
  wire  _T_1247; // @[package.scala 96:25:@63784.4 package.scala 96:25:@63785.4]
  wire  _T_1265; // @[package.scala 96:25:@63826.4 package.scala 96:25:@63827.4]
  wire  _T_1271; // @[package.scala 96:25:@63834.4 package.scala 96:25:@63835.4]
  wire  _T_1274; // @[SpatialBlocks.scala 137:99:@63837.4]
  wire  _T_1342; // @[package.scala 100:49:@64459.4]
  reg  _T_1345; // @[package.scala 48:56:@64460.4]
  reg [31:0] _RAND_2;
  wire  _T_1348; // @[package.scala 96:25:@64469.4 package.scala 96:25:@64470.4]
  wire  _T_1352; // @[package.scala 96:25:@64479.4 package.scala 96:25:@64480.4]
  wire  x623_inr_UnitPipe_mySignalsIn_mask; // @[sm_x653_outr_Reduce.scala 181:60:@64492.4]
  wire  _T_1369; // @[package.scala 96:25:@64515.4 package.scala 96:25:@64516.4]
  wire  _T_1375; // @[package.scala 96:25:@64523.4 package.scala 96:25:@64524.4]
  wire  _T_1378; // @[SpatialBlocks.scala 137:99:@64526.4]
  wire  _T_1450; // @[package.scala 96:25:@65054.4 package.scala 96:25:@65055.4]
  wire  _T_1454; // @[package.scala 96:25:@65063.4 package.scala 96:25:@65064.4]
  wire  _T_1458; // @[package.scala 96:25:@65073.4 package.scala 96:25:@65074.4]
  wire  x639_inr_Foreach_mySignalsIn_mask; // @[sm_x653_outr_Reduce.scala 196:94:@65087.4]
  wire  _T_1475; // @[package.scala 96:25:@65115.4 package.scala 96:25:@65116.4]
  wire  _T_1481; // @[package.scala 96:25:@65123.4 package.scala 96:25:@65124.4]
  wire  _T_1484; // @[SpatialBlocks.scala 137:99:@65126.4]
  wire  _T_1486; // @[SpatialBlocks.scala 156:36:@65135.4]
  wire  _T_1487; // @[SpatialBlocks.scala 156:78:@65136.4]
  wire  _T_1490; // @[SpatialBlocks.scala 157:128:@65142.4]
  wire  x639_inr_Foreach_mySignalsIn_iiDone; // @[SpatialBlocks.scala 157:126:@65143.4]
  wire  _T_1556; // @[package.scala 96:25:@65678.4 package.scala 96:25:@65679.4]
  wire  _T_1560; // @[package.scala 96:25:@65687.4 package.scala 96:25:@65688.4]
  wire  _T_1564; // @[package.scala 96:25:@65697.4 package.scala 96:25:@65698.4]
  wire  _T_1581; // @[package.scala 96:25:@65738.4 package.scala 96:25:@65739.4]
  wire  _T_1587; // @[package.scala 96:25:@65746.4 package.scala 96:25:@65747.4]
  wire  _T_1590; // @[SpatialBlocks.scala 137:99:@65749.4]
  wire  _T_1592; // @[SpatialBlocks.scala 156:36:@65758.4]
  wire  _T_1593; // @[SpatialBlocks.scala 156:78:@65759.4]
  wire  _T_1605; // @[package.scala 96:25:@65983.4 package.scala 96:25:@65984.4]
  _ _ ( // @[Math.scala 720:24:@61152.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  b550_chain b550_chain ( // @[sm_x653_outr_Reduce.scala 85:30:@61160.4]
    .clock(b550_chain_clock),
    .reset(b550_chain_reset),
    .io_rPort_5_output_0(b550_chain_io_rPort_5_output_0),
    .io_rPort_4_output_0(b550_chain_io_rPort_4_output_0),
    .io_rPort_3_output_0(b550_chain_io_rPort_3_output_0),
    .io_rPort_2_output_0(b550_chain_io_rPort_2_output_0),
    .io_rPort_1_output_0(b550_chain_io_rPort_1_output_0),
    .io_rPort_0_output_0(b550_chain_io_rPort_0_output_0),
    .io_wPort_0_data_0(b550_chain_io_wPort_0_data_0),
    .io_wPort_0_reset(b550_chain_io_wPort_0_reset),
    .io_wPort_0_en_0(b550_chain_io_wPort_0_en_0),
    .io_sEn_0(b550_chain_io_sEn_0),
    .io_sEn_1(b550_chain_io_sEn_1),
    .io_sEn_2(b550_chain_io_sEn_2),
    .io_sEn_3(b550_chain_io_sEn_3),
    .io_sEn_4(b550_chain_io_sEn_4),
    .io_sEn_5(b550_chain_io_sEn_5),
    .io_sEn_6(b550_chain_io_sEn_6),
    .io_sDone_0(b550_chain_io_sDone_0),
    .io_sDone_1(b550_chain_io_sDone_1),
    .io_sDone_2(b550_chain_io_sDone_2),
    .io_sDone_3(b550_chain_io_sDone_3),
    .io_sDone_4(b550_chain_io_sDone_4),
    .io_sDone_5(b550_chain_io_sDone_5),
    .io_sDone_6(b550_chain_io_sDone_6)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@61224.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  _ __1 ( // @[Math.scala 720:24:@61236.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  _ __2 ( // @[Math.scala 720:24:@61247.4]
    .io_b(__2_io_b),
    .io_result(__2_io_result)
  );
  _ __3 ( // @[Math.scala 720:24:@61258.4]
    .io_b(__3_io_b),
    .io_result(__3_io_result)
  );
  _ __4 ( // @[Math.scala 720:24:@61269.4]
    .io_b(__4_io_b),
    .io_result(__4_io_result)
  );
  _ __5 ( // @[Math.scala 720:24:@61280.4]
    .io_b(__5_io_b),
    .io_result(__5_io_result)
  );
  _ __6 ( // @[Math.scala 720:24:@61291.4]
    .io_b(__6_io_b),
    .io_result(__6_io_result)
  );
  b552_chain b552_chain ( // @[sm_x653_outr_Reduce.scala 94:30:@61300.4]
    .clock(b552_chain_clock),
    .reset(b552_chain_reset),
    .io_rPort_4_output_0(b552_chain_io_rPort_4_output_0),
    .io_rPort_3_output_0(b552_chain_io_rPort_3_output_0),
    .io_rPort_1_output_0(b552_chain_io_rPort_1_output_0),
    .io_rPort_0_output_0(b552_chain_io_rPort_0_output_0),
    .io_wPort_0_data_0(b552_chain_io_wPort_0_data_0),
    .io_wPort_0_reset(b552_chain_io_wPort_0_reset),
    .io_wPort_0_en_0(b552_chain_io_wPort_0_en_0),
    .io_sEn_0(b552_chain_io_sEn_0),
    .io_sEn_1(b552_chain_io_sEn_1),
    .io_sEn_2(b552_chain_io_sEn_2),
    .io_sEn_3(b552_chain_io_sEn_3),
    .io_sEn_4(b552_chain_io_sEn_4),
    .io_sEn_5(b552_chain_io_sEn_5),
    .io_sEn_6(b552_chain_io_sEn_6),
    .io_sDone_0(b552_chain_io_sDone_0),
    .io_sDone_1(b552_chain_io_sDone_1),
    .io_sDone_2(b552_chain_io_sDone_2),
    .io_sDone_3(b552_chain_io_sDone_3),
    .io_sDone_4(b552_chain_io_sDone_4),
    .io_sDone_5(b552_chain_io_sDone_5),
    .io_sDone_6(b552_chain_io_sDone_6)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@61364.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x554_tmp_0 x554_tmp_0 ( // @[m_x554_tmp_0.scala 28:22:@61379.4]
    .clock(x554_tmp_0_clock),
    .reset(x554_tmp_0_reset),
    .io_rPort_0_ofs_0(x554_tmp_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x554_tmp_0_io_rPort_0_en_0),
    .io_rPort_0_output_0(x554_tmp_0_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(x554_tmp_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x554_tmp_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x554_tmp_0_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(x554_tmp_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x554_tmp_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x554_tmp_0_io_wPort_0_en_0),
    .io_sEn_0(x554_tmp_0_io_sEn_0),
    .io_sEn_1(x554_tmp_0_io_sEn_1),
    .io_sEn_2(x554_tmp_0_io_sEn_2),
    .io_sEn_3(x554_tmp_0_io_sEn_3),
    .io_sEn_4(x554_tmp_0_io_sEn_4),
    .io_sEn_5(x554_tmp_0_io_sEn_5),
    .io_sDone_0(x554_tmp_0_io_sDone_0),
    .io_sDone_1(x554_tmp_0_io_sDone_1),
    .io_sDone_2(x554_tmp_0_io_sDone_2),
    .io_sDone_3(x554_tmp_0_io_sDone_3),
    .io_sDone_4(x554_tmp_0_io_sDone_4),
    .io_sDone_5(x554_tmp_0_io_sDone_5)
  );
  x554_tmp_0 x555_tmp_1 ( // @[m_x555_tmp_1.scala 28:22:@61426.4]
    .clock(x555_tmp_1_clock),
    .reset(x555_tmp_1_reset),
    .io_rPort_0_ofs_0(x555_tmp_1_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x555_tmp_1_io_rPort_0_en_0),
    .io_rPort_0_output_0(x555_tmp_1_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(x555_tmp_1_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x555_tmp_1_io_wPort_1_data_0),
    .io_wPort_1_en_0(x555_tmp_1_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(x555_tmp_1_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x555_tmp_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(x555_tmp_1_io_wPort_0_en_0),
    .io_sEn_0(x555_tmp_1_io_sEn_0),
    .io_sEn_1(x555_tmp_1_io_sEn_1),
    .io_sEn_2(x555_tmp_1_io_sEn_2),
    .io_sEn_3(x555_tmp_1_io_sEn_3),
    .io_sEn_4(x555_tmp_1_io_sEn_4),
    .io_sEn_5(x555_tmp_1_io_sEn_5),
    .io_sDone_0(x555_tmp_1_io_sDone_0),
    .io_sDone_1(x555_tmp_1_io_sDone_1),
    .io_sDone_2(x555_tmp_1_io_sDone_2),
    .io_sDone_3(x555_tmp_1_io_sDone_3),
    .io_sDone_4(x555_tmp_1_io_sDone_4),
    .io_sDone_5(x555_tmp_1_io_sDone_5)
  );
  x554_tmp_0 x556_tmp_2 ( // @[m_x556_tmp_2.scala 28:22:@61473.4]
    .clock(x556_tmp_2_clock),
    .reset(x556_tmp_2_reset),
    .io_rPort_0_ofs_0(x556_tmp_2_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x556_tmp_2_io_rPort_0_en_0),
    .io_rPort_0_output_0(x556_tmp_2_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(x556_tmp_2_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x556_tmp_2_io_wPort_1_data_0),
    .io_wPort_1_en_0(x556_tmp_2_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(x556_tmp_2_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x556_tmp_2_io_wPort_0_data_0),
    .io_wPort_0_en_0(x556_tmp_2_io_wPort_0_en_0),
    .io_sEn_0(x556_tmp_2_io_sEn_0),
    .io_sEn_1(x556_tmp_2_io_sEn_1),
    .io_sEn_2(x556_tmp_2_io_sEn_2),
    .io_sEn_3(x556_tmp_2_io_sEn_3),
    .io_sEn_4(x556_tmp_2_io_sEn_4),
    .io_sEn_5(x556_tmp_2_io_sEn_5),
    .io_sDone_0(x556_tmp_2_io_sDone_0),
    .io_sDone_1(x556_tmp_2_io_sDone_1),
    .io_sDone_2(x556_tmp_2_io_sDone_2),
    .io_sDone_3(x556_tmp_2_io_sDone_3),
    .io_sDone_4(x556_tmp_2_io_sDone_4),
    .io_sDone_5(x556_tmp_2_io_sDone_5)
  );
  x557_tmp_3 x557_tmp_3 ( // @[m_x557_tmp_3.scala 28:22:@61520.4]
    .clock(x557_tmp_3_clock),
    .reset(x557_tmp_3_reset),
    .io_rPort_0_ofs_0(x557_tmp_3_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x557_tmp_3_io_rPort_0_en_0),
    .io_rPort_0_output_0(x557_tmp_3_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(x557_tmp_3_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x557_tmp_3_io_wPort_1_data_0),
    .io_wPort_1_en_0(x557_tmp_3_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(x557_tmp_3_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x557_tmp_3_io_wPort_0_data_0),
    .io_wPort_0_en_0(x557_tmp_3_io_wPort_0_en_0),
    .io_sEn_0(x557_tmp_3_io_sEn_0),
    .io_sEn_1(x557_tmp_3_io_sEn_1),
    .io_sEn_2(x557_tmp_3_io_sEn_2),
    .io_sEn_3(x557_tmp_3_io_sEn_3),
    .io_sEn_4(x557_tmp_3_io_sEn_4),
    .io_sEn_5(x557_tmp_3_io_sEn_5),
    .io_sDone_0(x557_tmp_3_io_sDone_0),
    .io_sDone_1(x557_tmp_3_io_sDone_1),
    .io_sDone_2(x557_tmp_3_io_sDone_2),
    .io_sDone_3(x557_tmp_3_io_sDone_3),
    .io_sDone_4(x557_tmp_3_io_sDone_4),
    .io_sDone_5(x557_tmp_3_io_sDone_5)
  );
  x558_tmp_4 x558_tmp_4 ( // @[m_x558_tmp_4.scala 28:22:@61567.4]
    .clock(x558_tmp_4_clock),
    .reset(x558_tmp_4_reset),
    .io_rPort_0_ofs_0(x558_tmp_4_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x558_tmp_4_io_rPort_0_en_0),
    .io_rPort_0_output_0(x558_tmp_4_io_rPort_0_output_0),
    .io_wPort_1_ofs_0(x558_tmp_4_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x558_tmp_4_io_wPort_1_data_0),
    .io_wPort_1_en_0(x558_tmp_4_io_wPort_1_en_0),
    .io_wPort_0_ofs_0(x558_tmp_4_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x558_tmp_4_io_wPort_0_data_0),
    .io_wPort_0_en_0(x558_tmp_4_io_wPort_0_en_0),
    .io_sEn_0(x558_tmp_4_io_sEn_0),
    .io_sEn_1(x558_tmp_4_io_sEn_1),
    .io_sEn_2(x558_tmp_4_io_sEn_2),
    .io_sEn_3(x558_tmp_4_io_sEn_3),
    .io_sEn_4(x558_tmp_4_io_sEn_4),
    .io_sEn_5(x558_tmp_4_io_sEn_5),
    .io_sEn_6(x558_tmp_4_io_sEn_6),
    .io_sDone_0(x558_tmp_4_io_sDone_0),
    .io_sDone_1(x558_tmp_4_io_sDone_1),
    .io_sDone_2(x558_tmp_4_io_sDone_2),
    .io_sDone_3(x558_tmp_4_io_sDone_3),
    .io_sDone_4(x558_tmp_4_io_sDone_4),
    .io_sDone_5(x558_tmp_4_io_sDone_5),
    .io_sDone_6(x558_tmp_4_io_sDone_6)
  );
  x549_ctrchain x560_ctrchain ( // @[SpatialBlocks.scala 37:22:@61616.4]
    .clock(x560_ctrchain_clock),
    .reset(x560_ctrchain_reset),
    .io_input_reset(x560_ctrchain_io_input_reset),
    .io_input_enable(x560_ctrchain_io_input_enable),
    .io_output_counts_0(x560_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x560_ctrchain_io_output_oobs_0),
    .io_output_done(x560_ctrchain_io_output_done)
  );
  x579_inr_Foreach_sm x579_inr_Foreach_sm ( // @[sm_x579_inr_Foreach.scala 35:18:@61669.4]
    .clock(x579_inr_Foreach_sm_clock),
    .reset(x579_inr_Foreach_sm_reset),
    .io_enable(x579_inr_Foreach_sm_io_enable),
    .io_done(x579_inr_Foreach_sm_io_done),
    .io_ctrDone(x579_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x579_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x579_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x579_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x579_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x579_inr_Foreach_sm_io_backpressure),
    .io_break(x579_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@61698.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@61707.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@61717.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@61759.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@61767.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x579_inr_Foreach_kernelx579_inr_Foreach_concrete1 x579_inr_Foreach_kernelx579_inr_Foreach_concrete1 ( // @[sm_x579_inr_Foreach.scala 180:24:@61801.4]
    .clock(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_clock),
    .reset(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_reset),
    .io_in_x555_tmp_1_wPort_0_ofs_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_ofs_0),
    .io_in_x555_tmp_1_wPort_0_data_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_data_0),
    .io_in_x555_tmp_1_wPort_0_en_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_en_0),
    .io_in_x555_tmp_1_sEn_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_sEn_0),
    .io_in_x555_tmp_1_sDone_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_sDone_0),
    .io_in_b550_number(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b550_number),
    .io_in_x472_A_sram_1_rPort_0_ofs_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0),
    .io_in_x472_A_sram_1_rPort_0_en_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_en_0),
    .io_in_x472_A_sram_1_rPort_0_output_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_output_0),
    .io_in_b542_number(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b542_number),
    .io_in_x471_A_sram_0_rPort_0_ofs_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0),
    .io_in_x471_A_sram_0_rPort_0_en_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_en_0),
    .io_in_x471_A_sram_0_rPort_0_output_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_output_0),
    .io_in_x554_tmp_0_wPort_0_ofs_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_ofs_0),
    .io_in_x554_tmp_0_wPort_0_data_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_data_0),
    .io_in_x554_tmp_0_wPort_0_en_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_en_0),
    .io_in_x554_tmp_0_sEn_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_sEn_0),
    .io_in_x554_tmp_0_sDone_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_sDone_0),
    .io_in_x558_tmp_4_wPort_0_ofs_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_ofs_0),
    .io_in_x558_tmp_4_wPort_0_data_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_data_0),
    .io_in_x558_tmp_4_wPort_0_en_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_en_0),
    .io_in_x558_tmp_4_sEn_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_0),
    .io_in_x558_tmp_4_sDone_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_0),
    .io_in_b552(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b552),
    .io_in_x557_tmp_3_wPort_0_ofs_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_ofs_0),
    .io_in_x557_tmp_3_wPort_0_data_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_data_0),
    .io_in_x557_tmp_3_wPort_0_en_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_en_0),
    .io_in_x557_tmp_3_sEn_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_sEn_0),
    .io_in_x557_tmp_3_sDone_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_sDone_0),
    .io_in_x556_tmp_2_wPort_0_ofs_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_ofs_0),
    .io_in_x556_tmp_2_wPort_0_data_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_data_0),
    .io_in_x556_tmp_2_wPort_0_en_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_en_0),
    .io_in_x556_tmp_2_sEn_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_sEn_0),
    .io_in_x556_tmp_2_sDone_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_sDone_0),
    .io_in_b543(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b543),
    .io_sigsIn_done(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_datapathEn(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_rr)
  );
  x580_r_0 x580_r_0 ( // @[m_x580_r_0.scala 28:22:@62245.4]
    .clock(x580_r_0_clock),
    .reset(x580_r_0_reset),
    .io_rPort_1_en_0(x580_r_0_io_rPort_1_en_0),
    .io_rPort_1_output_0(x580_r_0_io_rPort_1_output_0),
    .io_rPort_0_en_0(x580_r_0_io_rPort_0_en_0),
    .io_rPort_0_output_0(x580_r_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(x580_r_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x580_r_0_io_wPort_0_en_0),
    .io_sEn_0(x580_r_0_io_sEn_0),
    .io_sEn_1(x580_r_0_io_sEn_1),
    .io_sEn_2(x580_r_0_io_sEn_2),
    .io_sDone_0(x580_r_0_io_sDone_0),
    .io_sDone_1(x580_r_0_io_sDone_1),
    .io_sDone_2(x580_r_0_io_sDone_2)
  );
  x593_inr_UnitPipe_sm x593_inr_UnitPipe_sm ( // @[sm_x593_inr_UnitPipe.scala 33:18:@62320.4]
    .clock(x593_inr_UnitPipe_sm_clock),
    .reset(x593_inr_UnitPipe_sm_reset),
    .io_enable(x593_inr_UnitPipe_sm_io_enable),
    .io_done(x593_inr_UnitPipe_sm_io_done),
    .io_ctrDone(x593_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x593_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x593_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x593_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x593_inr_UnitPipe_sm_io_backpressure),
    .io_break(x593_inr_UnitPipe_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@62353.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@62363.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@62399.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@62407.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1 x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1 ( // @[sm_x593_inr_UnitPipe.scala 134:24:@62436.4]
    .clock(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_clock),
    .reset(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_reset),
    .io_in_x555_tmp_1_rPort_0_en_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_rPort_0_en_0),
    .io_in_x555_tmp_1_rPort_0_output_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_rPort_0_output_0),
    .io_in_x555_tmp_1_sEn_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_1),
    .io_in_x555_tmp_1_sDone_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_1),
    .io_in_x554_tmp_0_rPort_0_en_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_rPort_0_en_0),
    .io_in_x554_tmp_0_rPort_0_output_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_rPort_0_output_0),
    .io_in_x554_tmp_0_sEn_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_1),
    .io_in_x554_tmp_0_sDone_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_1),
    .io_in_x558_tmp_4_sEn_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_1),
    .io_in_x558_tmp_4_sDone_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_1),
    .io_in_x557_tmp_3_sEn_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_1),
    .io_in_x557_tmp_3_sDone_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_1),
    .io_in_x580_r_0_wPort_0_data_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_wPort_0_data_0),
    .io_in_x580_r_0_wPort_0_en_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_wPort_0_en_0),
    .io_in_x580_r_0_sEn_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_sEn_0),
    .io_in_x580_r_0_sDone_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_sDone_0),
    .io_in_x556_tmp_2_rPort_0_en_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_rPort_0_en_0),
    .io_in_x556_tmp_2_rPort_0_output_0(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_rPort_0_output_0),
    .io_in_x556_tmp_2_sEn_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_1),
    .io_in_x556_tmp_2_sDone_1(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_1),
    .io_sigsIn_done(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_done),
    .io_sigsIn_datapathEn(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_break),
    .io_rr(x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_rr)
  );
  x594_force_0 x594_force_0 ( // @[m_x594_force_0.scala 27:22:@62880.4]
    .clock(x594_force_0_clock),
    .reset(x594_force_0_reset),
    .io_rPort_0_en_0(x594_force_0_io_rPort_0_en_0),
    .io_rPort_0_output_0(x594_force_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(x594_force_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x594_force_0_io_wPort_0_en_0),
    .io_sEn_0(x594_force_0_io_sEn_0),
    .io_sEn_1(x594_force_0_io_sEn_1),
    .io_sDone_0(x594_force_0_io_sDone_0),
    .io_sDone_1(x594_force_0_io_sDone_1)
  );
  x595_reg x595_reg ( // @[m_x595_reg.scala 28:22:@62910.4]
    .clock(x595_reg_clock),
    .reset(x595_reg_reset),
    .io_rPort_1_output_0(x595_reg_io_rPort_1_output_0),
    .io_rPort_0_output_0(x595_reg_io_rPort_0_output_0),
    .io_wPort_0_data_0(x595_reg_io_wPort_0_data_0),
    .io_wPort_0_reset(x595_reg_io_wPort_0_reset),
    .io_wPort_0_en_0(x595_reg_io_wPort_0_en_0),
    .io_sEn_0(x595_reg_io_sEn_0),
    .io_sEn_1(x595_reg_io_sEn_1),
    .io_sDone_0(x595_reg_io_sDone_0),
    .io_sDone_1(x595_reg_io_sDone_1)
  );
  x596_reg x596_reg ( // @[m_x596_reg.scala 27:22:@62947.4]
    .clock(x596_reg_clock),
    .reset(x596_reg_reset),
    .io_rPort_0_output_0(x596_reg_io_rPort_0_output_0),
    .io_wPort_0_data_0(x596_reg_io_wPort_0_data_0),
    .io_wPort_0_reset(x596_reg_io_wPort_0_reset),
    .io_wPort_0_en_0(x596_reg_io_wPort_0_en_0),
    .io_sEn_0(x596_reg_io_sEn_0),
    .io_sEn_1(x596_reg_io_sEn_1),
    .io_sDone_0(x596_reg_io_sDone_0),
    .io_sDone_1(x596_reg_io_sDone_1)
  );
  x536_inr_Foreach_sm x605_inr_UnitPipe_sm ( // @[sm_x605_inr_UnitPipe.scala 33:18:@63013.4]
    .clock(x605_inr_UnitPipe_sm_clock),
    .reset(x605_inr_UnitPipe_sm_reset),
    .io_enable(x605_inr_UnitPipe_sm_io_enable),
    .io_done(x605_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x605_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x605_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x605_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x605_inr_UnitPipe_sm_io_ctrInc),
    .io_ctrRst(x605_inr_UnitPipe_sm_io_ctrRst),
    .io_parentAck(x605_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x605_inr_UnitPipe_sm_io_backpressure),
    .io_break(x605_inr_UnitPipe_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_11 ( // @[package.scala 93:22:@63046.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper RetimeWrapper_12 ( // @[package.scala 93:22:@63056.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper RetimeWrapper_13 ( // @[package.scala 93:22:@63092.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@63100.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1 x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1 ( // @[sm_x605_inr_UnitPipe.scala 129:24:@63129.4]
    .clock(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_clock),
    .reset(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_reset),
    .io_in_x555_tmp_1_sEn_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_2),
    .io_in_x555_tmp_1_sDone_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_2),
    .io_in_x554_tmp_0_sEn_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_2),
    .io_in_x554_tmp_0_sDone_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_2),
    .io_in_x558_tmp_4_sEn_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_2),
    .io_in_x558_tmp_4_sDone_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_2),
    .io_in_x557_tmp_3_sEn_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_2),
    .io_in_x557_tmp_3_sDone_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_2),
    .io_in_x580_r_0_rPort_0_en_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_rPort_0_en_0),
    .io_in_x580_r_0_rPort_0_output_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_rPort_0_output_0),
    .io_in_x580_r_0_sEn_1(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_sEn_1),
    .io_in_x580_r_0_sDone_1(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_sDone_1),
    .io_in_x595_reg_wPort_0_data_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_data_0),
    .io_in_x595_reg_wPort_0_reset(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_reset),
    .io_in_x595_reg_wPort_0_en_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_en_0),
    .io_in_x595_reg_reset(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_reset),
    .io_in_x595_reg_sEn_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_sEn_0),
    .io_in_x595_reg_sDone_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_sDone_0),
    .io_in_x556_tmp_2_sEn_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_2),
    .io_in_x556_tmp_2_sDone_2(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_2),
    .io_in_x596_reg_wPort_0_data_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_data_0),
    .io_in_x596_reg_wPort_0_reset(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_reset),
    .io_in_x596_reg_wPort_0_en_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_en_0),
    .io_in_x596_reg_reset(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_reset),
    .io_in_x596_reg_sEn_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_sEn_0),
    .io_in_x596_reg_sDone_0(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_sDone_0),
    .io_sigsIn_done(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_done),
    .io_sigsIn_datapathEn(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_break),
    .io_rr(x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_rr)
  );
  x621_inr_Switch_sm x621_inr_Switch_sm ( // @[sm_x621_inr_Switch.scala 33:18:@63732.4]
    .clock(x621_inr_Switch_sm_clock),
    .reset(x621_inr_Switch_sm_reset),
    .io_enable(x621_inr_Switch_sm_io_enable),
    .io_done(x621_inr_Switch_sm_io_done),
    .io_parentAck(x621_inr_Switch_sm_io_parentAck),
    .io_backpressure(x621_inr_Switch_sm_io_backpressure),
    .io_doneIn_0(x621_inr_Switch_sm_io_doneIn_0),
    .io_doneIn_1(x621_inr_Switch_sm_io_doneIn_1),
    .io_childAck_0(x621_inr_Switch_sm_io_childAck_0),
    .io_childAck_1(x621_inr_Switch_sm_io_childAck_1),
    .io_selectsIn_0(x621_inr_Switch_sm_io_selectsIn_0),
    .io_selectsIn_1(x621_inr_Switch_sm_io_selectsIn_1),
    .io_selectsOut_0(x621_inr_Switch_sm_io_selectsOut_0),
    .io_selectsOut_1(x621_inr_Switch_sm_io_selectsOut_1)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@63769.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 ( // @[package.scala 93:22:@63779.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper RetimeWrapper_17 ( // @[package.scala 93:22:@63821.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 ( // @[package.scala 93:22:@63829.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  x621_inr_Switch_kernelx621_inr_Switch_concrete1 x621_inr_Switch_kernelx621_inr_Switch_concrete1 ( // @[sm_x621_inr_Switch.scala 132:24:@63858.4]
    .clock(x621_inr_Switch_kernelx621_inr_Switch_concrete1_clock),
    .reset(x621_inr_Switch_kernelx621_inr_Switch_concrete1_reset),
    .io_in_x555_tmp_1_sEn_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x555_tmp_1_sEn_3),
    .io_in_x555_tmp_1_sDone_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x555_tmp_1_sDone_3),
    .io_in_x554_tmp_0_sEn_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x554_tmp_0_sEn_3),
    .io_in_x554_tmp_0_sDone_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x554_tmp_0_sDone_3),
    .io_in_x558_tmp_4_sEn_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x558_tmp_4_sEn_3),
    .io_in_x558_tmp_4_sDone_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x558_tmp_4_sDone_3),
    .io_in_x736_rd_x596(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x736_rd_x596),
    .io_in_x557_tmp_3_sEn_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x557_tmp_3_sEn_3),
    .io_in_x557_tmp_3_sDone_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x557_tmp_3_sDone_3),
    .io_in_x580_r_0_rPort_1_en_0(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_rPort_1_en_0),
    .io_in_x580_r_0_rPort_1_output_0(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_rPort_1_output_0),
    .io_in_x580_r_0_sEn_2(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_sEn_2),
    .io_in_x580_r_0_sDone_2(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_sDone_2),
    .io_in_x595_reg_rPort_1_output_0(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_rPort_1_output_0),
    .io_in_x595_reg_sEn_1(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_sEn_1),
    .io_in_x595_reg_sDone_1(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_sDone_1),
    .io_in_x556_tmp_2_sEn_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x556_tmp_2_sEn_3),
    .io_in_x556_tmp_2_sDone_3(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x556_tmp_2_sDone_3),
    .io_in_x735_rd_x595(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x735_rd_x595),
    .io_in_x596_reg_sEn_1(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x596_reg_sEn_1),
    .io_in_x596_reg_sDone_1(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x596_reg_sDone_1),
    .io_sigsIn_done(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smSelectsOut_0(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smSelectsOut_0),
    .io_sigsIn_smSelectsOut_1(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smSelectsOut_1),
    .io_sigsIn_smChildAcks_0(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_rr),
    .io_ret_number(x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_ret_number)
  );
  x516_inr_UnitPipe_sm x623_inr_UnitPipe_sm ( // @[sm_x623_inr_UnitPipe.scala 34:18:@64431.4]
    .clock(x623_inr_UnitPipe_sm_clock),
    .reset(x623_inr_UnitPipe_sm_reset),
    .io_enable(x623_inr_UnitPipe_sm_io_enable),
    .io_done(x623_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x623_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x623_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x623_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x623_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x623_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x623_inr_UnitPipe_sm_io_backpressure),
    .io_break(x623_inr_UnitPipe_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_19 ( // @[package.scala 93:22:@64464.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper RetimeWrapper_20 ( // @[package.scala 93:22:@64474.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper RetimeWrapper_21 ( // @[package.scala 93:22:@64510.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper RetimeWrapper_22 ( // @[package.scala 93:22:@64518.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1 x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1 ( // @[sm_x623_inr_UnitPipe.scala 102:24:@64547.4]
    .clock(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_clock),
    .reset(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_reset),
    .io_in_x555_tmp_1_sEn_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_4),
    .io_in_x555_tmp_1_sDone_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_4),
    .io_in_x554_tmp_0_sEn_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_4),
    .io_in_x554_tmp_0_sDone_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_4),
    .io_in_x558_tmp_4_sEn_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_4),
    .io_in_x558_tmp_4_sDone_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_4),
    .io_in_x594_force_0_wPort_0_data_0(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_wPort_0_data_0),
    .io_in_x594_force_0_wPort_0_en_0(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_wPort_0_en_0),
    .io_in_x594_force_0_sEn_0(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_sEn_0),
    .io_in_x594_force_0_sDone_0(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_sDone_0),
    .io_in_x621_inr_Switch_number(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x621_inr_Switch_number),
    .io_in_x557_tmp_3_sEn_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_4),
    .io_in_x557_tmp_3_sDone_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_4),
    .io_in_x556_tmp_2_sEn_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_4),
    .io_in_x556_tmp_2_sDone_4(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_4),
    .io_sigsIn_done(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_done),
    .io_sigsIn_datapathEn(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_break),
    .io_rr(x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_rr)
  );
  x549_ctrchain x625_ctrchain ( // @[SpatialBlocks.scala 37:22:@64967.4]
    .clock(x625_ctrchain_clock),
    .reset(x625_ctrchain_reset),
    .io_input_reset(x625_ctrchain_io_input_reset),
    .io_input_enable(x625_ctrchain_io_input_enable),
    .io_output_counts_0(x625_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x625_ctrchain_io_output_oobs_0),
    .io_output_done(x625_ctrchain_io_output_done)
  );
  x639_inr_Foreach_sm x639_inr_Foreach_sm ( // @[sm_x639_inr_Foreach.scala 33:18:@65020.4]
    .clock(x639_inr_Foreach_sm_clock),
    .reset(x639_inr_Foreach_sm_reset),
    .io_enable(x639_inr_Foreach_sm_io_enable),
    .io_done(x639_inr_Foreach_sm_io_done),
    .io_rst(x639_inr_Foreach_sm_io_rst),
    .io_ctrDone(x639_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x639_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x639_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x639_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x639_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x639_inr_Foreach_sm_io_backpressure),
    .io_break(x639_inr_Foreach_sm_io_break)
  );
  x639_inr_Foreach_iiCtr x639_inr_Foreach_iiCtr ( // @[sm_x639_inr_Foreach.scala 34:21:@65045.4]
    .clock(x639_inr_Foreach_iiCtr_clock),
    .reset(x639_inr_Foreach_iiCtr_reset),
    .io_input_enable(x639_inr_Foreach_iiCtr_io_input_enable),
    .io_input_reset(x639_inr_Foreach_iiCtr_io_input_reset),
    .io_output_issue(x639_inr_Foreach_iiCtr_io_output_issue),
    .io_output_done(x639_inr_Foreach_iiCtr_io_output_done)
  );
  RetimeWrapper RetimeWrapper_23 ( // @[package.scala 93:22:@65049.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper RetimeWrapper_24 ( // @[package.scala 93:22:@65058.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@65068.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper RetimeWrapper_26 ( // @[package.scala 93:22:@65110.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper RetimeWrapper_27 ( // @[package.scala 93:22:@65118.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  x639_inr_Foreach_kernelx639_inr_Foreach_concrete1 x639_inr_Foreach_kernelx639_inr_Foreach_concrete1 ( // @[sm_x639_inr_Foreach.scala 151:24:@65152.4]
    .clock(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_clock),
    .reset(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_reset),
    .io_in_x555_tmp_1_wPort_1_ofs_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_ofs_0),
    .io_in_x555_tmp_1_wPort_1_data_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_data_0),
    .io_in_x555_tmp_1_wPort_1_en_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_en_0),
    .io_in_x555_tmp_1_sEn_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_sEn_5),
    .io_in_x555_tmp_1_sDone_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_sDone_5),
    .io_in_x554_tmp_0_wPort_1_ofs_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_ofs_0),
    .io_in_x554_tmp_0_wPort_1_data_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_data_0),
    .io_in_x554_tmp_0_wPort_1_en_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_en_0),
    .io_in_x554_tmp_0_sEn_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_sEn_5),
    .io_in_x554_tmp_0_sDone_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_sDone_5),
    .io_in_x558_tmp_4_wPort_1_ofs_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_ofs_0),
    .io_in_x558_tmp_4_wPort_1_data_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_data_0),
    .io_in_x558_tmp_4_wPort_1_en_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_en_0),
    .io_in_x558_tmp_4_sEn_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_5),
    .io_in_x558_tmp_4_sDone_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_5),
    .io_in_b552(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_b552),
    .io_in_x594_force_0_rPort_0_en_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_rPort_0_en_0),
    .io_in_x594_force_0_rPort_0_output_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_rPort_0_output_0),
    .io_in_x594_force_0_sEn_1(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_sEn_1),
    .io_in_x594_force_0_sDone_1(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_sDone_1),
    .io_in_x557_tmp_3_rPort_0_ofs_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_ofs_0),
    .io_in_x557_tmp_3_rPort_0_en_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_en_0),
    .io_in_x557_tmp_3_rPort_0_output_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_output_0),
    .io_in_x557_tmp_3_wPort_1_ofs_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_ofs_0),
    .io_in_x557_tmp_3_wPort_1_data_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_data_0),
    .io_in_x557_tmp_3_wPort_1_en_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_en_0),
    .io_in_x557_tmp_3_sEn_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_sEn_5),
    .io_in_x557_tmp_3_sDone_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_sDone_5),
    .io_in_x556_tmp_2_wPort_1_ofs_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_ofs_0),
    .io_in_x556_tmp_2_wPort_1_data_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_data_0),
    .io_in_x556_tmp_2_wPort_1_en_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_en_0),
    .io_in_x556_tmp_2_sEn_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_sEn_5),
    .io_in_x556_tmp_2_sDone_5(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_sDone_5),
    .io_in_b543(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_b543),
    .io_sigsIn_done(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_iiIssue(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_iiIssue),
    .io_sigsIn_datapathEn(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_rr)
  );
  x652_inr_Foreach_sm x652_inr_Foreach_sm ( // @[sm_x652_inr_Foreach.scala 35:18:@65644.4]
    .clock(x652_inr_Foreach_sm_clock),
    .reset(x652_inr_Foreach_sm_reset),
    .io_enable(x652_inr_Foreach_sm_io_enable),
    .io_done(x652_inr_Foreach_sm_io_done),
    .io_doneLatch(x652_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x652_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x652_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x652_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x652_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x652_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x652_inr_Foreach_sm_io_backpressure),
    .io_break(x652_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_28 ( // @[package.scala 93:22:@65673.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper RetimeWrapper_29 ( // @[package.scala 93:22:@65682.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper RetimeWrapper_30 ( // @[package.scala 93:22:@65692.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper RetimeWrapper_31 ( // @[package.scala 93:22:@65733.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper RetimeWrapper_32 ( // @[package.scala 93:22:@65741.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  x652_inr_Foreach_kernelx652_inr_Foreach_concrete1 x652_inr_Foreach_kernelx652_inr_Foreach_concrete1 ( // @[sm_x652_inr_Foreach.scala 123:24:@65775.4]
    .clock(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_clock),
    .reset(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_reset),
    .io_in_b550_number(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_b550_number),
    .io_in_x558_tmp_4_rPort_0_ofs_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_ofs_0),
    .io_in_x558_tmp_4_rPort_0_en_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_en_0),
    .io_in_x558_tmp_4_rPort_0_output_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_output_0),
    .io_in_x558_tmp_4_sEn_6(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_6),
    .io_in_x558_tmp_4_sDone_6(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_6),
    .io_in_x545_accum_1_wPort_0_ofs_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_ofs_0),
    .io_in_x545_accum_1_wPort_0_data_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_data_0),
    .io_in_x545_accum_1_wPort_0_en_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_en_0),
    .io_in_x544_accum_0_rPort_0_ofs_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_ofs_0),
    .io_in_x544_accum_0_rPort_0_en_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_en_0),
    .io_in_x544_accum_0_rPort_0_output_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_output_0),
    .io_in_x544_accum_0_wPort_0_ofs_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_ofs_0),
    .io_in_x544_accum_0_wPort_0_data_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_data_0),
    .io_in_x544_accum_0_wPort_0_en_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_en_0),
    .io_in_b543(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_b543),
    .io_sigsIn_done(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_datapathEn(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_rr)
  );
  RetimeWrapper RetimeWrapper_33 ( // @[package.scala 93:22:@65978.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  assign b552 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x653_outr_Reduce.scala 93:18:@61299.4]
  assign b552_chain_read_1 = b552_chain_io_rPort_0_output_0; // @[sm_x653_outr_Reduce.scala 96:61:@61373.4]
  assign b552_chain_read_2 = b552_chain_io_rPort_1_output_0; // @[sm_x653_outr_Reduce.scala 97:61:@61374.4]
  assign b552_chain_read_4 = b552_chain_io_rPort_3_output_0; // @[sm_x653_outr_Reduce.scala 99:61:@61376.4]
  assign b552_chain_read_5 = b552_chain_io_rPort_4_output_0; // @[sm_x653_outr_Reduce.scala 100:61:@61377.4]
  assign _T_897 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@61703.4 package.scala 96:25:@61704.4]
  assign _T_901 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@61712.4 package.scala 96:25:@61713.4]
  assign _T_905 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@61722.4 package.scala 96:25:@61723.4]
  assign x579_inr_Foreach_mySignalsIn_mask = b552 & io_in_b543; // @[sm_x653_outr_Reduce.scala 119:81:@61736.4]
  assign _T_922 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@61764.4 package.scala 96:25:@61765.4]
  assign _T_928 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@61772.4 package.scala 96:25:@61773.4]
  assign _T_931 = ~ _T_928; // @[SpatialBlocks.scala 137:99:@61775.4]
  assign _T_933 = x579_inr_Foreach_sm_io_datapathEn & x579_inr_Foreach_mySignalsIn_mask; // @[SpatialBlocks.scala 156:36:@61784.4]
  assign _T_934 = ~ x579_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 156:78:@61785.4]
  assign _T_1002 = x593_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@62348.4]
  assign _T_1008 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@62358.4 package.scala 96:25:@62359.4]
  assign _T_1012 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@62368.4 package.scala 96:25:@62369.4]
  assign x593_inr_UnitPipe_mySignalsIn_mask = b552_chain_read_1 & io_in_b543; // @[sm_x653_outr_Reduce.scala 131:60:@62381.4]
  assign _T_1029 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@62404.4 package.scala 96:25:@62405.4]
  assign _T_1035 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@62412.4 package.scala 96:25:@62413.4]
  assign _T_1038 = ~ _T_1035; // @[SpatialBlocks.scala 137:99:@62415.4]
  assign _T_1109 = x605_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@63041.4]
  assign _T_1115 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@63051.4 package.scala 96:25:@63052.4]
  assign _T_1119 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@63061.4 package.scala 96:25:@63062.4]
  assign x605_inr_UnitPipe_mySignalsIn_mask = b552_chain_read_2 & io_in_b543; // @[sm_x653_outr_Reduce.scala 145:60:@63074.4]
  assign _T_1136 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@63097.4 package.scala 96:25:@63098.4]
  assign _T_1142 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@63105.4 package.scala 96:25:@63106.4]
  assign _T_1145 = ~ _T_1142; // @[SpatialBlocks.scala 137:99:@63108.4]
  assign _T_1243 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@63774.4 package.scala 96:25:@63775.4]
  assign _T_1247 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@63784.4 package.scala 96:25:@63785.4]
  assign _T_1265 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@63826.4 package.scala 96:25:@63827.4]
  assign _T_1271 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@63834.4 package.scala 96:25:@63835.4]
  assign _T_1274 = ~ _T_1271; // @[SpatialBlocks.scala 137:99:@63837.4]
  assign _T_1342 = x623_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@64459.4]
  assign _T_1348 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@64469.4 package.scala 96:25:@64470.4]
  assign _T_1352 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@64479.4 package.scala 96:25:@64480.4]
  assign x623_inr_UnitPipe_mySignalsIn_mask = b552_chain_read_4 & io_in_b543; // @[sm_x653_outr_Reduce.scala 181:60:@64492.4]
  assign _T_1369 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@64515.4 package.scala 96:25:@64516.4]
  assign _T_1375 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@64523.4 package.scala 96:25:@64524.4]
  assign _T_1378 = ~ _T_1375; // @[SpatialBlocks.scala 137:99:@64526.4]
  assign _T_1450 = RetimeWrapper_23_io_out; // @[package.scala 96:25:@65054.4 package.scala 96:25:@65055.4]
  assign _T_1454 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@65063.4 package.scala 96:25:@65064.4]
  assign _T_1458 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@65073.4 package.scala 96:25:@65074.4]
  assign x639_inr_Foreach_mySignalsIn_mask = b552_chain_read_5 & io_in_b543; // @[sm_x653_outr_Reduce.scala 196:94:@65087.4]
  assign _T_1475 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@65115.4 package.scala 96:25:@65116.4]
  assign _T_1481 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@65123.4 package.scala 96:25:@65124.4]
  assign _T_1484 = ~ _T_1481; // @[SpatialBlocks.scala 137:99:@65126.4]
  assign _T_1486 = x639_inr_Foreach_sm_io_datapathEn & x639_inr_Foreach_mySignalsIn_mask; // @[SpatialBlocks.scala 156:36:@65135.4]
  assign _T_1487 = ~ x639_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 156:78:@65136.4]
  assign _T_1490 = ~ x639_inr_Foreach_mySignalsIn_mask; // @[SpatialBlocks.scala 157:128:@65142.4]
  assign x639_inr_Foreach_mySignalsIn_iiDone = x639_inr_Foreach_iiCtr_io_output_done | _T_1490; // @[SpatialBlocks.scala 157:126:@65143.4]
  assign _T_1556 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@65678.4 package.scala 96:25:@65679.4]
  assign _T_1560 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@65687.4 package.scala 96:25:@65688.4]
  assign _T_1564 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@65697.4 package.scala 96:25:@65698.4]
  assign _T_1581 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@65738.4 package.scala 96:25:@65739.4]
  assign _T_1587 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@65746.4 package.scala 96:25:@65747.4]
  assign _T_1590 = ~ _T_1587; // @[SpatialBlocks.scala 137:99:@65749.4]
  assign _T_1592 = x652_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 156:36:@65758.4]
  assign _T_1593 = ~ x652_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 156:78:@65759.4]
  assign _T_1605 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@65983.4 package.scala 96:25:@65984.4]
  assign io_in_x472_A_sram_1_rPort_0_ofs_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@62108.4]
  assign io_in_x472_A_sram_1_rPort_0_en_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@62107.4]
  assign io_in_x471_A_sram_0_rPort_0_ofs_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@62114.4]
  assign io_in_x471_A_sram_0_rPort_0_en_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@62113.4]
  assign io_in_x545_accum_1_wPort_0_ofs_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@65935.4]
  assign io_in_x545_accum_1_wPort_0_data_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@65934.4]
  assign io_in_x545_accum_1_wPort_0_en_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x545_accum_1_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@65930.4]
  assign io_in_x545_accum_1_sEn_0 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@65986.4]
  assign io_in_x545_accum_1_sDone_0 = io_rr ? _T_1605 : 1'h0; // @[MemInterfaceType.scala 197:17:@65987.4]
  assign io_in_x544_accum_0_rPort_0_ofs_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@65940.4]
  assign io_in_x544_accum_0_rPort_0_en_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@65939.4]
  assign io_in_x544_accum_0_wPort_0_ofs_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@65947.4]
  assign io_in_x544_accum_0_wPort_0_data_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@65946.4]
  assign io_in_x544_accum_0_wPort_0_en_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@65942.4]
  assign io_in_x549_ctrchain_input_reset = x652_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@65774.4]
  assign io_in_x549_ctrchain_input_enable = x652_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 158:42:@65773.4]
  assign io_sigsOut_smDoneIn_0 = x579_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@61782.4]
  assign io_sigsOut_smDoneIn_1 = x593_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 155:56:@62422.4]
  assign io_sigsOut_smDoneIn_2 = x605_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 155:56:@63115.4]
  assign io_sigsOut_smDoneIn_3 = x621_inr_Switch_sm_io_done; // @[SpatialBlocks.scala 155:56:@63844.4]
  assign io_sigsOut_smDoneIn_4 = x623_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 155:56:@64533.4]
  assign io_sigsOut_smDoneIn_5 = x639_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@65133.4]
  assign io_sigsOut_smDoneIn_6 = x652_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@65756.4]
  assign io_sigsOut_smMaskIn_0 = b552 & io_in_b543; // @[SpatialBlocks.scala 155:86:@61783.4]
  assign io_sigsOut_smMaskIn_1 = b552_chain_read_1 & io_in_b543; // @[SpatialBlocks.scala 155:86:@62423.4]
  assign io_sigsOut_smMaskIn_2 = b552_chain_read_2 & io_in_b543; // @[SpatialBlocks.scala 155:86:@63116.4]
  assign io_sigsOut_smMaskIn_4 = b552_chain_read_4 & io_in_b543; // @[SpatialBlocks.scala 155:86:@64534.4]
  assign io_sigsOut_smMaskIn_5 = b552_chain_read_5 & io_in_b543; // @[SpatialBlocks.scala 155:86:@65134.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@61155.4]
  assign b550_chain_clock = clock; // @[:@61161.4]
  assign b550_chain_reset = reset; // @[:@61162.4]
  assign b550_chain_io_wPort_0_data_0 = __io_result; // @[NBuffers.scala 309:54:@61222.4]
  assign b550_chain_io_wPort_0_reset = RetimeWrapper_io_out; // @[NBuffers.scala 312:23:@61231.4]
  assign b550_chain_io_wPort_0_en_0 = io_sigsOut_smDoneIn_0; // @[NBuffers.scala 311:25:@61223.4]
  assign b550_chain_io_sEn_0 = _T_922 & _T_931; // @[NBuffers.scala 302:18:@61715.4]
  assign b550_chain_io_sEn_1 = _T_1029 & _T_1038; // @[NBuffers.scala 302:18:@62361.4]
  assign b550_chain_io_sEn_2 = _T_1136 & _T_1145; // @[NBuffers.scala 302:18:@63054.4]
  assign b550_chain_io_sEn_3 = _T_1265 & _T_1274; // @[NBuffers.scala 302:18:@63777.4]
  assign b550_chain_io_sEn_4 = _T_1369 & _T_1378; // @[NBuffers.scala 302:18:@64472.4]
  assign b550_chain_io_sEn_5 = _T_1475 & _T_1484; // @[NBuffers.scala 302:18:@65066.4]
  assign b550_chain_io_sEn_6 = _T_1581 & _T_1590; // @[NBuffers.scala 302:18:@65690.4]
  assign b550_chain_io_sDone_0 = io_rr ? _T_901 : 1'h0; // @[NBuffers.scala 303:20:@61716.4]
  assign b550_chain_io_sDone_1 = io_rr ? _T_1008 : 1'h0; // @[NBuffers.scala 303:20:@62362.4]
  assign b550_chain_io_sDone_2 = io_rr ? _T_1115 : 1'h0; // @[NBuffers.scala 303:20:@63055.4]
  assign b550_chain_io_sDone_3 = io_rr ? _T_1243 : 1'h0; // @[NBuffers.scala 303:20:@63778.4]
  assign b550_chain_io_sDone_4 = io_rr ? _T_1348 : 1'h0; // @[NBuffers.scala 303:20:@64473.4]
  assign b550_chain_io_sDone_5 = io_rr ? _T_1454 : 1'h0; // @[NBuffers.scala 303:20:@65067.4]
  assign b550_chain_io_sDone_6 = io_rr ? _T_1560 : 1'h0; // @[NBuffers.scala 303:20:@65691.4]
  assign RetimeWrapper_clock = clock; // @[:@61225.4]
  assign RetimeWrapper_reset = reset; // @[:@61226.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@61228.4]
  assign RetimeWrapper_io_in = b550_chain_reset; // @[package.scala 94:16:@61227.4]
  assign __1_io_b = b550_chain_io_rPort_0_output_0; // @[Math.scala 721:17:@61239.4]
  assign __2_io_b = b550_chain_io_rPort_1_output_0; // @[Math.scala 721:17:@61250.4]
  assign __3_io_b = b550_chain_io_rPort_2_output_0; // @[Math.scala 721:17:@61261.4]
  assign __4_io_b = b550_chain_io_rPort_3_output_0; // @[Math.scala 721:17:@61272.4]
  assign __5_io_b = b550_chain_io_rPort_4_output_0; // @[Math.scala 721:17:@61283.4]
  assign __6_io_b = b550_chain_io_rPort_5_output_0; // @[Math.scala 721:17:@61294.4]
  assign b552_chain_clock = clock; // @[:@61301.4]
  assign b552_chain_reset = reset; // @[:@61302.4]
  assign b552_chain_io_wPort_0_data_0 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[NBuffers.scala 308:54:@61362.4]
  assign b552_chain_io_wPort_0_reset = RetimeWrapper_1_io_out; // @[NBuffers.scala 312:23:@61371.4]
  assign b552_chain_io_wPort_0_en_0 = io_sigsOut_smDoneIn_0; // @[NBuffers.scala 311:25:@61363.4]
  assign b552_chain_io_sEn_0 = _T_922 & _T_931; // @[NBuffers.scala 302:18:@61725.4]
  assign b552_chain_io_sEn_1 = _T_1029 & _T_1038; // @[NBuffers.scala 302:18:@62371.4]
  assign b552_chain_io_sEn_2 = _T_1136 & _T_1145; // @[NBuffers.scala 302:18:@63064.4]
  assign b552_chain_io_sEn_3 = _T_1265 & _T_1274; // @[NBuffers.scala 302:18:@63787.4]
  assign b552_chain_io_sEn_4 = _T_1369 & _T_1378; // @[NBuffers.scala 302:18:@64482.4]
  assign b552_chain_io_sEn_5 = _T_1475 & _T_1484; // @[NBuffers.scala 302:18:@65076.4]
  assign b552_chain_io_sEn_6 = _T_1581 & _T_1590; // @[NBuffers.scala 302:18:@65700.4]
  assign b552_chain_io_sDone_0 = io_rr ? _T_905 : 1'h0; // @[NBuffers.scala 303:20:@61726.4]
  assign b552_chain_io_sDone_1 = io_rr ? _T_1012 : 1'h0; // @[NBuffers.scala 303:20:@62372.4]
  assign b552_chain_io_sDone_2 = io_rr ? _T_1119 : 1'h0; // @[NBuffers.scala 303:20:@63065.4]
  assign b552_chain_io_sDone_3 = io_rr ? _T_1247 : 1'h0; // @[NBuffers.scala 303:20:@63788.4]
  assign b552_chain_io_sDone_4 = io_rr ? _T_1352 : 1'h0; // @[NBuffers.scala 303:20:@64483.4]
  assign b552_chain_io_sDone_5 = io_rr ? _T_1458 : 1'h0; // @[NBuffers.scala 303:20:@65077.4]
  assign b552_chain_io_sDone_6 = io_rr ? _T_1564 : 1'h0; // @[NBuffers.scala 303:20:@65701.4]
  assign RetimeWrapper_1_clock = clock; // @[:@61365.4]
  assign RetimeWrapper_1_reset = reset; // @[:@61366.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@61368.4]
  assign RetimeWrapper_1_io_in = b552_chain_reset; // @[package.scala 94:16:@61367.4]
  assign x554_tmp_0_clock = clock; // @[:@61380.4]
  assign x554_tmp_0_reset = reset; // @[:@61381.4]
  assign x554_tmp_0_io_rPort_0_ofs_0 = 2'h0; // @[MemInterfaceType.scala 66:44:@62765.4]
  assign x554_tmp_0_io_rPort_0_en_0 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@62764.4]
  assign x554_tmp_0_io_wPort_1_ofs_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_ofs_0; // @[MemInterfaceType.scala 67:44:@65476.4]
  assign x554_tmp_0_io_wPort_1_data_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_data_0; // @[MemInterfaceType.scala 67:44:@65475.4]
  assign x554_tmp_0_io_wPort_1_en_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_1_en_0; // @[MemInterfaceType.scala 67:44:@65471.4]
  assign x554_tmp_0_io_wPort_0_ofs_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@62139.4]
  assign x554_tmp_0_io_wPort_0_data_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@62138.4]
  assign x554_tmp_0_io_wPort_0_en_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@62134.4]
  assign x554_tmp_0_io_sEn_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_sEn_0; // @[MemInterfaceType.scala 189:41:@62124.4]
  assign x554_tmp_0_io_sEn_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_1; // @[MemInterfaceType.scala 189:41:@62752.4]
  assign x554_tmp_0_io_sEn_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_2; // @[MemInterfaceType.scala 189:41:@63499.4]
  assign x554_tmp_0_io_sEn_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x554_tmp_0_sEn_3; // @[MemInterfaceType.scala 189:41:@64234.4]
  assign x554_tmp_0_io_sEn_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sEn_4; // @[MemInterfaceType.scala 189:41:@64850.4]
  assign x554_tmp_0_io_sEn_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_sEn_5; // @[MemInterfaceType.scala 189:41:@65461.4]
  assign x554_tmp_0_io_sDone_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x554_tmp_0_sDone_0; // @[MemInterfaceType.scala 189:64:@62125.4]
  assign x554_tmp_0_io_sDone_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_1; // @[MemInterfaceType.scala 189:64:@62753.4]
  assign x554_tmp_0_io_sDone_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_2; // @[MemInterfaceType.scala 189:64:@63500.4]
  assign x554_tmp_0_io_sDone_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x554_tmp_0_sDone_3; // @[MemInterfaceType.scala 189:64:@64235.4]
  assign x554_tmp_0_io_sDone_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x554_tmp_0_sDone_4; // @[MemInterfaceType.scala 189:64:@64851.4]
  assign x554_tmp_0_io_sDone_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x554_tmp_0_sDone_5; // @[MemInterfaceType.scala 189:64:@65462.4]
  assign x555_tmp_1_clock = clock; // @[:@61427.4]
  assign x555_tmp_1_reset = reset; // @[:@61428.4]
  assign x555_tmp_1_io_rPort_0_ofs_0 = 2'h1; // @[MemInterfaceType.scala 66:44:@62742.4]
  assign x555_tmp_1_io_rPort_0_en_0 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@62741.4]
  assign x555_tmp_1_io_wPort_1_ofs_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_ofs_0; // @[MemInterfaceType.scala 67:44:@65451.4]
  assign x555_tmp_1_io_wPort_1_data_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_data_0; // @[MemInterfaceType.scala 67:44:@65450.4]
  assign x555_tmp_1_io_wPort_1_en_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_1_en_0; // @[MemInterfaceType.scala 67:44:@65446.4]
  assign x555_tmp_1_io_wPort_0_ofs_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@62102.4]
  assign x555_tmp_1_io_wPort_0_data_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@62101.4]
  assign x555_tmp_1_io_wPort_0_en_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@62097.4]
  assign x555_tmp_1_io_sEn_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_sEn_0; // @[MemInterfaceType.scala 189:41:@62087.4]
  assign x555_tmp_1_io_sEn_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_1; // @[MemInterfaceType.scala 189:41:@62729.4]
  assign x555_tmp_1_io_sEn_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_2; // @[MemInterfaceType.scala 189:41:@63481.4]
  assign x555_tmp_1_io_sEn_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x555_tmp_1_sEn_3; // @[MemInterfaceType.scala 189:41:@64216.4]
  assign x555_tmp_1_io_sEn_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sEn_4; // @[MemInterfaceType.scala 189:41:@64832.4]
  assign x555_tmp_1_io_sEn_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_sEn_5; // @[MemInterfaceType.scala 189:41:@65436.4]
  assign x555_tmp_1_io_sDone_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x555_tmp_1_sDone_0; // @[MemInterfaceType.scala 189:64:@62088.4]
  assign x555_tmp_1_io_sDone_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_1; // @[MemInterfaceType.scala 189:64:@62730.4]
  assign x555_tmp_1_io_sDone_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_2; // @[MemInterfaceType.scala 189:64:@63482.4]
  assign x555_tmp_1_io_sDone_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x555_tmp_1_sDone_3; // @[MemInterfaceType.scala 189:64:@64217.4]
  assign x555_tmp_1_io_sDone_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x555_tmp_1_sDone_4; // @[MemInterfaceType.scala 189:64:@64833.4]
  assign x555_tmp_1_io_sDone_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x555_tmp_1_sDone_5; // @[MemInterfaceType.scala 189:64:@65437.4]
  assign x556_tmp_2_clock = clock; // @[:@61474.4]
  assign x556_tmp_2_reset = reset; // @[:@61475.4]
  assign x556_tmp_2_io_rPort_0_ofs_0 = 2'h2; // @[MemInterfaceType.scala 66:44:@62850.4]
  assign x556_tmp_2_io_rPort_0_en_0 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@62849.4]
  assign x556_tmp_2_io_wPort_1_ofs_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_ofs_0; // @[MemInterfaceType.scala 67:44:@65578.4]
  assign x556_tmp_2_io_wPort_1_data_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_data_0; // @[MemInterfaceType.scala 67:44:@65577.4]
  assign x556_tmp_2_io_wPort_1_en_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_1_en_0; // @[MemInterfaceType.scala 67:44:@65573.4]
  assign x556_tmp_2_io_wPort_0_ofs_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@62215.4]
  assign x556_tmp_2_io_wPort_0_data_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@62214.4]
  assign x556_tmp_2_io_wPort_0_en_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@62210.4]
  assign x556_tmp_2_io_sEn_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_sEn_0; // @[MemInterfaceType.scala 189:41:@62200.4]
  assign x556_tmp_2_io_sEn_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_1; // @[MemInterfaceType.scala 189:41:@62837.4]
  assign x556_tmp_2_io_sEn_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_2; // @[MemInterfaceType.scala 189:41:@63602.4]
  assign x556_tmp_2_io_sEn_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x556_tmp_2_sEn_3; // @[MemInterfaceType.scala 189:41:@64335.4]
  assign x556_tmp_2_io_sEn_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sEn_4; // @[MemInterfaceType.scala 189:41:@64929.4]
  assign x556_tmp_2_io_sEn_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_sEn_5; // @[MemInterfaceType.scala 189:41:@65563.4]
  assign x556_tmp_2_io_sDone_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x556_tmp_2_sDone_0; // @[MemInterfaceType.scala 189:64:@62201.4]
  assign x556_tmp_2_io_sDone_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_1; // @[MemInterfaceType.scala 189:64:@62838.4]
  assign x556_tmp_2_io_sDone_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_2; // @[MemInterfaceType.scala 189:64:@63603.4]
  assign x556_tmp_2_io_sDone_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x556_tmp_2_sDone_3; // @[MemInterfaceType.scala 189:64:@64336.4]
  assign x556_tmp_2_io_sDone_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x556_tmp_2_sDone_4; // @[MemInterfaceType.scala 189:64:@64930.4]
  assign x556_tmp_2_io_sDone_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x556_tmp_2_sDone_5; // @[MemInterfaceType.scala 189:64:@65564.4]
  assign x557_tmp_3_clock = clock; // @[:@61521.4]
  assign x557_tmp_3_reset = reset; // @[:@61522.4]
  assign x557_tmp_3_io_rPort_0_ofs_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@65546.4]
  assign x557_tmp_3_io_rPort_0_en_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@65545.4]
  assign x557_tmp_3_io_wPort_1_ofs_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_ofs_0; // @[MemInterfaceType.scala 67:44:@65553.4]
  assign x557_tmp_3_io_wPort_1_data_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_data_0; // @[MemInterfaceType.scala 67:44:@65552.4]
  assign x557_tmp_3_io_wPort_1_en_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_1_en_0; // @[MemInterfaceType.scala 67:44:@65548.4]
  assign x557_tmp_3_io_wPort_0_ofs_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@62190.4]
  assign x557_tmp_3_io_wPort_0_data_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@62189.4]
  assign x557_tmp_3_io_wPort_0_en_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@62185.4]
  assign x557_tmp_3_io_sEn_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_sEn_0; // @[MemInterfaceType.scala 189:41:@62175.4]
  assign x557_tmp_3_io_sEn_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_1; // @[MemInterfaceType.scala 189:41:@62794.4]
  assign x557_tmp_3_io_sEn_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_2; // @[MemInterfaceType.scala 189:41:@63536.4]
  assign x557_tmp_3_io_sEn_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x557_tmp_3_sEn_3; // @[MemInterfaceType.scala 189:41:@64271.4]
  assign x557_tmp_3_io_sEn_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sEn_4; // @[MemInterfaceType.scala 189:41:@64911.4]
  assign x557_tmp_3_io_sEn_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_sEn_5; // @[MemInterfaceType.scala 189:41:@65533.4]
  assign x557_tmp_3_io_sDone_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x557_tmp_3_sDone_0; // @[MemInterfaceType.scala 189:64:@62176.4]
  assign x557_tmp_3_io_sDone_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_1; // @[MemInterfaceType.scala 189:64:@62795.4]
  assign x557_tmp_3_io_sDone_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_2; // @[MemInterfaceType.scala 189:64:@63537.4]
  assign x557_tmp_3_io_sDone_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x557_tmp_3_sDone_3; // @[MemInterfaceType.scala 189:64:@64272.4]
  assign x557_tmp_3_io_sDone_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x557_tmp_3_sDone_4; // @[MemInterfaceType.scala 189:64:@64912.4]
  assign x557_tmp_3_io_sDone_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_sDone_5; // @[MemInterfaceType.scala 189:64:@65534.4]
  assign x558_tmp_4_clock = clock; // @[:@61568.4]
  assign x558_tmp_4_reset = reset; // @[:@61569.4]
  assign x558_tmp_4_io_rPort_0_ofs_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@65914.4]
  assign x558_tmp_4_io_rPort_0_en_0 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@65913.4]
  assign x558_tmp_4_io_wPort_1_ofs_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_ofs_0; // @[MemInterfaceType.scala 67:44:@65501.4]
  assign x558_tmp_4_io_wPort_1_data_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_data_0; // @[MemInterfaceType.scala 67:44:@65500.4]
  assign x558_tmp_4_io_wPort_1_en_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_1_en_0; // @[MemInterfaceType.scala 67:44:@65496.4]
  assign x558_tmp_4_io_wPort_0_ofs_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@62164.4]
  assign x558_tmp_4_io_wPort_0_data_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@62163.4]
  assign x558_tmp_4_io_wPort_0_en_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@62159.4]
  assign x558_tmp_4_io_sEn_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_0; // @[MemInterfaceType.scala 189:41:@62149.4]
  assign x558_tmp_4_io_sEn_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_1; // @[MemInterfaceType.scala 189:41:@62775.4]
  assign x558_tmp_4_io_sEn_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_2; // @[MemInterfaceType.scala 189:41:@63517.4]
  assign x558_tmp_4_io_sEn_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x558_tmp_4_sEn_3; // @[MemInterfaceType.scala 189:41:@64252.4]
  assign x558_tmp_4_io_sEn_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sEn_4; // @[MemInterfaceType.scala 189:41:@64868.4]
  assign x558_tmp_4_io_sEn_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_5; // @[MemInterfaceType.scala 189:41:@65486.4]
  assign x558_tmp_4_io_sEn_6 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_sEn_6; // @[MemInterfaceType.scala 189:41:@65901.4]
  assign x558_tmp_4_io_sDone_0 = x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_0; // @[MemInterfaceType.scala 189:64:@62150.4]
  assign x558_tmp_4_io_sDone_1 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_1; // @[MemInterfaceType.scala 189:64:@62776.4]
  assign x558_tmp_4_io_sDone_2 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_2; // @[MemInterfaceType.scala 189:64:@63518.4]
  assign x558_tmp_4_io_sDone_3 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x558_tmp_4_sDone_3; // @[MemInterfaceType.scala 189:64:@64253.4]
  assign x558_tmp_4_io_sDone_4 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x558_tmp_4_sDone_4; // @[MemInterfaceType.scala 189:64:@64869.4]
  assign x558_tmp_4_io_sDone_5 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_5; // @[MemInterfaceType.scala 189:64:@65487.4]
  assign x558_tmp_4_io_sDone_6 = x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_sDone_6; // @[MemInterfaceType.scala 189:64:@65902.4]
  assign x560_ctrchain_clock = clock; // @[:@61617.4]
  assign x560_ctrchain_reset = reset; // @[:@61618.4]
  assign x560_ctrchain_io_input_reset = x579_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@61800.4]
  assign x560_ctrchain_io_input_enable = x579_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 158:42:@61799.4]
  assign x579_inr_Foreach_sm_clock = clock; // @[:@61670.4]
  assign x579_inr_Foreach_sm_reset = reset; // @[:@61671.4]
  assign x579_inr_Foreach_sm_io_enable = _T_922 & _T_931; // @[SpatialBlocks.scala 139:18:@61779.4]
  assign x579_inr_Foreach_sm_io_ctrDone = io_rr ? _T_897 : 1'h0; // @[sm_x653_outr_Reduce.scala 112:38:@61706.4]
  assign x579_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@61781.4]
  assign x579_inr_Foreach_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@61753.4]
  assign x579_inr_Foreach_sm_io_break = 1'h0; // @[sm_x653_outr_Reduce.scala 118:36:@61733.4]
  assign RetimeWrapper_2_clock = clock; // @[:@61699.4]
  assign RetimeWrapper_2_reset = reset; // @[:@61700.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@61702.4]
  assign RetimeWrapper_2_io_in = x560_ctrchain_io_output_done; // @[package.scala 94:16:@61701.4]
  assign RetimeWrapper_3_clock = clock; // @[:@61708.4]
  assign RetimeWrapper_3_reset = reset; // @[:@61709.4]
  assign RetimeWrapper_3_io_flow = x579_inr_Foreach_sm_io_backpressure; // @[package.scala 95:18:@61711.4]
  assign RetimeWrapper_3_io_in = x579_inr_Foreach_sm_io_done; // @[package.scala 94:16:@61710.4]
  assign RetimeWrapper_4_clock = clock; // @[:@61718.4]
  assign RetimeWrapper_4_reset = reset; // @[:@61719.4]
  assign RetimeWrapper_4_io_flow = x579_inr_Foreach_sm_io_backpressure; // @[package.scala 95:18:@61721.4]
  assign RetimeWrapper_4_io_in = x579_inr_Foreach_sm_io_done; // @[package.scala 94:16:@61720.4]
  assign RetimeWrapper_5_clock = clock; // @[:@61760.4]
  assign RetimeWrapper_5_reset = reset; // @[:@61761.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@61763.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@61762.4]
  assign RetimeWrapper_6_clock = clock; // @[:@61768.4]
  assign RetimeWrapper_6_reset = reset; // @[:@61769.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@61771.4]
  assign RetimeWrapper_6_io_in = x579_inr_Foreach_sm_io_done; // @[package.scala 94:16:@61770.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_clock = clock; // @[:@61802.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_reset = reset; // @[:@61803.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b550_number = __io_result; // @[sm_x579_inr_Foreach.scala 70:23:@62104.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_output_0 = io_in_x472_A_sram_1_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@62105.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b542_number = io_in_b542_number; // @[sm_x579_inr_Foreach.scala 72:23:@62110.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_output_0 = io_in_x471_A_sram_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@62111.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b552 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x579_inr_Foreach.scala 76:23:@62166.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_in_b543 = io_in_b543; // @[sm_x579_inr_Foreach.scala 79:23:@62217.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_done = x579_inr_Foreach_sm_io_done; // @[sm_x579_inr_Foreach.scala 185:22:@62237.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_933 & _T_934; // @[sm_x579_inr_Foreach.scala 185:22:@62230.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_baseEn = _T_922 & _T_931; // @[sm_x579_inr_Foreach.scala 185:22:@62229.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_break = x579_inr_Foreach_sm_io_break; // @[sm_x579_inr_Foreach.scala 185:22:@62228.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{28{x560_ctrchain_io_output_counts_0[3]}},x560_ctrchain_io_output_counts_0}; // @[sm_x579_inr_Foreach.scala 185:22:@62223.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x560_ctrchain_io_output_oobs_0; // @[sm_x579_inr_Foreach.scala 185:22:@62222.4]
  assign x579_inr_Foreach_kernelx579_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x579_inr_Foreach.scala 184:18:@62218.4]
  assign x580_r_0_clock = clock; // @[:@62246.4]
  assign x580_r_0_reset = reset; // @[:@62247.4]
  assign x580_r_0_io_rPort_1_en_0 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_rPort_1_en_0; // @[MemInterfaceType.scala 66:44:@64301.4]
  assign x580_r_0_io_rPort_0_en_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@63566.4]
  assign x580_r_0_io_wPort_0_data_0 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@62826.4]
  assign x580_r_0_io_wPort_0_en_0 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@62822.4]
  assign x580_r_0_io_sEn_0 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_sEn_0; // @[MemInterfaceType.scala 189:41:@62812.4]
  assign x580_r_0_io_sEn_1 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_sEn_1; // @[MemInterfaceType.scala 189:41:@63554.4]
  assign x580_r_0_io_sEn_2 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_sEn_2; // @[MemInterfaceType.scala 189:41:@64289.4]
  assign x580_r_0_io_sDone_0 = x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x580_r_0_sDone_0; // @[MemInterfaceType.scala 189:64:@62813.4]
  assign x580_r_0_io_sDone_1 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_sDone_1; // @[MemInterfaceType.scala 189:64:@63555.4]
  assign x580_r_0_io_sDone_2 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_sDone_2; // @[MemInterfaceType.scala 189:64:@64290.4]
  assign x593_inr_UnitPipe_sm_clock = clock; // @[:@62321.4]
  assign x593_inr_UnitPipe_sm_reset = reset; // @[:@62322.4]
  assign x593_inr_UnitPipe_sm_io_enable = _T_1029 & _T_1038; // @[SpatialBlocks.scala 139:18:@62419.4]
  assign x593_inr_UnitPipe_sm_io_ctrDone = x593_inr_UnitPipe_sm_io_ctrInc & _T_1005; // @[sm_x653_outr_Reduce.scala 124:39:@62352.4]
  assign x593_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 141:21:@62421.4]
  assign x593_inr_UnitPipe_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@62393.4]
  assign x593_inr_UnitPipe_sm_io_break = 1'h0; // @[sm_x653_outr_Reduce.scala 130:37:@62379.4]
  assign RetimeWrapper_7_clock = clock; // @[:@62354.4]
  assign RetimeWrapper_7_reset = reset; // @[:@62355.4]
  assign RetimeWrapper_7_io_flow = x593_inr_UnitPipe_sm_io_backpressure; // @[package.scala 95:18:@62357.4]
  assign RetimeWrapper_7_io_in = x593_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@62356.4]
  assign RetimeWrapper_8_clock = clock; // @[:@62364.4]
  assign RetimeWrapper_8_reset = reset; // @[:@62365.4]
  assign RetimeWrapper_8_io_flow = x593_inr_UnitPipe_sm_io_backpressure; // @[package.scala 95:18:@62367.4]
  assign RetimeWrapper_8_io_in = x593_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@62366.4]
  assign RetimeWrapper_9_clock = clock; // @[:@62400.4]
  assign RetimeWrapper_9_reset = reset; // @[:@62401.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@62403.4]
  assign RetimeWrapper_9_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@62402.4]
  assign RetimeWrapper_10_clock = clock; // @[:@62408.4]
  assign RetimeWrapper_10_reset = reset; // @[:@62409.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@62411.4]
  assign RetimeWrapper_10_io_in = x593_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@62410.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_clock = clock; // @[:@62437.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_reset = reset; // @[:@62438.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x555_tmp_1_rPort_0_output_0 = x555_tmp_1_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@62739.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x554_tmp_0_rPort_0_output_0 = x554_tmp_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@62762.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_in_x556_tmp_2_rPort_0_output_0 = x556_tmp_2_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@62847.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_done = x593_inr_UnitPipe_sm_io_done; // @[sm_x593_inr_UnitPipe.scala 139:22:@62872.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x593_inr_UnitPipe_sm_io_datapathEn & x593_inr_UnitPipe_mySignalsIn_mask; // @[sm_x593_inr_UnitPipe.scala 139:22:@62865.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_baseEn = _T_1029 & _T_1038; // @[sm_x593_inr_UnitPipe.scala 139:22:@62864.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_sigsIn_break = x593_inr_UnitPipe_sm_io_break; // @[sm_x593_inr_UnitPipe.scala 139:22:@62863.4]
  assign x593_inr_UnitPipe_kernelx593_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x593_inr_UnitPipe.scala 138:18:@62853.4]
  assign x594_force_0_clock = clock; // @[:@62881.4]
  assign x594_force_0_reset = reset; // @[:@62882.4]
  assign x594_force_0_io_rPort_0_en_0 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@65522.4]
  assign x594_force_0_io_wPort_0_data_0 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@64899.4]
  assign x594_force_0_io_wPort_0_en_0 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@64895.4]
  assign x594_force_0_io_sEn_0 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_sEn_0; // @[MemInterfaceType.scala 189:41:@64886.4]
  assign x594_force_0_io_sEn_1 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_sEn_1; // @[MemInterfaceType.scala 189:41:@65511.4]
  assign x594_force_0_io_sDone_0 = x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x594_force_0_sDone_0; // @[MemInterfaceType.scala 189:64:@64887.4]
  assign x594_force_0_io_sDone_1 = x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_sDone_1; // @[MemInterfaceType.scala 189:64:@65512.4]
  assign x595_reg_clock = clock; // @[:@62911.4]
  assign x595_reg_reset = reset; // @[:@62912.4]
  assign x595_reg_io_wPort_0_data_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@63591.4]
  assign x595_reg_io_wPort_0_reset = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_reset; // @[MemInterfaceType.scala 67:44:@63590.4]
  assign x595_reg_io_wPort_0_en_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@63587.4]
  assign x595_reg_io_sEn_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_sEn_0; // @[MemInterfaceType.scala 189:41:@63577.4]
  assign x595_reg_io_sEn_1 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_sEn_1; // @[MemInterfaceType.scala 189:41:@64312.4]
  assign x595_reg_io_sDone_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x595_reg_sDone_0; // @[MemInterfaceType.scala 189:64:@63578.4]
  assign x595_reg_io_sDone_1 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_sDone_1; // @[MemInterfaceType.scala 189:64:@64313.4]
  assign x596_reg_clock = clock; // @[:@62948.4]
  assign x596_reg_reset = reset; // @[:@62949.4]
  assign x596_reg_io_wPort_0_data_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@63632.4]
  assign x596_reg_io_wPort_0_reset = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_reset; // @[MemInterfaceType.scala 67:44:@63631.4]
  assign x596_reg_io_wPort_0_en_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@63628.4]
  assign x596_reg_io_sEn_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_sEn_0; // @[MemInterfaceType.scala 189:41:@63619.4]
  assign x596_reg_io_sEn_1 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x596_reg_sEn_1; // @[MemInterfaceType.scala 189:41:@64353.4]
  assign x596_reg_io_sDone_0 = x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x596_reg_sDone_0; // @[MemInterfaceType.scala 189:64:@63620.4]
  assign x596_reg_io_sDone_1 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x596_reg_sDone_1; // @[MemInterfaceType.scala 189:64:@64354.4]
  assign x605_inr_UnitPipe_sm_clock = clock; // @[:@63014.4]
  assign x605_inr_UnitPipe_sm_reset = reset; // @[:@63015.4]
  assign x605_inr_UnitPipe_sm_io_enable = _T_1136 & _T_1145; // @[SpatialBlocks.scala 139:18:@63112.4]
  assign x605_inr_UnitPipe_sm_io_ctrDone = x605_inr_UnitPipe_sm_io_ctrInc & _T_1112; // @[sm_x653_outr_Reduce.scala 138:39:@63045.4]
  assign x605_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 141:21:@63114.4]
  assign x605_inr_UnitPipe_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@63086.4]
  assign x605_inr_UnitPipe_sm_io_break = 1'h0; // @[sm_x653_outr_Reduce.scala 144:37:@63072.4]
  assign RetimeWrapper_11_clock = clock; // @[:@63047.4]
  assign RetimeWrapper_11_reset = reset; // @[:@63048.4]
  assign RetimeWrapper_11_io_flow = x605_inr_UnitPipe_sm_io_backpressure; // @[package.scala 95:18:@63050.4]
  assign RetimeWrapper_11_io_in = x605_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@63049.4]
  assign RetimeWrapper_12_clock = clock; // @[:@63057.4]
  assign RetimeWrapper_12_reset = reset; // @[:@63058.4]
  assign RetimeWrapper_12_io_flow = x605_inr_UnitPipe_sm_io_backpressure; // @[package.scala 95:18:@63060.4]
  assign RetimeWrapper_12_io_in = x605_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@63059.4]
  assign RetimeWrapper_13_clock = clock; // @[:@63093.4]
  assign RetimeWrapper_13_reset = reset; // @[:@63094.4]
  assign RetimeWrapper_13_io_flow = 1'h1; // @[package.scala 95:18:@63096.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@63095.4]
  assign RetimeWrapper_14_clock = clock; // @[:@63101.4]
  assign RetimeWrapper_14_reset = reset; // @[:@63102.4]
  assign RetimeWrapper_14_io_flow = 1'h1; // @[package.scala 95:18:@63104.4]
  assign RetimeWrapper_14_io_in = x605_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@63103.4]
  assign x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_clock = clock; // @[:@63130.4]
  assign x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_reset = reset; // @[:@63131.4]
  assign x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_in_x580_r_0_rPort_0_output_0 = x580_r_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@63564.4]
  assign x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_done = x605_inr_UnitPipe_sm_io_done; // @[sm_x605_inr_UnitPipe.scala 134:22:@63655.4]
  assign x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x605_inr_UnitPipe_sm_io_datapathEn & x605_inr_UnitPipe_mySignalsIn_mask; // @[sm_x605_inr_UnitPipe.scala 134:22:@63648.4]
  assign x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_baseEn = _T_1136 & _T_1145; // @[sm_x605_inr_UnitPipe.scala 134:22:@63647.4]
  assign x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_sigsIn_break = x605_inr_UnitPipe_sm_io_break; // @[sm_x605_inr_UnitPipe.scala 134:22:@63646.4]
  assign x605_inr_UnitPipe_kernelx605_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x605_inr_UnitPipe.scala 133:18:@63636.4]
  assign x621_inr_Switch_sm_clock = clock; // @[:@63733.4]
  assign x621_inr_Switch_sm_reset = reset; // @[:@63734.4]
  assign x621_inr_Switch_sm_io_enable = _T_1265 & _T_1274; // @[SpatialBlocks.scala 139:18:@63841.4]
  assign x621_inr_Switch_sm_io_parentAck = io_sigsIn_smChildAcks_3; // @[SpatialBlocks.scala 141:21:@63843.4]
  assign x621_inr_Switch_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@63815.4]
  assign x621_inr_Switch_sm_io_doneIn_0 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@63811.4]
  assign x621_inr_Switch_sm_io_doneIn_1 = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:72:@63812.4]
  assign x621_inr_Switch_sm_io_selectsIn_0 = x595_reg_io_rPort_0_output_0; // @[sm_x653_outr_Reduce.scala 161:46:@63767.4]
  assign x621_inr_Switch_sm_io_selectsIn_1 = x596_reg_io_rPort_0_output_0; // @[sm_x653_outr_Reduce.scala 162:46:@63768.4]
  assign RetimeWrapper_15_clock = clock; // @[:@63770.4]
  assign RetimeWrapper_15_reset = reset; // @[:@63771.4]
  assign RetimeWrapper_15_io_flow = x621_inr_Switch_sm_io_backpressure; // @[package.scala 95:18:@63773.4]
  assign RetimeWrapper_15_io_in = x621_inr_Switch_sm_io_done; // @[package.scala 94:16:@63772.4]
  assign RetimeWrapper_16_clock = clock; // @[:@63780.4]
  assign RetimeWrapper_16_reset = reset; // @[:@63781.4]
  assign RetimeWrapper_16_io_flow = x621_inr_Switch_sm_io_backpressure; // @[package.scala 95:18:@63783.4]
  assign RetimeWrapper_16_io_in = x621_inr_Switch_sm_io_done; // @[package.scala 94:16:@63782.4]
  assign RetimeWrapper_17_clock = clock; // @[:@63822.4]
  assign RetimeWrapper_17_reset = reset; // @[:@63823.4]
  assign RetimeWrapper_17_io_flow = 1'h1; // @[package.scala 95:18:@63825.4]
  assign RetimeWrapper_17_io_in = io_sigsIn_smEnableOuts_3; // @[package.scala 94:16:@63824.4]
  assign RetimeWrapper_18_clock = clock; // @[:@63830.4]
  assign RetimeWrapper_18_reset = reset; // @[:@63831.4]
  assign RetimeWrapper_18_io_flow = 1'h1; // @[package.scala 95:18:@63833.4]
  assign RetimeWrapper_18_io_in = x621_inr_Switch_sm_io_done; // @[package.scala 94:16:@63832.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_clock = clock; // @[:@63859.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_reset = reset; // @[:@63860.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x736_rd_x596 = x596_reg_io_rPort_0_output_0; // @[sm_x621_inr_Switch.scala 69:31:@64262.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x580_r_0_rPort_1_output_0 = x580_r_0_io_rPort_1_output_0; // @[MemInterfaceType.scala 66:44:@64299.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x595_reg_rPort_1_output_0 = x595_reg_io_rPort_1_output_0; // @[MemInterfaceType.scala 66:44:@64322.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_in_x735_rd_x595 = x595_reg_io_rPort_0_output_0; // @[sm_x621_inr_Switch.scala 74:31:@64345.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_done = x621_inr_Switch_sm_io_done; // @[sm_x621_inr_Switch.scala 137:22:@64384.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_baseEn = _T_1265 & _T_1274; // @[sm_x621_inr_Switch.scala 137:22:@64376.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smSelectsOut_0 = x621_inr_Switch_sm_io_selectsOut_0; // @[sm_x621_inr_Switch.scala 137:22:@64370.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smSelectsOut_1 = x621_inr_Switch_sm_io_selectsOut_1; // @[sm_x621_inr_Switch.scala 137:22:@64371.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smChildAcks_0 = x621_inr_Switch_sm_io_childAck_0; // @[sm_x621_inr_Switch.scala 137:22:@64368.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_sigsIn_smChildAcks_1 = x621_inr_Switch_sm_io_childAck_1; // @[sm_x621_inr_Switch.scala 137:22:@64369.4]
  assign x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_rr = io_rr; // @[sm_x621_inr_Switch.scala 136:18:@64362.4]
  assign x623_inr_UnitPipe_sm_clock = clock; // @[:@64432.4]
  assign x623_inr_UnitPipe_sm_reset = reset; // @[:@64433.4]
  assign x623_inr_UnitPipe_sm_io_enable = _T_1369 & _T_1378; // @[SpatialBlocks.scala 139:18:@64530.4]
  assign x623_inr_UnitPipe_sm_io_ctrDone = x623_inr_UnitPipe_sm_io_ctrInc & _T_1345; // @[sm_x653_outr_Reduce.scala 174:39:@64463.4]
  assign x623_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_4; // @[SpatialBlocks.scala 141:21:@64532.4]
  assign x623_inr_UnitPipe_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@64504.4]
  assign x623_inr_UnitPipe_sm_io_break = 1'h0; // @[sm_x653_outr_Reduce.scala 180:37:@64490.4]
  assign RetimeWrapper_19_clock = clock; // @[:@64465.4]
  assign RetimeWrapper_19_reset = reset; // @[:@64466.4]
  assign RetimeWrapper_19_io_flow = x623_inr_UnitPipe_sm_io_backpressure; // @[package.scala 95:18:@64468.4]
  assign RetimeWrapper_19_io_in = x623_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@64467.4]
  assign RetimeWrapper_20_clock = clock; // @[:@64475.4]
  assign RetimeWrapper_20_reset = reset; // @[:@64476.4]
  assign RetimeWrapper_20_io_flow = x623_inr_UnitPipe_sm_io_backpressure; // @[package.scala 95:18:@64478.4]
  assign RetimeWrapper_20_io_in = x623_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@64477.4]
  assign RetimeWrapper_21_clock = clock; // @[:@64511.4]
  assign RetimeWrapper_21_reset = reset; // @[:@64512.4]
  assign RetimeWrapper_21_io_flow = 1'h1; // @[package.scala 95:18:@64514.4]
  assign RetimeWrapper_21_io_in = io_sigsIn_smEnableOuts_4; // @[package.scala 94:16:@64513.4]
  assign RetimeWrapper_22_clock = clock; // @[:@64519.4]
  assign RetimeWrapper_22_reset = reset; // @[:@64520.4]
  assign RetimeWrapper_22_io_flow = 1'h1; // @[package.scala 95:18:@64522.4]
  assign RetimeWrapper_22_io_in = x623_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@64521.4]
  assign x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_clock = clock; // @[:@64548.4]
  assign x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_reset = reset; // @[:@64549.4]
  assign x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_in_x621_inr_Switch_number = x621_inr_Switch_kernelx621_inr_Switch_concrete1_io_ret_number; // @[sm_x623_inr_UnitPipe.scala 69:34:@64902.4]
  assign x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_done = x623_inr_UnitPipe_sm_io_done; // @[sm_x623_inr_UnitPipe.scala 107:22:@64959.4]
  assign x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x623_inr_UnitPipe_sm_io_datapathEn & x623_inr_UnitPipe_mySignalsIn_mask; // @[sm_x623_inr_UnitPipe.scala 107:22:@64952.4]
  assign x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_baseEn = _T_1369 & _T_1378; // @[sm_x623_inr_UnitPipe.scala 107:22:@64951.4]
  assign x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_sigsIn_break = x623_inr_UnitPipe_sm_io_break; // @[sm_x623_inr_UnitPipe.scala 107:22:@64950.4]
  assign x623_inr_UnitPipe_kernelx623_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x623_inr_UnitPipe.scala 106:18:@64940.4]
  assign x625_ctrchain_clock = clock; // @[:@64968.4]
  assign x625_ctrchain_reset = reset; // @[:@64969.4]
  assign x625_ctrchain_io_input_reset = x639_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@65151.4]
  assign x625_ctrchain_io_input_enable = x639_inr_Foreach_sm_io_ctrInc & x639_inr_Foreach_mySignalsIn_iiDone; // @[SpatialBlocks.scala 158:42:@65150.4]
  assign x639_inr_Foreach_sm_clock = clock; // @[:@65021.4]
  assign x639_inr_Foreach_sm_reset = reset; // @[:@65022.4]
  assign x639_inr_Foreach_sm_io_enable = _T_1475 & _T_1484; // @[SpatialBlocks.scala 139:18:@65130.4]
  assign x639_inr_Foreach_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 133:15:@65105.4]
  assign x639_inr_Foreach_sm_io_ctrDone = io_rr ? _T_1450 : 1'h0; // @[sm_x653_outr_Reduce.scala 189:38:@65057.4]
  assign x639_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_5; // @[SpatialBlocks.scala 141:21:@65132.4]
  assign x639_inr_Foreach_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@65104.4]
  assign x639_inr_Foreach_sm_io_break = 1'h0; // @[sm_x653_outr_Reduce.scala 195:36:@65084.4]
  assign x639_inr_Foreach_iiCtr_clock = clock; // @[:@65046.4]
  assign x639_inr_Foreach_iiCtr_reset = reset; // @[:@65047.4]
  assign x639_inr_Foreach_iiCtr_io_input_enable = _T_1486 & _T_1487; // @[SpatialBlocks.scala 157:27:@65139.4]
  assign x639_inr_Foreach_iiCtr_io_input_reset = x639_inr_Foreach_sm_io_rst | x639_inr_Foreach_sm_io_parentAck; // @[SpatialBlocks.scala 157:63:@65141.4]
  assign RetimeWrapper_23_clock = clock; // @[:@65050.4]
  assign RetimeWrapper_23_reset = reset; // @[:@65051.4]
  assign RetimeWrapper_23_io_flow = 1'h1; // @[package.scala 95:18:@65053.4]
  assign RetimeWrapper_23_io_in = x625_ctrchain_io_output_done; // @[package.scala 94:16:@65052.4]
  assign RetimeWrapper_24_clock = clock; // @[:@65059.4]
  assign RetimeWrapper_24_reset = reset; // @[:@65060.4]
  assign RetimeWrapper_24_io_flow = x639_inr_Foreach_sm_io_backpressure; // @[package.scala 95:18:@65062.4]
  assign RetimeWrapper_24_io_in = x639_inr_Foreach_sm_io_done; // @[package.scala 94:16:@65061.4]
  assign RetimeWrapper_25_clock = clock; // @[:@65069.4]
  assign RetimeWrapper_25_reset = reset; // @[:@65070.4]
  assign RetimeWrapper_25_io_flow = x639_inr_Foreach_sm_io_backpressure; // @[package.scala 95:18:@65072.4]
  assign RetimeWrapper_25_io_in = x639_inr_Foreach_sm_io_done; // @[package.scala 94:16:@65071.4]
  assign RetimeWrapper_26_clock = clock; // @[:@65111.4]
  assign RetimeWrapper_26_reset = reset; // @[:@65112.4]
  assign RetimeWrapper_26_io_flow = 1'h1; // @[package.scala 95:18:@65114.4]
  assign RetimeWrapper_26_io_in = io_sigsIn_smEnableOuts_5; // @[package.scala 94:16:@65113.4]
  assign RetimeWrapper_27_clock = clock; // @[:@65119.4]
  assign RetimeWrapper_27_reset = reset; // @[:@65120.4]
  assign RetimeWrapper_27_io_flow = 1'h1; // @[package.scala 95:18:@65122.4]
  assign RetimeWrapper_27_io_in = x639_inr_Foreach_sm_io_done; // @[package.scala 94:16:@65121.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_clock = clock; // @[:@65153.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_reset = reset; // @[:@65154.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_b552 = b552_chain_io_rPort_4_output_0; // @[sm_x639_inr_Foreach.scala 64:23:@65503.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x594_force_0_rPort_0_output_0 = x594_force_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@65520.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_x557_tmp_3_rPort_0_output_0 = x557_tmp_3_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@65543.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_in_b543 = io_in_b543; // @[sm_x639_inr_Foreach.scala 68:23:@65580.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_done = x639_inr_Foreach_sm_io_done; // @[sm_x639_inr_Foreach.scala 156:22:@65600.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_iiIssue = x639_inr_Foreach_iiCtr_io_output_issue | _T_1490; // @[sm_x639_inr_Foreach.scala 156:22:@65597.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_1486 & _T_1487; // @[sm_x639_inr_Foreach.scala 156:22:@65593.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_baseEn = _T_1475 & _T_1484; // @[sm_x639_inr_Foreach.scala 156:22:@65592.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_break = x639_inr_Foreach_sm_io_break; // @[sm_x639_inr_Foreach.scala 156:22:@65591.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{28{x625_ctrchain_io_output_counts_0[3]}},x625_ctrchain_io_output_counts_0}; // @[sm_x639_inr_Foreach.scala 156:22:@65586.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x625_ctrchain_io_output_oobs_0; // @[sm_x639_inr_Foreach.scala 156:22:@65585.4]
  assign x639_inr_Foreach_kernelx639_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x639_inr_Foreach.scala 155:18:@65581.4]
  assign x652_inr_Foreach_sm_clock = clock; // @[:@65645.4]
  assign x652_inr_Foreach_sm_reset = reset; // @[:@65646.4]
  assign x652_inr_Foreach_sm_io_enable = _T_1581 & _T_1590; // @[SpatialBlocks.scala 139:18:@65753.4]
  assign x652_inr_Foreach_sm_io_ctrDone = io_rr ? _T_1556 : 1'h0; // @[sm_x653_outr_Reduce.scala 200:38:@65681.4]
  assign x652_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_6; // @[SpatialBlocks.scala 141:21:@65755.4]
  assign x652_inr_Foreach_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@65727.4]
  assign x652_inr_Foreach_sm_io_break = 1'h0; // @[sm_x653_outr_Reduce.scala 206:36:@65708.4]
  assign RetimeWrapper_28_clock = clock; // @[:@65674.4]
  assign RetimeWrapper_28_reset = reset; // @[:@65675.4]
  assign RetimeWrapper_28_io_flow = 1'h1; // @[package.scala 95:18:@65677.4]
  assign RetimeWrapper_28_io_in = io_in_x549_ctrchain_output_done; // @[package.scala 94:16:@65676.4]
  assign RetimeWrapper_29_clock = clock; // @[:@65683.4]
  assign RetimeWrapper_29_reset = reset; // @[:@65684.4]
  assign RetimeWrapper_29_io_flow = x652_inr_Foreach_sm_io_backpressure; // @[package.scala 95:18:@65686.4]
  assign RetimeWrapper_29_io_in = x652_inr_Foreach_sm_io_done; // @[package.scala 94:16:@65685.4]
  assign RetimeWrapper_30_clock = clock; // @[:@65693.4]
  assign RetimeWrapper_30_reset = reset; // @[:@65694.4]
  assign RetimeWrapper_30_io_flow = x652_inr_Foreach_sm_io_backpressure; // @[package.scala 95:18:@65696.4]
  assign RetimeWrapper_30_io_in = x652_inr_Foreach_sm_io_done; // @[package.scala 94:16:@65695.4]
  assign RetimeWrapper_31_clock = clock; // @[:@65734.4]
  assign RetimeWrapper_31_reset = reset; // @[:@65735.4]
  assign RetimeWrapper_31_io_flow = 1'h1; // @[package.scala 95:18:@65737.4]
  assign RetimeWrapper_31_io_in = io_sigsIn_smEnableOuts_6; // @[package.scala 94:16:@65736.4]
  assign RetimeWrapper_32_clock = clock; // @[:@65742.4]
  assign RetimeWrapper_32_reset = reset; // @[:@65743.4]
  assign RetimeWrapper_32_io_flow = 1'h1; // @[package.scala 95:18:@65745.4]
  assign RetimeWrapper_32_io_in = x652_inr_Foreach_sm_io_done; // @[package.scala 94:16:@65744.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_clock = clock; // @[:@65776.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_reset = reset; // @[:@65777.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_b550_number = __6_io_result; // @[sm_x652_inr_Foreach.scala 57:23:@65892.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x558_tmp_4_rPort_0_output_0 = x558_tmp_4_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@65911.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_x544_accum_0_rPort_0_output_0 = io_in_x544_accum_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@65937.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_in_b543 = io_in_b543; // @[sm_x652_inr_Foreach.scala 61:23:@65949.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_done = x652_inr_Foreach_sm_io_done; // @[sm_x652_inr_Foreach.scala 128:22:@65969.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_1592 & _T_1593; // @[sm_x652_inr_Foreach.scala 128:22:@65962.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_baseEn = _T_1581 & _T_1590; // @[sm_x652_inr_Foreach.scala 128:22:@65961.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_break = x652_inr_Foreach_sm_io_break; // @[sm_x652_inr_Foreach.scala 128:22:@65960.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{28{io_in_x549_ctrchain_output_counts_0[3]}},io_in_x549_ctrchain_output_counts_0}; // @[sm_x652_inr_Foreach.scala 128:22:@65955.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = io_in_x549_ctrchain_output_oobs_0; // @[sm_x652_inr_Foreach.scala 128:22:@65954.4]
  assign x652_inr_Foreach_kernelx652_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x652_inr_Foreach.scala 127:18:@65950.4]
  assign RetimeWrapper_33_clock = clock; // @[:@65979.4]
  assign RetimeWrapper_33_reset = reset; // @[:@65980.4]
  assign RetimeWrapper_33_io_flow = 1'h1; // @[package.scala 95:18:@65982.4]
  assign RetimeWrapper_33_io_in = io_sigsIn_done; // @[package.scala 94:16:@65981.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1005 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1112 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1345 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1005 <= 1'h0;
    end else begin
      _T_1005 <= _T_1002;
    end
    if (reset) begin
      _T_1112 <= 1'h0;
    end else begin
      _T_1112 <= _T_1109;
    end
    if (reset) begin
      _T_1345 <= 1'h0;
    end else begin
      _T_1345 <= _T_1342;
    end
  end
endmodule
module x667_inr_Foreach_kernelx667_inr_Foreach_concrete1( // @[:@67547.2]
  input         clock, // @[:@67548.4]
  input         reset, // @[:@67549.4]
  input  [31:0] io_in_b542_number, // @[:@67550.4]
  output [1:0]  io_in_x545_accum_1_rPort_0_ofs_0, // @[:@67550.4]
  output        io_in_x545_accum_1_rPort_0_en_0, // @[:@67550.4]
  input  [31:0] io_in_x545_accum_1_rPort_0_output_0, // @[:@67550.4]
  output        io_in_x545_accum_1_sEn_1, // @[:@67550.4]
  output        io_in_x545_accum_1_sDone_1, // @[:@67550.4]
  output [8:0]  io_in_x473_A_sram_2_rPort_0_ofs_0, // @[:@67550.4]
  output        io_in_x473_A_sram_2_rPort_0_en_0, // @[:@67550.4]
  input  [31:0] io_in_x473_A_sram_2_rPort_0_output_0, // @[:@67550.4]
  output [8:0]  io_in_x539_out_sram_0_wPort_0_ofs_0, // @[:@67550.4]
  output [31:0] io_in_x539_out_sram_0_wPort_0_data_0, // @[:@67550.4]
  output        io_in_x539_out_sram_0_wPort_0_en_0, // @[:@67550.4]
  input         io_in_b543, // @[:@67550.4]
  input         io_sigsIn_done, // @[:@67550.4]
  input         io_sigsIn_datapathEn, // @[:@67550.4]
  input         io_sigsIn_baseEn, // @[:@67550.4]
  input         io_sigsIn_break, // @[:@67550.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@67550.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@67550.4]
  input         io_rr // @[:@67550.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@67616.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@67616.4]
  wire  x751_sum_1_clock; // @[Math.scala 150:24:@67652.4]
  wire  x751_sum_1_reset; // @[Math.scala 150:24:@67652.4]
  wire [31:0] x751_sum_1_io_a; // @[Math.scala 150:24:@67652.4]
  wire [31:0] x751_sum_1_io_b; // @[Math.scala 150:24:@67652.4]
  wire  x751_sum_1_io_flow; // @[Math.scala 150:24:@67652.4]
  wire [31:0] x751_sum_1_io_result; // @[Math.scala 150:24:@67652.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@67663.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@67663.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@67663.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@67663.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@67663.4]
  wire  x662_sum_1_clock; // @[Math.scala 150:24:@67672.4]
  wire  x662_sum_1_reset; // @[Math.scala 150:24:@67672.4]
  wire [31:0] x662_sum_1_io_a; // @[Math.scala 150:24:@67672.4]
  wire [31:0] x662_sum_1_io_b; // @[Math.scala 150:24:@67672.4]
  wire  x662_sum_1_io_flow; // @[Math.scala 150:24:@67672.4]
  wire [31:0] x662_sum_1_io_result; // @[Math.scala 150:24:@67672.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@67683.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@67683.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@67683.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@67683.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@67683.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@67693.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@67693.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@67693.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@67693.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@67693.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@67705.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@67705.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@67705.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@67705.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@67705.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@67717.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@67717.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@67717.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@67717.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@67717.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@67738.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@67738.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@67738.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@67738.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@67738.4]
  wire  x665_sum_1_clock; // @[Math.scala 150:24:@67747.4]
  wire  x665_sum_1_reset; // @[Math.scala 150:24:@67747.4]
  wire [31:0] x665_sum_1_io_a; // @[Math.scala 150:24:@67747.4]
  wire [31:0] x665_sum_1_io_b; // @[Math.scala 150:24:@67747.4]
  wire [31:0] x665_sum_1_io_result; // @[Math.scala 150:24:@67747.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@67758.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@67758.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@67758.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@67758.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@67758.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@67768.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@67768.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@67768.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@67768.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@67778.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@67778.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@67778.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@67778.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@67778.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@67792.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@67792.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@67792.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@67792.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@67792.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@67812.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@67812.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@67812.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@67812.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@67812.4]
  wire  b657; // @[sm_x667_inr_Foreach.scala 76:18:@67624.4]
  wire  _T_604; // @[sm_x667_inr_Foreach.scala 81:114:@67630.4]
  wire  _T_605; // @[sm_x667_inr_Foreach.scala 81:111:@67631.4]
  wire  _T_610; // @[implicits.scala 56:10:@67634.4]
  wire  _T_611; // @[sm_x667_inr_Foreach.scala 81:131:@67635.4]
  wire  _T_612; // @[sm_x667_inr_Foreach.scala 81:228:@67636.4]
  wire [32:0] _GEN_0; // @[Math.scala 461:32:@67648.4]
  wire [32:0] _T_618; // @[Math.scala 461:32:@67648.4]
  wire  _T_655; // @[package.scala 96:25:@67710.4 package.scala 96:25:@67711.4]
  wire  _T_657; // @[implicits.scala 56:10:@67712.4]
  wire  _T_659; // @[sm_x667_inr_Foreach.scala 102:111:@67714.4]
  wire  _T_664; // @[package.scala 96:25:@67722.4 package.scala 96:25:@67723.4]
  wire  _T_666; // @[implicits.scala 56:10:@67724.4]
  wire  _T_667; // @[sm_x667_inr_Foreach.scala 102:131:@67725.4]
  wire  x796_b657_D2; // @[package.scala 96:25:@67698.4 package.scala 96:25:@67699.4]
  wire  _T_668; // @[sm_x667_inr_Foreach.scala 102:228:@67726.4]
  wire  x795_b543_D2; // @[package.scala 96:25:@67688.4 package.scala 96:25:@67689.4]
  wire  _T_705; // @[package.scala 96:25:@67797.4 package.scala 96:25:@67798.4]
  wire  _T_707; // @[implicits.scala 56:10:@67799.4]
  wire  _T_708; // @[sm_x667_inr_Foreach.scala 121:120:@67800.4]
  wire  _T_710; // @[sm_x667_inr_Foreach.scala 121:217:@67802.4]
  wire  x800_b657_D5; // @[package.scala 96:25:@67783.4 package.scala 96:25:@67784.4]
  wire  _T_712; // @[sm_x667_inr_Foreach.scala 121:262:@67804.4]
  wire  x798_b543_D5; // @[package.scala 96:25:@67763.4 package.scala 96:25:@67764.4]
  wire  _T_717; // @[package.scala 96:25:@67817.4 package.scala 96:25:@67818.4]
  wire [31:0] b656_number; // @[Math.scala 723:22:@67621.4 Math.scala 724:14:@67622.4]
  wire [31:0] x662_sum_number; // @[Math.scala 154:22:@67678.4 Math.scala 155:14:@67679.4]
  wire [31:0] x799_x662_sum_D3_number; // @[package.scala 96:25:@67773.4 package.scala 96:25:@67774.4]
  _ _ ( // @[Math.scala 720:24:@67616.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x739_sum x751_sum_1 ( // @[Math.scala 150:24:@67652.4]
    .clock(x751_sum_1_clock),
    .reset(x751_sum_1_reset),
    .io_a(x751_sum_1_io_a),
    .io_b(x751_sum_1_io_b),
    .io_flow(x751_sum_1_io_flow),
    .io_result(x751_sum_1_io_result)
  );
  RetimeWrapper_31 RetimeWrapper ( // @[package.scala 93:22:@67663.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x739_sum x662_sum_1 ( // @[Math.scala 150:24:@67672.4]
    .clock(x662_sum_1_clock),
    .reset(x662_sum_1_reset),
    .io_a(x662_sum_1_io_a),
    .io_b(x662_sum_1_io_b),
    .io_flow(x662_sum_1_io_flow),
    .io_result(x662_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@67683.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@67693.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@67705.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@67717.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_5 ( // @[package.scala 93:22:@67738.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  x648_sum x665_sum_1 ( // @[Math.scala 150:24:@67747.4]
    .clock(x665_sum_1_clock),
    .reset(x665_sum_1_reset),
    .io_a(x665_sum_1_io_a),
    .io_b(x665_sum_1_io_b),
    .io_result(x665_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_6 ( // @[package.scala 93:22:@67758.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_705 RetimeWrapper_7 ( // @[package.scala 93:22:@67768.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_8 ( // @[package.scala 93:22:@67778.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_9 ( // @[package.scala 93:22:@67792.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@67812.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign b657 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x667_inr_Foreach.scala 76:18:@67624.4]
  assign _T_604 = ~ io_sigsIn_break; // @[sm_x667_inr_Foreach.scala 81:114:@67630.4]
  assign _T_605 = io_rr & _T_604; // @[sm_x667_inr_Foreach.scala 81:111:@67631.4]
  assign _T_610 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 56:10:@67634.4]
  assign _T_611 = _T_605 & _T_610; // @[sm_x667_inr_Foreach.scala 81:131:@67635.4]
  assign _T_612 = _T_611 & b657; // @[sm_x667_inr_Foreach.scala 81:228:@67636.4]
  assign _GEN_0 = {{1'd0}, io_in_b542_number}; // @[Math.scala 461:32:@67648.4]
  assign _T_618 = _GEN_0 << 1; // @[Math.scala 461:32:@67648.4]
  assign _T_655 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@67710.4 package.scala 96:25:@67711.4]
  assign _T_657 = io_rr ? _T_655 : 1'h0; // @[implicits.scala 56:10:@67712.4]
  assign _T_659 = _T_657 & _T_604; // @[sm_x667_inr_Foreach.scala 102:111:@67714.4]
  assign _T_664 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@67722.4 package.scala 96:25:@67723.4]
  assign _T_666 = io_rr ? _T_664 : 1'h0; // @[implicits.scala 56:10:@67724.4]
  assign _T_667 = _T_659 & _T_666; // @[sm_x667_inr_Foreach.scala 102:131:@67725.4]
  assign x796_b657_D2 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@67698.4 package.scala 96:25:@67699.4]
  assign _T_668 = _T_667 & x796_b657_D2; // @[sm_x667_inr_Foreach.scala 102:228:@67726.4]
  assign x795_b543_D2 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@67688.4 package.scala 96:25:@67689.4]
  assign _T_705 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@67797.4 package.scala 96:25:@67798.4]
  assign _T_707 = io_rr ? _T_705 : 1'h0; // @[implicits.scala 56:10:@67799.4]
  assign _T_708 = _T_604 & _T_707; // @[sm_x667_inr_Foreach.scala 121:120:@67800.4]
  assign _T_710 = _T_708 & _T_604; // @[sm_x667_inr_Foreach.scala 121:217:@67802.4]
  assign x800_b657_D5 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@67783.4 package.scala 96:25:@67784.4]
  assign _T_712 = _T_710 & x800_b657_D5; // @[sm_x667_inr_Foreach.scala 121:262:@67804.4]
  assign x798_b543_D5 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@67763.4 package.scala 96:25:@67764.4]
  assign _T_717 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@67817.4 package.scala 96:25:@67818.4]
  assign b656_number = __io_result; // @[Math.scala 723:22:@67621.4 Math.scala 724:14:@67622.4]
  assign x662_sum_number = x662_sum_1_io_result; // @[Math.scala 154:22:@67678.4 Math.scala 155:14:@67679.4]
  assign x799_x662_sum_D3_number = RetimeWrapper_7_io_out; // @[package.scala 96:25:@67773.4 package.scala 96:25:@67774.4]
  assign io_in_x545_accum_1_rPort_0_ofs_0 = b656_number[1:0]; // @[MemInterfaceType.scala 107:54:@67640.4]
  assign io_in_x545_accum_1_rPort_0_en_0 = _T_612 & io_in_b543; // @[MemInterfaceType.scala 110:79:@67642.4]
  assign io_in_x545_accum_1_sEn_1 = io_sigsIn_baseEn; // @[MemInterfaceType.scala 196:15:@67820.4]
  assign io_in_x545_accum_1_sDone_1 = io_rr ? _T_717 : 1'h0; // @[MemInterfaceType.scala 197:17:@67821.4]
  assign io_in_x473_A_sram_2_rPort_0_ofs_0 = x662_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@67730.4]
  assign io_in_x473_A_sram_2_rPort_0_en_0 = _T_668 & x795_b543_D2; // @[MemInterfaceType.scala 110:79:@67732.4]
  assign io_in_x539_out_sram_0_wPort_0_ofs_0 = x799_x662_sum_D3_number[8:0]; // @[MemInterfaceType.scala 89:54:@67807.4]
  assign io_in_x539_out_sram_0_wPort_0_data_0 = x665_sum_1_io_result; // @[MemInterfaceType.scala 90:56:@67808.4]
  assign io_in_x539_out_sram_0_wPort_0_en_0 = _T_712 & x798_b543_D5; // @[MemInterfaceType.scala 93:57:@67810.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@67619.4]
  assign x751_sum_1_clock = clock; // @[:@67653.4]
  assign x751_sum_1_reset = reset; // @[:@67654.4]
  assign x751_sum_1_io_a = _T_618[31:0]; // @[Math.scala 151:17:@67655.4]
  assign x751_sum_1_io_b = io_in_b542_number; // @[Math.scala 152:17:@67656.4]
  assign x751_sum_1_io_flow = 1'h1; // @[Math.scala 153:20:@67657.4]
  assign RetimeWrapper_clock = clock; // @[:@67664.4]
  assign RetimeWrapper_reset = reset; // @[:@67665.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@67667.4]
  assign RetimeWrapper_io_in = __io_result; // @[package.scala 94:16:@67666.4]
  assign x662_sum_1_clock = clock; // @[:@67673.4]
  assign x662_sum_1_reset = reset; // @[:@67674.4]
  assign x662_sum_1_io_a = x751_sum_1_io_result; // @[Math.scala 151:17:@67675.4]
  assign x662_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@67676.4]
  assign x662_sum_1_io_flow = 1'h1; // @[Math.scala 153:20:@67677.4]
  assign RetimeWrapper_1_clock = clock; // @[:@67684.4]
  assign RetimeWrapper_1_reset = reset; // @[:@67685.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@67687.4]
  assign RetimeWrapper_1_io_in = io_in_b543; // @[package.scala 94:16:@67686.4]
  assign RetimeWrapper_2_clock = clock; // @[:@67694.4]
  assign RetimeWrapper_2_reset = reset; // @[:@67695.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@67697.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@67696.4]
  assign RetimeWrapper_3_clock = clock; // @[:@67706.4]
  assign RetimeWrapper_3_reset = reset; // @[:@67707.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@67709.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@67708.4]
  assign RetimeWrapper_4_clock = clock; // @[:@67718.4]
  assign RetimeWrapper_4_reset = reset; // @[:@67719.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@67721.4]
  assign RetimeWrapper_4_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@67720.4]
  assign RetimeWrapper_5_clock = clock; // @[:@67739.4]
  assign RetimeWrapper_5_reset = reset; // @[:@67740.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@67742.4]
  assign RetimeWrapper_5_io_in = io_in_x545_accum_1_rPort_0_output_0; // @[package.scala 94:16:@67741.4]
  assign x665_sum_1_clock = clock; // @[:@67748.4]
  assign x665_sum_1_reset = reset; // @[:@67749.4]
  assign x665_sum_1_io_a = RetimeWrapper_5_io_out; // @[Math.scala 151:17:@67750.4]
  assign x665_sum_1_io_b = io_in_x473_A_sram_2_rPort_0_output_0; // @[Math.scala 152:17:@67751.4]
  assign RetimeWrapper_6_clock = clock; // @[:@67759.4]
  assign RetimeWrapper_6_reset = reset; // @[:@67760.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@67762.4]
  assign RetimeWrapper_6_io_in = io_in_b543; // @[package.scala 94:16:@67761.4]
  assign RetimeWrapper_7_clock = clock; // @[:@67769.4]
  assign RetimeWrapper_7_reset = reset; // @[:@67770.4]
  assign RetimeWrapper_7_io_in = x662_sum_1_io_result; // @[package.scala 94:16:@67771.4]
  assign RetimeWrapper_8_clock = clock; // @[:@67779.4]
  assign RetimeWrapper_8_reset = reset; // @[:@67780.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@67782.4]
  assign RetimeWrapper_8_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@67781.4]
  assign RetimeWrapper_9_clock = clock; // @[:@67793.4]
  assign RetimeWrapper_9_reset = reset; // @[:@67794.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@67796.4]
  assign RetimeWrapper_9_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@67795.4]
  assign RetimeWrapper_10_clock = clock; // @[:@67813.4]
  assign RetimeWrapper_10_reset = reset; // @[:@67814.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@67816.4]
  assign RetimeWrapper_10_io_in = io_sigsIn_done; // @[package.scala 94:16:@67815.4]
endmodule
module x668_outr_Foreach_kernelx668_outr_Foreach_concrete1( // @[:@67823.2]
  input         clock, // @[:@67824.4]
  input         reset, // @[:@67825.4]
  output [8:0]  io_in_x472_A_sram_1_rPort_0_ofs_0, // @[:@67826.4]
  output        io_in_x472_A_sram_1_rPort_0_en_0, // @[:@67826.4]
  input  [31:0] io_in_x472_A_sram_1_rPort_0_output_0, // @[:@67826.4]
  output [8:0]  io_in_x471_A_sram_0_rPort_0_ofs_0, // @[:@67826.4]
  output        io_in_x471_A_sram_0_rPort_0_en_0, // @[:@67826.4]
  input  [31:0] io_in_x471_A_sram_0_rPort_0_output_0, // @[:@67826.4]
  output [8:0]  io_in_x473_A_sram_2_rPort_0_ofs_0, // @[:@67826.4]
  output        io_in_x473_A_sram_2_rPort_0_en_0, // @[:@67826.4]
  input  [31:0] io_in_x473_A_sram_2_rPort_0_output_0, // @[:@67826.4]
  output [8:0]  io_in_x539_out_sram_0_wPort_0_ofs_0, // @[:@67826.4]
  output [31:0] io_in_x539_out_sram_0_wPort_0_data_0, // @[:@67826.4]
  output        io_in_x539_out_sram_0_wPort_0_en_0, // @[:@67826.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@67826.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@67826.4]
  input         io_sigsIn_smChildAcks_0, // @[:@67826.4]
  input         io_sigsIn_smChildAcks_1, // @[:@67826.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@67826.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@67826.4]
  output        io_sigsOut_smDoneIn_0, // @[:@67826.4]
  output        io_sigsOut_smDoneIn_1, // @[:@67826.4]
  output        io_sigsOut_smMaskIn_0, // @[:@67826.4]
  output        io_sigsOut_smMaskIn_1, // @[:@67826.4]
  input         io_rr // @[:@67826.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@67894.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@67894.4]
  wire  b542_chain_clock; // @[sm_x668_outr_Foreach.scala 69:30:@67902.4]
  wire  b542_chain_reset; // @[sm_x668_outr_Foreach.scala 69:30:@67902.4]
  wire [31:0] b542_chain_io_rPort_0_output_0; // @[sm_x668_outr_Foreach.scala 69:30:@67902.4]
  wire [31:0] b542_chain_io_wPort_0_data_0; // @[sm_x668_outr_Foreach.scala 69:30:@67902.4]
  wire  b542_chain_io_wPort_0_reset; // @[sm_x668_outr_Foreach.scala 69:30:@67902.4]
  wire  b542_chain_io_wPort_0_en_0; // @[sm_x668_outr_Foreach.scala 69:30:@67902.4]
  wire  b542_chain_io_sEn_0; // @[sm_x668_outr_Foreach.scala 69:30:@67902.4]
  wire  b542_chain_io_sEn_1; // @[sm_x668_outr_Foreach.scala 69:30:@67902.4]
  wire  b542_chain_io_sDone_0; // @[sm_x668_outr_Foreach.scala 69:30:@67902.4]
  wire  b542_chain_io_sDone_1; // @[sm_x668_outr_Foreach.scala 69:30:@67902.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@67931.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@67931.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@67931.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@67931.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@67931.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@67943.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@67943.4]
  wire  b543_chain_clock; // @[sm_x668_outr_Foreach.scala 73:30:@67952.4]
  wire  b543_chain_reset; // @[sm_x668_outr_Foreach.scala 73:30:@67952.4]
  wire  b543_chain_io_rPort_0_output_0; // @[sm_x668_outr_Foreach.scala 73:30:@67952.4]
  wire  b543_chain_io_wPort_0_data_0; // @[sm_x668_outr_Foreach.scala 73:30:@67952.4]
  wire  b543_chain_io_wPort_0_reset; // @[sm_x668_outr_Foreach.scala 73:30:@67952.4]
  wire  b543_chain_io_wPort_0_en_0; // @[sm_x668_outr_Foreach.scala 73:30:@67952.4]
  wire  b543_chain_io_sEn_0; // @[sm_x668_outr_Foreach.scala 73:30:@67952.4]
  wire  b543_chain_io_sEn_1; // @[sm_x668_outr_Foreach.scala 73:30:@67952.4]
  wire  b543_chain_io_sDone_0; // @[sm_x668_outr_Foreach.scala 73:30:@67952.4]
  wire  b543_chain_io_sDone_1; // @[sm_x668_outr_Foreach.scala 73:30:@67952.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@67981.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@67981.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@67981.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@67981.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@67981.4]
  wire  x544_accum_0_clock; // @[m_x544_accum_0.scala 27:22:@67991.4]
  wire  x544_accum_0_reset; // @[m_x544_accum_0.scala 27:22:@67991.4]
  wire [1:0] x544_accum_0_io_rPort_0_ofs_0; // @[m_x544_accum_0.scala 27:22:@67991.4]
  wire  x544_accum_0_io_rPort_0_en_0; // @[m_x544_accum_0.scala 27:22:@67991.4]
  wire [31:0] x544_accum_0_io_rPort_0_output_0; // @[m_x544_accum_0.scala 27:22:@67991.4]
  wire [1:0] x544_accum_0_io_wPort_0_ofs_0; // @[m_x544_accum_0.scala 27:22:@67991.4]
  wire [31:0] x544_accum_0_io_wPort_0_data_0; // @[m_x544_accum_0.scala 27:22:@67991.4]
  wire  x544_accum_0_io_wPort_0_en_0; // @[m_x544_accum_0.scala 27:22:@67991.4]
  wire  x545_accum_1_clock; // @[m_x545_accum_1.scala 27:22:@68008.4]
  wire  x545_accum_1_reset; // @[m_x545_accum_1.scala 27:22:@68008.4]
  wire [1:0] x545_accum_1_io_rPort_0_ofs_0; // @[m_x545_accum_1.scala 27:22:@68008.4]
  wire  x545_accum_1_io_rPort_0_en_0; // @[m_x545_accum_1.scala 27:22:@68008.4]
  wire [31:0] x545_accum_1_io_rPort_0_output_0; // @[m_x545_accum_1.scala 27:22:@68008.4]
  wire [1:0] x545_accum_1_io_wPort_0_ofs_0; // @[m_x545_accum_1.scala 27:22:@68008.4]
  wire [31:0] x545_accum_1_io_wPort_0_data_0; // @[m_x545_accum_1.scala 27:22:@68008.4]
  wire  x545_accum_1_io_wPort_0_en_0; // @[m_x545_accum_1.scala 27:22:@68008.4]
  wire  x545_accum_1_io_sEn_0; // @[m_x545_accum_1.scala 27:22:@68008.4]
  wire  x545_accum_1_io_sEn_1; // @[m_x545_accum_1.scala 27:22:@68008.4]
  wire  x545_accum_1_io_sDone_0; // @[m_x545_accum_1.scala 27:22:@68008.4]
  wire  x545_accum_1_io_sDone_1; // @[m_x545_accum_1.scala 27:22:@68008.4]
  wire  x547_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@68038.4]
  wire  x547_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@68038.4]
  wire  x547_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@68038.4]
  wire  x547_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@68038.4]
  wire [8:0] x547_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@68038.4]
  wire  x547_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@68038.4]
  wire  x547_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@68038.4]
  wire  x549_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@68055.4]
  wire  x549_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@68055.4]
  wire  x549_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@68055.4]
  wire  x549_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@68055.4]
  wire [3:0] x549_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@68055.4]
  wire  x549_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@68055.4]
  wire  x549_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@68055.4]
  wire  x653_outr_Reduce_sm_clock; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_reset; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_enable; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_done; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_ctrDone; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_ctrInc; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_ctrRst; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_parentAck; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_backpressure; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_doneIn_0; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_doneIn_1; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_doneIn_2; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_doneIn_3; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_doneIn_4; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_doneIn_5; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_doneIn_6; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_maskIn_0; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_maskIn_1; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_maskIn_2; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_maskIn_4; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_maskIn_5; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_enableOut_0; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_enableOut_1; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_enableOut_2; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_enableOut_3; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_enableOut_4; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_enableOut_5; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_enableOut_6; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_childAck_0; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_childAck_1; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_childAck_2; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_childAck_3; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_childAck_4; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_childAck_5; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  x653_outr_Reduce_sm_io_childAck_6; // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@68197.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@68197.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@68197.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@68197.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@68197.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@68206.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@68206.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@68206.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@68206.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@68206.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@68216.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@68216.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@68216.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@68216.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@68216.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@68287.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@68287.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@68287.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@68287.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@68287.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@68295.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@68295.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@68295.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@68295.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@68295.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_clock; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_reset; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire [8:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_en_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire [31:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_output_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire [31:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_b542_number; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire [8:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_en_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire [31:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_output_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire [1:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_ofs_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire [31:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_data_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_en_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_sEn_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_sDone_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire [1:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_ofs_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_en_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire [31:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_output_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire [1:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_ofs_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire [31:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_data_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_en_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_input_reset; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_input_enable; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire [3:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_counts_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_oobs_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_done; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_b543; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_done; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_baseEn; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_3; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_4; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_5; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_6; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_3; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_4; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_5; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_6; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire [31:0] x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_3; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_4; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_5; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_6; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_0; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_1; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_2; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_4; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_5; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_rr; // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
  wire  x655_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@68580.4]
  wire  x655_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@68580.4]
  wire  x655_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@68580.4]
  wire  x655_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@68580.4]
  wire [3:0] x655_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@68580.4]
  wire  x655_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@68580.4]
  wire  x655_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@68580.4]
  wire  x667_inr_Foreach_sm_clock; // @[sm_x667_inr_Foreach.scala 35:18:@68633.4]
  wire  x667_inr_Foreach_sm_reset; // @[sm_x667_inr_Foreach.scala 35:18:@68633.4]
  wire  x667_inr_Foreach_sm_io_enable; // @[sm_x667_inr_Foreach.scala 35:18:@68633.4]
  wire  x667_inr_Foreach_sm_io_done; // @[sm_x667_inr_Foreach.scala 35:18:@68633.4]
  wire  x667_inr_Foreach_sm_io_ctrDone; // @[sm_x667_inr_Foreach.scala 35:18:@68633.4]
  wire  x667_inr_Foreach_sm_io_datapathEn; // @[sm_x667_inr_Foreach.scala 35:18:@68633.4]
  wire  x667_inr_Foreach_sm_io_ctrInc; // @[sm_x667_inr_Foreach.scala 35:18:@68633.4]
  wire  x667_inr_Foreach_sm_io_ctrRst; // @[sm_x667_inr_Foreach.scala 35:18:@68633.4]
  wire  x667_inr_Foreach_sm_io_parentAck; // @[sm_x667_inr_Foreach.scala 35:18:@68633.4]
  wire  x667_inr_Foreach_sm_io_backpressure; // @[sm_x667_inr_Foreach.scala 35:18:@68633.4]
  wire  x667_inr_Foreach_sm_io_break; // @[sm_x667_inr_Foreach.scala 35:18:@68633.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@68662.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@68662.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@68662.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@68662.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@68662.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@68671.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@68671.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@68671.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@68671.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@68671.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@68681.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@68681.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@68681.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@68681.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@68681.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@68722.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@68722.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@68722.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@68722.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@68722.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@68730.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@68730.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@68730.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@68730.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@68730.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_clock; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_reset; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire [31:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_b542_number; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire [1:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_ofs_0; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_en_0; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire [31:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_output_0; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_sEn_1; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_sDone_1; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire [8:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_ofs_0; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_en_0; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire [31:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_output_0; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire [8:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_ofs_0; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire [31:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_data_0; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_en_0; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_b543; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_done; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_baseEn; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire [31:0] x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_rr; // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
  wire  b543_chain_read_1; // @[sm_x668_outr_Foreach.scala 75:61:@67990.4]
  wire  _T_708; // @[package.scala 96:25:@68202.4 package.scala 96:25:@68203.4]
  wire  _T_712; // @[package.scala 96:25:@68211.4 package.scala 96:25:@68212.4]
  wire  _T_716; // @[package.scala 96:25:@68221.4 package.scala 96:25:@68222.4]
  wire  _T_732; // @[package.scala 96:25:@68292.4 package.scala 96:25:@68293.4]
  wire  _T_738; // @[package.scala 96:25:@68300.4 package.scala 96:25:@68301.4]
  wire  _T_741; // @[SpatialBlocks.scala 137:99:@68303.4]
  wire  _T_815; // @[package.scala 96:25:@68667.4 package.scala 96:25:@68668.4]
  wire  _T_819; // @[package.scala 96:25:@68676.4 package.scala 96:25:@68677.4]
  wire  _T_823; // @[package.scala 96:25:@68686.4 package.scala 96:25:@68687.4]
  wire  _T_839; // @[package.scala 96:25:@68727.4 package.scala 96:25:@68728.4]
  wire  _T_845; // @[package.scala 96:25:@68735.4 package.scala 96:25:@68736.4]
  wire  _T_848; // @[SpatialBlocks.scala 137:99:@68738.4]
  wire  _T_850; // @[SpatialBlocks.scala 156:36:@68747.4]
  wire  _T_851; // @[SpatialBlocks.scala 156:78:@68748.4]
  _ _ ( // @[Math.scala 720:24:@67894.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  b542_chain b542_chain ( // @[sm_x668_outr_Foreach.scala 69:30:@67902.4]
    .clock(b542_chain_clock),
    .reset(b542_chain_reset),
    .io_rPort_0_output_0(b542_chain_io_rPort_0_output_0),
    .io_wPort_0_data_0(b542_chain_io_wPort_0_data_0),
    .io_wPort_0_reset(b542_chain_io_wPort_0_reset),
    .io_wPort_0_en_0(b542_chain_io_wPort_0_en_0),
    .io_sEn_0(b542_chain_io_sEn_0),
    .io_sEn_1(b542_chain_io_sEn_1),
    .io_sDone_0(b542_chain_io_sDone_0),
    .io_sDone_1(b542_chain_io_sDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@67931.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  _ __1 ( // @[Math.scala 720:24:@67943.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  b543_chain b543_chain ( // @[sm_x668_outr_Foreach.scala 73:30:@67952.4]
    .clock(b543_chain_clock),
    .reset(b543_chain_reset),
    .io_rPort_0_output_0(b543_chain_io_rPort_0_output_0),
    .io_wPort_0_data_0(b543_chain_io_wPort_0_data_0),
    .io_wPort_0_reset(b543_chain_io_wPort_0_reset),
    .io_wPort_0_en_0(b543_chain_io_wPort_0_en_0),
    .io_sEn_0(b543_chain_io_sEn_0),
    .io_sEn_1(b543_chain_io_sEn_1),
    .io_sDone_0(b543_chain_io_sDone_0),
    .io_sDone_1(b543_chain_io_sDone_1)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@67981.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x544_accum_0 x544_accum_0 ( // @[m_x544_accum_0.scala 27:22:@67991.4]
    .clock(x544_accum_0_clock),
    .reset(x544_accum_0_reset),
    .io_rPort_0_ofs_0(x544_accum_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x544_accum_0_io_rPort_0_en_0),
    .io_rPort_0_output_0(x544_accum_0_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(x544_accum_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x544_accum_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x544_accum_0_io_wPort_0_en_0)
  );
  x545_accum_1 x545_accum_1 ( // @[m_x545_accum_1.scala 27:22:@68008.4]
    .clock(x545_accum_1_clock),
    .reset(x545_accum_1_reset),
    .io_rPort_0_ofs_0(x545_accum_1_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x545_accum_1_io_rPort_0_en_0),
    .io_rPort_0_output_0(x545_accum_1_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(x545_accum_1_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x545_accum_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(x545_accum_1_io_wPort_0_en_0),
    .io_sEn_0(x545_accum_1_io_sEn_0),
    .io_sEn_1(x545_accum_1_io_sEn_1),
    .io_sDone_0(x545_accum_1_io_sDone_0),
    .io_sDone_1(x545_accum_1_io_sDone_1)
  );
  x478_ctrchain x547_ctrchain ( // @[SpatialBlocks.scala 37:22:@68038.4]
    .clock(x547_ctrchain_clock),
    .reset(x547_ctrchain_reset),
    .io_input_reset(x547_ctrchain_io_input_reset),
    .io_input_enable(x547_ctrchain_io_input_enable),
    .io_output_counts_0(x547_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x547_ctrchain_io_output_oobs_0),
    .io_output_done(x547_ctrchain_io_output_done)
  );
  x549_ctrchain x549_ctrchain ( // @[SpatialBlocks.scala 37:22:@68055.4]
    .clock(x549_ctrchain_clock),
    .reset(x549_ctrchain_reset),
    .io_input_reset(x549_ctrchain_io_input_reset),
    .io_input_enable(x549_ctrchain_io_input_enable),
    .io_output_counts_0(x549_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x549_ctrchain_io_output_oobs_0),
    .io_output_done(x549_ctrchain_io_output_done)
  );
  x653_outr_Reduce_sm x653_outr_Reduce_sm ( // @[sm_x653_outr_Reduce.scala 36:18:@68138.4]
    .clock(x653_outr_Reduce_sm_clock),
    .reset(x653_outr_Reduce_sm_reset),
    .io_enable(x653_outr_Reduce_sm_io_enable),
    .io_done(x653_outr_Reduce_sm_io_done),
    .io_ctrDone(x653_outr_Reduce_sm_io_ctrDone),
    .io_ctrInc(x653_outr_Reduce_sm_io_ctrInc),
    .io_ctrRst(x653_outr_Reduce_sm_io_ctrRst),
    .io_parentAck(x653_outr_Reduce_sm_io_parentAck),
    .io_backpressure(x653_outr_Reduce_sm_io_backpressure),
    .io_doneIn_0(x653_outr_Reduce_sm_io_doneIn_0),
    .io_doneIn_1(x653_outr_Reduce_sm_io_doneIn_1),
    .io_doneIn_2(x653_outr_Reduce_sm_io_doneIn_2),
    .io_doneIn_3(x653_outr_Reduce_sm_io_doneIn_3),
    .io_doneIn_4(x653_outr_Reduce_sm_io_doneIn_4),
    .io_doneIn_5(x653_outr_Reduce_sm_io_doneIn_5),
    .io_doneIn_6(x653_outr_Reduce_sm_io_doneIn_6),
    .io_maskIn_0(x653_outr_Reduce_sm_io_maskIn_0),
    .io_maskIn_1(x653_outr_Reduce_sm_io_maskIn_1),
    .io_maskIn_2(x653_outr_Reduce_sm_io_maskIn_2),
    .io_maskIn_4(x653_outr_Reduce_sm_io_maskIn_4),
    .io_maskIn_5(x653_outr_Reduce_sm_io_maskIn_5),
    .io_enableOut_0(x653_outr_Reduce_sm_io_enableOut_0),
    .io_enableOut_1(x653_outr_Reduce_sm_io_enableOut_1),
    .io_enableOut_2(x653_outr_Reduce_sm_io_enableOut_2),
    .io_enableOut_3(x653_outr_Reduce_sm_io_enableOut_3),
    .io_enableOut_4(x653_outr_Reduce_sm_io_enableOut_4),
    .io_enableOut_5(x653_outr_Reduce_sm_io_enableOut_5),
    .io_enableOut_6(x653_outr_Reduce_sm_io_enableOut_6),
    .io_childAck_0(x653_outr_Reduce_sm_io_childAck_0),
    .io_childAck_1(x653_outr_Reduce_sm_io_childAck_1),
    .io_childAck_2(x653_outr_Reduce_sm_io_childAck_2),
    .io_childAck_3(x653_outr_Reduce_sm_io_childAck_3),
    .io_childAck_4(x653_outr_Reduce_sm_io_childAck_4),
    .io_childAck_5(x653_outr_Reduce_sm_io_childAck_5),
    .io_childAck_6(x653_outr_Reduce_sm_io_childAck_6)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@68197.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@68206.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@68216.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@68287.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@68295.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x653_outr_Reduce_kernelx653_outr_Reduce_concrete1 x653_outr_Reduce_kernelx653_outr_Reduce_concrete1 ( // @[sm_x653_outr_Reduce.scala 212:24:@68329.4]
    .clock(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_clock),
    .reset(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_reset),
    .io_in_x472_A_sram_1_rPort_0_ofs_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0),
    .io_in_x472_A_sram_1_rPort_0_en_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_en_0),
    .io_in_x472_A_sram_1_rPort_0_output_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_output_0),
    .io_in_b542_number(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_b542_number),
    .io_in_x471_A_sram_0_rPort_0_ofs_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0),
    .io_in_x471_A_sram_0_rPort_0_en_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_en_0),
    .io_in_x471_A_sram_0_rPort_0_output_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_output_0),
    .io_in_x545_accum_1_wPort_0_ofs_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_ofs_0),
    .io_in_x545_accum_1_wPort_0_data_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_data_0),
    .io_in_x545_accum_1_wPort_0_en_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_en_0),
    .io_in_x545_accum_1_sEn_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_sEn_0),
    .io_in_x545_accum_1_sDone_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_sDone_0),
    .io_in_x544_accum_0_rPort_0_ofs_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_ofs_0),
    .io_in_x544_accum_0_rPort_0_en_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_en_0),
    .io_in_x544_accum_0_rPort_0_output_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_output_0),
    .io_in_x544_accum_0_wPort_0_ofs_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_ofs_0),
    .io_in_x544_accum_0_wPort_0_data_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_data_0),
    .io_in_x544_accum_0_wPort_0_en_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_en_0),
    .io_in_x549_ctrchain_input_reset(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_input_reset),
    .io_in_x549_ctrchain_input_enable(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_input_enable),
    .io_in_x549_ctrchain_output_counts_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_counts_0),
    .io_in_x549_ctrchain_output_oobs_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_oobs_0),
    .io_in_x549_ctrchain_output_done(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_done),
    .io_in_b543(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_b543),
    .io_sigsIn_done(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_done),
    .io_sigsIn_baseEn(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_smEnableOuts_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smEnableOuts_3(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_3),
    .io_sigsIn_smEnableOuts_4(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_4),
    .io_sigsIn_smEnableOuts_5(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_5),
    .io_sigsIn_smEnableOuts_6(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_6),
    .io_sigsIn_smChildAcks_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsIn_smChildAcks_3(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_3),
    .io_sigsIn_smChildAcks_4(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_4),
    .io_sigsIn_smChildAcks_5(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_5),
    .io_sigsIn_smChildAcks_6(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_6),
    .io_sigsIn_cchainOutputs_0_counts_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsOut_smDoneIn_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smDoneIn_3(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_3),
    .io_sigsOut_smDoneIn_4(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_4),
    .io_sigsOut_smDoneIn_5(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_5),
    .io_sigsOut_smDoneIn_6(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_6),
    .io_sigsOut_smMaskIn_0(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_0),
    .io_sigsOut_smMaskIn_1(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_1),
    .io_sigsOut_smMaskIn_2(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_2),
    .io_sigsOut_smMaskIn_4(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_4),
    .io_sigsOut_smMaskIn_5(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_5),
    .io_rr(x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_rr)
  );
  x549_ctrchain x655_ctrchain ( // @[SpatialBlocks.scala 37:22:@68580.4]
    .clock(x655_ctrchain_clock),
    .reset(x655_ctrchain_reset),
    .io_input_reset(x655_ctrchain_io_input_reset),
    .io_input_enable(x655_ctrchain_io_input_enable),
    .io_output_counts_0(x655_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x655_ctrchain_io_output_oobs_0),
    .io_output_done(x655_ctrchain_io_output_done)
  );
  x579_inr_Foreach_sm x667_inr_Foreach_sm ( // @[sm_x667_inr_Foreach.scala 35:18:@68633.4]
    .clock(x667_inr_Foreach_sm_clock),
    .reset(x667_inr_Foreach_sm_reset),
    .io_enable(x667_inr_Foreach_sm_io_enable),
    .io_done(x667_inr_Foreach_sm_io_done),
    .io_ctrDone(x667_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x667_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x667_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x667_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x667_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x667_inr_Foreach_sm_io_backpressure),
    .io_break(x667_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@68662.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@68671.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@68681.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@68722.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper RetimeWrapper_11 ( // @[package.scala 93:22:@68730.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  x667_inr_Foreach_kernelx667_inr_Foreach_concrete1 x667_inr_Foreach_kernelx667_inr_Foreach_concrete1 ( // @[sm_x667_inr_Foreach.scala 124:24:@68764.4]
    .clock(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_clock),
    .reset(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_reset),
    .io_in_b542_number(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_b542_number),
    .io_in_x545_accum_1_rPort_0_ofs_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_ofs_0),
    .io_in_x545_accum_1_rPort_0_en_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_en_0),
    .io_in_x545_accum_1_rPort_0_output_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_output_0),
    .io_in_x545_accum_1_sEn_1(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_sEn_1),
    .io_in_x545_accum_1_sDone_1(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_sDone_1),
    .io_in_x473_A_sram_2_rPort_0_ofs_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_ofs_0),
    .io_in_x473_A_sram_2_rPort_0_en_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_en_0),
    .io_in_x473_A_sram_2_rPort_0_output_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_output_0),
    .io_in_x539_out_sram_0_wPort_0_ofs_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_ofs_0),
    .io_in_x539_out_sram_0_wPort_0_data_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_data_0),
    .io_in_x539_out_sram_0_wPort_0_en_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_en_0),
    .io_in_b543(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_b543),
    .io_sigsIn_done(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_done),
    .io_sigsIn_datapathEn(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_baseEn(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_baseEn),
    .io_sigsIn_break(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_rr)
  );
  assign b543_chain_read_1 = b543_chain_io_rPort_0_output_0; // @[sm_x668_outr_Foreach.scala 75:61:@67990.4]
  assign _T_708 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@68202.4 package.scala 96:25:@68203.4]
  assign _T_712 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@68211.4 package.scala 96:25:@68212.4]
  assign _T_716 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@68221.4 package.scala 96:25:@68222.4]
  assign _T_732 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@68292.4 package.scala 96:25:@68293.4]
  assign _T_738 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@68300.4 package.scala 96:25:@68301.4]
  assign _T_741 = ~ _T_738; // @[SpatialBlocks.scala 137:99:@68303.4]
  assign _T_815 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@68667.4 package.scala 96:25:@68668.4]
  assign _T_819 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@68676.4 package.scala 96:25:@68677.4]
  assign _T_823 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@68686.4 package.scala 96:25:@68687.4]
  assign _T_839 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@68727.4 package.scala 96:25:@68728.4]
  assign _T_845 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@68735.4 package.scala 96:25:@68736.4]
  assign _T_848 = ~ _T_845; // @[SpatialBlocks.scala 137:99:@68738.4]
  assign _T_850 = x667_inr_Foreach_sm_io_datapathEn & b543_chain_read_1; // @[SpatialBlocks.scala 156:36:@68747.4]
  assign _T_851 = ~ x667_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 156:78:@68748.4]
  assign io_in_x472_A_sram_1_rPort_0_ofs_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@68472.4]
  assign io_in_x472_A_sram_1_rPort_0_en_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@68471.4]
  assign io_in_x471_A_sram_0_rPort_0_ofs_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@68478.4]
  assign io_in_x471_A_sram_0_rPort_0_en_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@68477.4]
  assign io_in_x473_A_sram_2_rPort_0_ofs_0 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@68874.4]
  assign io_in_x473_A_sram_2_rPort_0_en_0 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@68873.4]
  assign io_in_x539_out_sram_0_wPort_0_ofs_0 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@68881.4]
  assign io_in_x539_out_sram_0_wPort_0_data_0 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@68880.4]
  assign io_in_x539_out_sram_0_wPort_0_en_0 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@68876.4]
  assign io_sigsOut_smDoneIn_0 = x653_outr_Reduce_sm_io_done; // @[SpatialBlocks.scala 155:56:@68310.4]
  assign io_sigsOut_smDoneIn_1 = x667_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@68745.4]
  assign io_sigsOut_smMaskIn_0 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[SpatialBlocks.scala 155:86:@68311.4]
  assign io_sigsOut_smMaskIn_1 = b543_chain_io_rPort_0_output_0; // @[SpatialBlocks.scala 155:86:@68746.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@67897.4]
  assign b542_chain_clock = clock; // @[:@67903.4]
  assign b542_chain_reset = reset; // @[:@67904.4]
  assign b542_chain_io_wPort_0_data_0 = __io_result; // @[NBuffers.scala 309:54:@67929.4]
  assign b542_chain_io_wPort_0_reset = RetimeWrapper_io_out; // @[NBuffers.scala 312:23:@67938.4]
  assign b542_chain_io_wPort_0_en_0 = io_sigsOut_smDoneIn_0; // @[NBuffers.scala 311:25:@67930.4]
  assign b542_chain_io_sEn_0 = _T_732 & _T_741; // @[NBuffers.scala 302:18:@68214.4]
  assign b542_chain_io_sEn_1 = _T_839 & _T_848; // @[NBuffers.scala 302:18:@68679.4]
  assign b542_chain_io_sDone_0 = io_rr ? _T_712 : 1'h0; // @[NBuffers.scala 303:20:@68215.4]
  assign b542_chain_io_sDone_1 = io_rr ? _T_819 : 1'h0; // @[NBuffers.scala 303:20:@68680.4]
  assign RetimeWrapper_clock = clock; // @[:@67932.4]
  assign RetimeWrapper_reset = reset; // @[:@67933.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@67935.4]
  assign RetimeWrapper_io_in = b542_chain_reset; // @[package.scala 94:16:@67934.4]
  assign __1_io_b = b542_chain_io_rPort_0_output_0; // @[Math.scala 721:17:@67946.4]
  assign b543_chain_clock = clock; // @[:@67953.4]
  assign b543_chain_reset = reset; // @[:@67954.4]
  assign b543_chain_io_wPort_0_data_0 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[NBuffers.scala 308:54:@67979.4]
  assign b543_chain_io_wPort_0_reset = RetimeWrapper_1_io_out; // @[NBuffers.scala 312:23:@67988.4]
  assign b543_chain_io_wPort_0_en_0 = io_sigsOut_smDoneIn_0; // @[NBuffers.scala 311:25:@67980.4]
  assign b543_chain_io_sEn_0 = _T_732 & _T_741; // @[NBuffers.scala 302:18:@68224.4]
  assign b543_chain_io_sEn_1 = _T_839 & _T_848; // @[NBuffers.scala 302:18:@68689.4]
  assign b543_chain_io_sDone_0 = io_rr ? _T_716 : 1'h0; // @[NBuffers.scala 303:20:@68225.4]
  assign b543_chain_io_sDone_1 = io_rr ? _T_823 : 1'h0; // @[NBuffers.scala 303:20:@68690.4]
  assign RetimeWrapper_1_clock = clock; // @[:@67982.4]
  assign RetimeWrapper_1_reset = reset; // @[:@67983.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@67985.4]
  assign RetimeWrapper_1_io_in = b543_chain_reset; // @[package.scala 94:16:@67984.4]
  assign x544_accum_0_clock = clock; // @[:@67992.4]
  assign x544_accum_0_reset = reset; // @[:@67993.4]
  assign x544_accum_0_io_rPort_0_ofs_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@68506.4]
  assign x544_accum_0_io_rPort_0_en_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@68505.4]
  assign x544_accum_0_io_wPort_0_ofs_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@68513.4]
  assign x544_accum_0_io_wPort_0_data_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@68512.4]
  assign x544_accum_0_io_wPort_0_en_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@68508.4]
  assign x545_accum_1_clock = clock; // @[:@68009.4]
  assign x545_accum_1_reset = reset; // @[:@68010.4]
  assign x545_accum_1_io_rPort_0_ofs_0 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@68869.4]
  assign x545_accum_1_io_rPort_0_en_0 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@68868.4]
  assign x545_accum_1_io_wPort_0_ofs_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@68501.4]
  assign x545_accum_1_io_wPort_0_data_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@68500.4]
  assign x545_accum_1_io_wPort_0_en_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@68496.4]
  assign x545_accum_1_io_sEn_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_sEn_0; // @[MemInterfaceType.scala 189:41:@68487.4]
  assign x545_accum_1_io_sEn_1 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_sEn_1; // @[MemInterfaceType.scala 189:41:@68857.4]
  assign x545_accum_1_io_sDone_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x545_accum_1_sDone_0; // @[MemInterfaceType.scala 189:64:@68488.4]
  assign x545_accum_1_io_sDone_1 = x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_sDone_1; // @[MemInterfaceType.scala 189:64:@68858.4]
  assign x547_ctrchain_clock = clock; // @[:@68039.4]
  assign x547_ctrchain_reset = reset; // @[:@68040.4]
  assign x547_ctrchain_io_input_reset = x653_outr_Reduce_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@68328.4]
  assign x547_ctrchain_io_input_enable = x653_outr_Reduce_sm_io_ctrInc; // @[SpatialBlocks.scala 158:42:@68327.4]
  assign x549_ctrchain_clock = clock; // @[:@68056.4]
  assign x549_ctrchain_reset = reset; // @[:@68057.4]
  assign x549_ctrchain_io_input_reset = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_input_reset; // @[sm_x653_outr_Reduce.scala 67:38:@68516.4]
  assign x549_ctrchain_io_input_enable = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_input_enable; // @[sm_x653_outr_Reduce.scala 67:38:@68515.4]
  assign x653_outr_Reduce_sm_clock = clock; // @[:@68139.4]
  assign x653_outr_Reduce_sm_reset = reset; // @[:@68140.4]
  assign x653_outr_Reduce_sm_io_enable = _T_732 & _T_741; // @[SpatialBlocks.scala 139:18:@68307.4]
  assign x653_outr_Reduce_sm_io_ctrDone = io_rr ? _T_708 : 1'h0; // @[sm_x668_outr_Foreach.scala 87:38:@68205.4]
  assign x653_outr_Reduce_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@68309.4]
  assign x653_outr_Reduce_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@68281.4]
  assign x653_outr_Reduce_sm_io_doneIn_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@68267.4]
  assign x653_outr_Reduce_sm_io_doneIn_1 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:72:@68268.4]
  assign x653_outr_Reduce_sm_io_doneIn_2 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:72:@68269.4]
  assign x653_outr_Reduce_sm_io_doneIn_3 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_3; // @[SpatialBlocks.scala 130:72:@68270.4]
  assign x653_outr_Reduce_sm_io_doneIn_4 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_4; // @[SpatialBlocks.scala 130:72:@68271.4]
  assign x653_outr_Reduce_sm_io_doneIn_5 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_5; // @[SpatialBlocks.scala 130:72:@68272.4]
  assign x653_outr_Reduce_sm_io_doneIn_6 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smDoneIn_6; // @[SpatialBlocks.scala 130:72:@68273.4]
  assign x653_outr_Reduce_sm_io_maskIn_0 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_0; // @[SpatialBlocks.scala 131:72:@68274.4]
  assign x653_outr_Reduce_sm_io_maskIn_1 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_1; // @[SpatialBlocks.scala 131:72:@68275.4]
  assign x653_outr_Reduce_sm_io_maskIn_2 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_2; // @[SpatialBlocks.scala 131:72:@68276.4]
  assign x653_outr_Reduce_sm_io_maskIn_4 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_4; // @[SpatialBlocks.scala 131:72:@68278.4]
  assign x653_outr_Reduce_sm_io_maskIn_5 = x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsOut_smMaskIn_5; // @[SpatialBlocks.scala 131:72:@68279.4]
  assign RetimeWrapper_2_clock = clock; // @[:@68198.4]
  assign RetimeWrapper_2_reset = reset; // @[:@68199.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@68201.4]
  assign RetimeWrapper_2_io_in = x547_ctrchain_io_output_done; // @[package.scala 94:16:@68200.4]
  assign RetimeWrapper_3_clock = clock; // @[:@68207.4]
  assign RetimeWrapper_3_reset = reset; // @[:@68208.4]
  assign RetimeWrapper_3_io_flow = x653_outr_Reduce_sm_io_backpressure; // @[package.scala 95:18:@68210.4]
  assign RetimeWrapper_3_io_in = x653_outr_Reduce_sm_io_done; // @[package.scala 94:16:@68209.4]
  assign RetimeWrapper_4_clock = clock; // @[:@68217.4]
  assign RetimeWrapper_4_reset = reset; // @[:@68218.4]
  assign RetimeWrapper_4_io_flow = x653_outr_Reduce_sm_io_backpressure; // @[package.scala 95:18:@68220.4]
  assign RetimeWrapper_4_io_in = x653_outr_Reduce_sm_io_done; // @[package.scala 94:16:@68219.4]
  assign RetimeWrapper_5_clock = clock; // @[:@68288.4]
  assign RetimeWrapper_5_reset = reset; // @[:@68289.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@68291.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@68290.4]
  assign RetimeWrapper_6_clock = clock; // @[:@68296.4]
  assign RetimeWrapper_6_reset = reset; // @[:@68297.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@68299.4]
  assign RetimeWrapper_6_io_in = x653_outr_Reduce_sm_io_done; // @[package.scala 94:16:@68298.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_clock = clock; // @[:@68330.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_reset = reset; // @[:@68331.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x472_A_sram_1_rPort_0_output_0 = io_in_x472_A_sram_1_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@68469.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_b542_number = __io_result; // @[sm_x653_outr_Reduce.scala 63:23:@68474.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x471_A_sram_0_rPort_0_output_0 = io_in_x471_A_sram_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@68475.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x544_accum_0_rPort_0_output_0 = x544_accum_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@68503.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_counts_0 = x549_ctrchain_io_output_counts_0; // @[sm_x653_outr_Reduce.scala 67:96:@68521.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_oobs_0 = x549_ctrchain_io_output_oobs_0; // @[sm_x653_outr_Reduce.scala 67:96:@68520.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_x549_ctrchain_output_done = x549_ctrchain_io_output_done; // @[sm_x653_outr_Reduce.scala 67:96:@68518.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_in_b543 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x653_outr_Reduce.scala 68:23:@68522.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_done = x653_outr_Reduce_sm_io_done; // @[sm_x653_outr_Reduce.scala 217:22:@68560.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_baseEn = _T_732 & _T_741; // @[sm_x653_outr_Reduce.scala 217:22:@68552.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_0 = x653_outr_Reduce_sm_io_enableOut_0; // @[sm_x653_outr_Reduce.scala 217:22:@68543.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_1 = x653_outr_Reduce_sm_io_enableOut_1; // @[sm_x653_outr_Reduce.scala 217:22:@68544.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_2 = x653_outr_Reduce_sm_io_enableOut_2; // @[sm_x653_outr_Reduce.scala 217:22:@68545.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_3 = x653_outr_Reduce_sm_io_enableOut_3; // @[sm_x653_outr_Reduce.scala 217:22:@68546.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_4 = x653_outr_Reduce_sm_io_enableOut_4; // @[sm_x653_outr_Reduce.scala 217:22:@68547.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_5 = x653_outr_Reduce_sm_io_enableOut_5; // @[sm_x653_outr_Reduce.scala 217:22:@68548.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smEnableOuts_6 = x653_outr_Reduce_sm_io_enableOut_6; // @[sm_x653_outr_Reduce.scala 217:22:@68549.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_0 = x653_outr_Reduce_sm_io_childAck_0; // @[sm_x653_outr_Reduce.scala 217:22:@68529.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_1 = x653_outr_Reduce_sm_io_childAck_1; // @[sm_x653_outr_Reduce.scala 217:22:@68530.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_2 = x653_outr_Reduce_sm_io_childAck_2; // @[sm_x653_outr_Reduce.scala 217:22:@68531.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_3 = x653_outr_Reduce_sm_io_childAck_3; // @[sm_x653_outr_Reduce.scala 217:22:@68532.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_4 = x653_outr_Reduce_sm_io_childAck_4; // @[sm_x653_outr_Reduce.scala 217:22:@68533.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_5 = x653_outr_Reduce_sm_io_childAck_5; // @[sm_x653_outr_Reduce.scala 217:22:@68534.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_smChildAcks_6 = x653_outr_Reduce_sm_io_childAck_6; // @[sm_x653_outr_Reduce.scala 217:22:@68535.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{23{x547_ctrchain_io_output_counts_0[8]}},x547_ctrchain_io_output_counts_0}; // @[sm_x653_outr_Reduce.scala 217:22:@68528.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x547_ctrchain_io_output_oobs_0; // @[sm_x653_outr_Reduce.scala 217:22:@68527.4]
  assign x653_outr_Reduce_kernelx653_outr_Reduce_concrete1_io_rr = io_rr; // @[sm_x653_outr_Reduce.scala 216:18:@68523.4]
  assign x655_ctrchain_clock = clock; // @[:@68581.4]
  assign x655_ctrchain_reset = reset; // @[:@68582.4]
  assign x655_ctrchain_io_input_reset = x667_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@68763.4]
  assign x655_ctrchain_io_input_enable = x667_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 158:42:@68762.4]
  assign x667_inr_Foreach_sm_clock = clock; // @[:@68634.4]
  assign x667_inr_Foreach_sm_reset = reset; // @[:@68635.4]
  assign x667_inr_Foreach_sm_io_enable = _T_839 & _T_848; // @[SpatialBlocks.scala 139:18:@68742.4]
  assign x667_inr_Foreach_sm_io_ctrDone = io_rr ? _T_815 : 1'h0; // @[sm_x668_outr_Foreach.scala 102:38:@68670.4]
  assign x667_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 141:21:@68744.4]
  assign x667_inr_Foreach_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@68716.4]
  assign x667_inr_Foreach_sm_io_break = 1'h0; // @[sm_x668_outr_Foreach.scala 108:36:@68697.4]
  assign RetimeWrapper_7_clock = clock; // @[:@68663.4]
  assign RetimeWrapper_7_reset = reset; // @[:@68664.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@68666.4]
  assign RetimeWrapper_7_io_in = x655_ctrchain_io_output_done; // @[package.scala 94:16:@68665.4]
  assign RetimeWrapper_8_clock = clock; // @[:@68672.4]
  assign RetimeWrapper_8_reset = reset; // @[:@68673.4]
  assign RetimeWrapper_8_io_flow = x667_inr_Foreach_sm_io_backpressure; // @[package.scala 95:18:@68675.4]
  assign RetimeWrapper_8_io_in = x667_inr_Foreach_sm_io_done; // @[package.scala 94:16:@68674.4]
  assign RetimeWrapper_9_clock = clock; // @[:@68682.4]
  assign RetimeWrapper_9_reset = reset; // @[:@68683.4]
  assign RetimeWrapper_9_io_flow = x667_inr_Foreach_sm_io_backpressure; // @[package.scala 95:18:@68685.4]
  assign RetimeWrapper_9_io_in = x667_inr_Foreach_sm_io_done; // @[package.scala 94:16:@68684.4]
  assign RetimeWrapper_10_clock = clock; // @[:@68723.4]
  assign RetimeWrapper_10_reset = reset; // @[:@68724.4]
  assign RetimeWrapper_10_io_flow = 1'h1; // @[package.scala 95:18:@68726.4]
  assign RetimeWrapper_10_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@68725.4]
  assign RetimeWrapper_11_clock = clock; // @[:@68731.4]
  assign RetimeWrapper_11_reset = reset; // @[:@68732.4]
  assign RetimeWrapper_11_io_flow = 1'h1; // @[package.scala 95:18:@68734.4]
  assign RetimeWrapper_11_io_in = x667_inr_Foreach_sm_io_done; // @[package.scala 94:16:@68733.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_clock = clock; // @[:@68765.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_reset = reset; // @[:@68766.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_b542_number = __1_io_result; // @[sm_x667_inr_Foreach.scala 57:23:@68849.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x545_accum_1_rPort_0_output_0 = x545_accum_1_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@68866.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_output_0 = io_in_x473_A_sram_2_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@68871.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_in_b543 = b543_chain_io_rPort_0_output_0; // @[sm_x667_inr_Foreach.scala 61:23:@68883.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_done = x667_inr_Foreach_sm_io_done; // @[sm_x667_inr_Foreach.scala 129:22:@68903.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_850 & _T_851; // @[sm_x667_inr_Foreach.scala 129:22:@68896.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_baseEn = _T_839 & _T_848; // @[sm_x667_inr_Foreach.scala 129:22:@68895.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_break = x667_inr_Foreach_sm_io_break; // @[sm_x667_inr_Foreach.scala 129:22:@68894.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{28{x655_ctrchain_io_output_counts_0[3]}},x655_ctrchain_io_output_counts_0}; // @[sm_x667_inr_Foreach.scala 129:22:@68889.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x655_ctrchain_io_output_oobs_0; // @[sm_x667_inr_Foreach.scala 129:22:@68888.4]
  assign x667_inr_Foreach_kernelx667_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x667_inr_Foreach.scala 128:18:@68884.4]
endmodule
module x724_outr_UnitPipe_DenseTransfer_sm( // @[:@69111.2]
  input   clock, // @[:@69112.4]
  input   reset, // @[:@69113.4]
  input   io_enable, // @[:@69114.4]
  output  io_done, // @[:@69114.4]
  input   io_parentAck, // @[:@69114.4]
  input   io_doneIn_0, // @[:@69114.4]
  output  io_enableOut_0, // @[:@69114.4]
  output  io_childAck_0, // @[:@69114.4]
  input   io_ctrCopyDone_0 // @[:@69114.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@69117.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@69117.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@69117.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@69117.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@69117.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@69117.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@69120.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@69120.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@69120.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@69120.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@69120.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@69120.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@69137.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@69137.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@69137.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@69137.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@69137.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@69137.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@69168.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@69168.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@69168.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@69168.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@69168.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@69182.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@69182.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@69182.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@69182.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@69182.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@69200.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@69200.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@69200.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@69200.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@69200.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@69237.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@69237.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@69237.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@69237.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@69237.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@69254.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@69254.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@69254.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@69254.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@69254.4]
  wire  _T_105; // @[Controllers.scala 165:35:@69152.4]
  wire  _T_107; // @[Controllers.scala 165:60:@69153.4]
  wire  _T_108; // @[Controllers.scala 165:58:@69154.4]
  wire  _T_110; // @[Controllers.scala 165:76:@69155.4]
  wire  _T_111; // @[Controllers.scala 165:74:@69156.4]
  wire  _T_115; // @[Controllers.scala 165:109:@69159.4]
  wire  _T_118; // @[Controllers.scala 165:141:@69161.4]
  wire  _T_126; // @[package.scala 96:25:@69173.4 package.scala 96:25:@69174.4]
  wire  _T_130; // @[Controllers.scala 167:54:@69176.4]
  wire  _T_131; // @[Controllers.scala 167:52:@69177.4]
  wire  _T_138; // @[package.scala 96:25:@69187.4 package.scala 96:25:@69188.4]
  wire  _T_156; // @[package.scala 96:25:@69205.4 package.scala 96:25:@69206.4]
  wire  _T_160; // @[Controllers.scala 169:67:@69208.4]
  wire  _T_161; // @[Controllers.scala 169:86:@69209.4]
  wire  _T_174; // @[Controllers.scala 213:68:@69223.4]
  wire  _T_176; // @[Controllers.scala 213:90:@69225.4]
  wire  _T_178; // @[Controllers.scala 213:132:@69227.4]
  reg  _T_186; // @[package.scala 48:56:@69233.4]
  reg [31:0] _RAND_0;
  wire  _T_187; // @[package.scala 100:41:@69235.4]
  reg  _T_200; // @[package.scala 48:56:@69251.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@69117.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@69120.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@69137.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@69168.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@69182.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@69200.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@69237.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@69254.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_105 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@69152.4]
  assign _T_107 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@69153.4]
  assign _T_108 = _T_105 & _T_107; // @[Controllers.scala 165:58:@69154.4]
  assign _T_110 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@69155.4]
  assign _T_111 = _T_108 & _T_110; // @[Controllers.scala 165:74:@69156.4]
  assign _T_115 = _T_111 & io_enable; // @[Controllers.scala 165:109:@69159.4]
  assign _T_118 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@69161.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@69173.4 package.scala 96:25:@69174.4]
  assign _T_130 = _T_126 == 1'h0; // @[Controllers.scala 167:54:@69176.4]
  assign _T_131 = io_doneIn_0 | _T_130; // @[Controllers.scala 167:52:@69177.4]
  assign _T_138 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@69187.4 package.scala 96:25:@69188.4]
  assign _T_156 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@69205.4 package.scala 96:25:@69206.4]
  assign _T_160 = _T_156 == 1'h0; // @[Controllers.scala 169:67:@69208.4]
  assign _T_161 = _T_160 & io_enable; // @[Controllers.scala 169:86:@69209.4]
  assign _T_174 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@69223.4]
  assign _T_176 = _T_174 & _T_105; // @[Controllers.scala 213:90:@69225.4]
  assign _T_178 = ~ done_0_io_output; // @[Controllers.scala 213:132:@69227.4]
  assign _T_187 = done_0_io_output & _T_186; // @[package.scala 100:41:@69235.4]
  assign io_done = RetimeWrapper_4_io_out; // @[Controllers.scala 245:13:@69261.4]
  assign io_enableOut_0 = _T_176 & _T_178; // @[Controllers.scala 213:55:@69231.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@69222.4]
  assign active_0_clock = clock; // @[:@69118.4]
  assign active_0_reset = reset; // @[:@69119.4]
  assign active_0_io_input_set = _T_115 & _T_118; // @[Controllers.scala 165:32:@69163.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@69167.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@69125.4]
  assign done_0_clock = clock; // @[:@69121.4]
  assign done_0_reset = reset; // @[:@69122.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_161; // @[Controllers.scala 169:30:@69213.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@69135.4 Controllers.scala 170:32:@69220.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@69126.4]
  assign iterDone_0_clock = clock; // @[:@69138.4]
  assign iterDone_0_reset = reset; // @[:@69139.4]
  assign iterDone_0_io_input_set = _T_131 & io_enable; // @[Controllers.scala 167:34:@69181.4]
  assign iterDone_0_io_input_reset = _T_138 | io_parentAck; // @[Controllers.scala 92:37:@69149.4 Controllers.scala 168:36:@69197.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@69140.4]
  assign RetimeWrapper_clock = clock; // @[:@69169.4]
  assign RetimeWrapper_reset = reset; // @[:@69170.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@69172.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@69171.4]
  assign RetimeWrapper_1_clock = clock; // @[:@69183.4]
  assign RetimeWrapper_1_reset = reset; // @[:@69184.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@69186.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@69185.4]
  assign RetimeWrapper_2_clock = clock; // @[:@69201.4]
  assign RetimeWrapper_2_reset = reset; // @[:@69202.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@69204.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@69203.4]
  assign RetimeWrapper_3_clock = clock; // @[:@69238.4]
  assign RetimeWrapper_3_reset = reset; // @[:@69239.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@69241.4]
  assign RetimeWrapper_3_io_in = _T_187 | io_parentAck; // @[package.scala 94:16:@69240.4]
  assign RetimeWrapper_4_clock = clock; // @[:@69255.4]
  assign RetimeWrapper_4_reset = reset; // @[:@69256.4]
  assign RetimeWrapper_4_io_flow = io_enable; // @[package.scala 95:18:@69258.4]
  assign RetimeWrapper_4_io_in = done_0_io_output & _T_200; // @[package.scala 94:16:@69257.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_200 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= _T_110;
    end
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_110;
    end
  end
endmodule
module x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1( // @[:@72154.2]
  input         clock, // @[:@72155.4]
  input         reset, // @[:@72156.4]
  output [31:0] io_in_x677_reg_wPort_0_data_0, // @[:@72157.4]
  output        io_in_x677_reg_wPort_0_reset, // @[:@72157.4]
  output        io_in_x677_reg_wPort_0_en_0, // @[:@72157.4]
  output        io_in_x677_reg_reset, // @[:@72157.4]
  output [31:0] io_in_x678_reg_wPort_0_data_0, // @[:@72157.4]
  output        io_in_x678_reg_wPort_0_reset, // @[:@72157.4]
  output        io_in_x678_reg_wPort_0_en_0, // @[:@72157.4]
  output        io_in_x678_reg_reset, // @[:@72157.4]
  input         io_in_x669_ready, // @[:@72157.4]
  output        io_in_x669_valid, // @[:@72157.4]
  output [63:0] io_in_x669_bits_addr, // @[:@72157.4]
  output [31:0] io_in_x669_bits_size, // @[:@72157.4]
  input  [31:0] io_in_b674_number, // @[:@72157.4]
  input  [63:0] io_in_x470_out_host_number, // @[:@72157.4]
  output [31:0] io_in_x676_reg_wPort_0_data_0, // @[:@72157.4]
  output        io_in_x676_reg_wPort_0_reset, // @[:@72157.4]
  output        io_in_x676_reg_wPort_0_en_0, // @[:@72157.4]
  output        io_in_x676_reg_reset, // @[:@72157.4]
  input         io_sigsIn_backpressure, // @[:@72157.4]
  input         io_sigsIn_datapathEn, // @[:@72157.4]
  input         io_sigsIn_break, // @[:@72157.4]
  input         io_rr // @[:@72157.4]
);
  wire  x753_sum_1_clock; // @[Math.scala 150:24:@72214.4]
  wire  x753_sum_1_reset; // @[Math.scala 150:24:@72214.4]
  wire [31:0] x753_sum_1_io_a; // @[Math.scala 150:24:@72214.4]
  wire [31:0] x753_sum_1_io_b; // @[Math.scala 150:24:@72214.4]
  wire  x753_sum_1_io_flow; // @[Math.scala 150:24:@72214.4]
  wire [31:0] x753_sum_1_io_result; // @[Math.scala 150:24:@72214.4]
  wire  x683_sub_1_clock; // @[Math.scala 191:24:@72251.4]
  wire  x683_sub_1_reset; // @[Math.scala 191:24:@72251.4]
  wire [31:0] x683_sub_1_io_a; // @[Math.scala 191:24:@72251.4]
  wire [31:0] x683_sub_1_io_b; // @[Math.scala 191:24:@72251.4]
  wire  x683_sub_1_io_flow; // @[Math.scala 191:24:@72251.4]
  wire [31:0] x683_sub_1_io_result; // @[Math.scala 191:24:@72251.4]
  wire  x684_sum_1_clock; // @[Math.scala 150:24:@72263.4]
  wire  x684_sum_1_reset; // @[Math.scala 150:24:@72263.4]
  wire [31:0] x684_sum_1_io_a; // @[Math.scala 150:24:@72263.4]
  wire [31:0] x684_sum_1_io_b; // @[Math.scala 150:24:@72263.4]
  wire  x684_sum_1_io_flow; // @[Math.scala 150:24:@72263.4]
  wire [31:0] x684_sum_1_io_result; // @[Math.scala 150:24:@72263.4]
  wire  x685_sum_1_clock; // @[Math.scala 150:24:@72275.4]
  wire  x685_sum_1_reset; // @[Math.scala 150:24:@72275.4]
  wire [31:0] x685_sum_1_io_a; // @[Math.scala 150:24:@72275.4]
  wire [31:0] x685_sum_1_io_b; // @[Math.scala 150:24:@72275.4]
  wire  x685_sum_1_io_flow; // @[Math.scala 150:24:@72275.4]
  wire [31:0] x685_sum_1_io_result; // @[Math.scala 150:24:@72275.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@72304.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@72304.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@72304.4]
  wire [35:0] RetimeWrapper_io_in; // @[package.scala 93:22:@72304.4]
  wire [35:0] RetimeWrapper_io_out; // @[package.scala 93:22:@72304.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@72316.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@72316.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@72316.4]
  wire [37:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@72316.4]
  wire [37:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@72316.4]
  wire [31:0] x689_1_io_b; // @[Math.scala 720:24:@72326.4]
  wire [63:0] x689_1_io_result; // @[Math.scala 720:24:@72326.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@72336.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@72336.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@72336.4]
  wire [63:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@72336.4]
  wire [63:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@72336.4]
  wire  x691_sum_1_clock; // @[Math.scala 150:24:@72345.4]
  wire  x691_sum_1_reset; // @[Math.scala 150:24:@72345.4]
  wire [63:0] x691_sum_1_io_a; // @[Math.scala 150:24:@72345.4]
  wire [63:0] x691_sum_1_io_b; // @[Math.scala 150:24:@72345.4]
  wire  x691_sum_1_io_flow; // @[Math.scala 150:24:@72345.4]
  wire [63:0] x691_sum_1_io_result; // @[Math.scala 150:24:@72345.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@72356.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@72356.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@72356.4]
  wire [63:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@72356.4]
  wire [63:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@72356.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@72370.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@72370.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@72370.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@72370.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@72370.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@72380.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@72380.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@72380.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@72380.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@72380.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@72399.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@72399.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@72399.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@72399.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@72399.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@72419.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@72419.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@72419.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@72419.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@72419.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@72439.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@72439.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@72439.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@72439.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@72439.4]
  wire [32:0] _GEN_0; // @[Math.scala 461:32:@72210.4]
  wire [32:0] _T_508; // @[Math.scala 461:32:@72210.4]
  wire [31:0] x753_sum_number; // @[Math.scala 154:22:@72220.4 Math.scala 155:14:@72221.4]
  wire  _T_514; // @[FixedPoint.scala 50:25:@72225.4]
  wire [3:0] _T_518; // @[Bitwise.scala 72:12:@72227.4]
  wire [27:0] _T_519; // @[FixedPoint.scala 18:52:@72228.4]
  wire  _T_525; // @[Math.scala 451:55:@72230.4]
  wire [3:0] _T_526; // @[FixedPoint.scala 18:52:@72231.4]
  wire  _T_532; // @[Math.scala 451:110:@72233.4]
  wire  _T_533; // @[Math.scala 451:94:@72234.4]
  wire [31:0] _T_535; // @[Cat.scala 30:58:@72236.4]
  wire [31:0] x680_1_number; // @[Math.scala 454:20:@72237.4]
  wire [35:0] _GEN_1; // @[Math.scala 461:32:@72242.4]
  wire [35:0] _T_540; // @[Math.scala 461:32:@72242.4]
  wire [37:0] _GEN_2; // @[Math.scala 461:32:@72247.4]
  wire [37:0] _T_543; // @[Math.scala 461:32:@72247.4]
  wire [31:0] x685_sum_number; // @[Math.scala 154:22:@72281.4 Math.scala 155:14:@72282.4]
  wire  _T_563; // @[FixedPoint.scala 50:25:@72286.4]
  wire [3:0] _T_567; // @[Bitwise.scala 72:12:@72288.4]
  wire [27:0] _T_568; // @[FixedPoint.scala 18:52:@72289.4]
  wire  _T_574; // @[Math.scala 451:55:@72291.4]
  wire [3:0] _T_575; // @[FixedPoint.scala 18:52:@72292.4]
  wire  _T_581; // @[Math.scala 451:110:@72294.4]
  wire  _T_582; // @[Math.scala 451:94:@72295.4]
  wire [31:0] _T_584; // @[Cat.scala 30:58:@72297.4]
  wire [31:0] x686_1_number; // @[Math.scala 454:20:@72298.4]
  wire [35:0] _GEN_3; // @[Math.scala 461:32:@72303.4]
  wire [37:0] _GEN_4; // @[Math.scala 461:32:@72315.4]
  wire [37:0] _T_596; // @[package.scala 96:25:@72321.4 package.scala 96:25:@72322.4]
  wire [31:0] x755_1_number; // @[Math.scala 459:22:@72314.4 Math.scala 461:14:@72323.4]
  wire [63:0] x802_x691_sum_D1_number; // @[package.scala 96:25:@72361.4 package.scala 96:25:@72362.4]
  wire [96:0] x692_tuple; // @[Cat.scala 30:58:@72366.4]
  wire  _T_626; // @[package.scala 96:25:@72385.4 package.scala 96:25:@72386.4]
  wire  _T_628; // @[implicits.scala 56:10:@72387.4]
  wire  x803_x693_D4; // @[package.scala 96:25:@72375.4 package.scala 96:25:@72376.4]
  wire  _T_629; // @[sm_x698_inr_UnitPipe.scala 116:121:@72388.4]
  wire  _T_633; // @[sm_x698_inr_UnitPipe.scala 123:116:@72395.4]
  wire  _T_639; // @[package.scala 96:25:@72404.4 package.scala 96:25:@72405.4]
  wire  _T_641; // @[implicits.scala 56:10:@72406.4]
  wire  _T_642; // @[sm_x698_inr_UnitPipe.scala 123:133:@72407.4]
  wire  _T_644; // @[sm_x698_inr_UnitPipe.scala 123:230:@72409.4]
  wire  _T_654; // @[package.scala 96:25:@72424.4 package.scala 96:25:@72425.4]
  wire  _T_656; // @[implicits.scala 56:10:@72426.4]
  wire  _T_657; // @[sm_x698_inr_UnitPipe.scala 128:133:@72427.4]
  wire  _T_659; // @[sm_x698_inr_UnitPipe.scala 128:230:@72429.4]
  wire  _T_669; // @[package.scala 96:25:@72444.4 package.scala 96:25:@72445.4]
  wire  _T_671; // @[implicits.scala 56:10:@72446.4]
  wire  _T_672; // @[sm_x698_inr_UnitPipe.scala 133:133:@72447.4]
  wire  _T_674; // @[sm_x698_inr_UnitPipe.scala 133:230:@72449.4]
  wire [35:0] _T_591; // @[package.scala 96:25:@72309.4 package.scala 96:25:@72310.4]
  x739_sum x753_sum_1 ( // @[Math.scala 150:24:@72214.4]
    .clock(x753_sum_1_clock),
    .reset(x753_sum_1_reset),
    .io_a(x753_sum_1_io_a),
    .io_b(x753_sum_1_io_b),
    .io_flow(x753_sum_1_io_flow),
    .io_result(x753_sum_1_io_result)
  );
  x485_sub x683_sub_1 ( // @[Math.scala 191:24:@72251.4]
    .clock(x683_sub_1_clock),
    .reset(x683_sub_1_reset),
    .io_a(x683_sub_1_io_a),
    .io_b(x683_sub_1_io_b),
    .io_flow(x683_sub_1_io_flow),
    .io_result(x683_sub_1_io_result)
  );
  x739_sum x684_sum_1 ( // @[Math.scala 150:24:@72263.4]
    .clock(x684_sum_1_clock),
    .reset(x684_sum_1_reset),
    .io_a(x684_sum_1_io_a),
    .io_b(x684_sum_1_io_b),
    .io_flow(x684_sum_1_io_flow),
    .io_result(x684_sum_1_io_result)
  );
  x739_sum x685_sum_1 ( // @[Math.scala 150:24:@72275.4]
    .clock(x685_sum_1_clock),
    .reset(x685_sum_1_reset),
    .io_a(x685_sum_1_io_a),
    .io_b(x685_sum_1_io_b),
    .io_flow(x685_sum_1_io_flow),
    .io_result(x685_sum_1_io_result)
  );
  RetimeWrapper_35 RetimeWrapper ( // @[package.scala 93:22:@72304.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_36 RetimeWrapper_1 ( // @[package.scala 93:22:@72316.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x491 x689_1 ( // @[Math.scala 720:24:@72326.4]
    .io_b(x689_1_io_b),
    .io_result(x689_1_io_result)
  );
  RetimeWrapper_37 RetimeWrapper_2 ( // @[package.scala 93:22:@72336.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x493_sum x691_sum_1 ( // @[Math.scala 150:24:@72345.4]
    .clock(x691_sum_1_clock),
    .reset(x691_sum_1_reset),
    .io_a(x691_sum_1_io_a),
    .io_b(x691_sum_1_io_b),
    .io_flow(x691_sum_1_io_flow),
    .io_result(x691_sum_1_io_result)
  );
  RetimeWrapper_37 RetimeWrapper_3 ( // @[package.scala 93:22:@72356.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@72370.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_5 ( // @[package.scala 93:22:@72380.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@72399.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_58 RetimeWrapper_7 ( // @[package.scala 93:22:@72419.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_8 ( // @[package.scala 93:22:@72439.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  assign _GEN_0 = {{1'd0}, io_in_b674_number}; // @[Math.scala 461:32:@72210.4]
  assign _T_508 = _GEN_0 << 1; // @[Math.scala 461:32:@72210.4]
  assign x753_sum_number = x753_sum_1_io_result; // @[Math.scala 154:22:@72220.4 Math.scala 155:14:@72221.4]
  assign _T_514 = x753_sum_number[31]; // @[FixedPoint.scala 50:25:@72225.4]
  assign _T_518 = _T_514 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@72227.4]
  assign _T_519 = x753_sum_number[31:4]; // @[FixedPoint.scala 18:52:@72228.4]
  assign _T_525 = _T_519 == 28'hfffffff; // @[Math.scala 451:55:@72230.4]
  assign _T_526 = x753_sum_number[3:0]; // @[FixedPoint.scala 18:52:@72231.4]
  assign _T_532 = _T_526 != 4'h0; // @[Math.scala 451:110:@72233.4]
  assign _T_533 = _T_525 & _T_532; // @[Math.scala 451:94:@72234.4]
  assign _T_535 = {_T_518,_T_519}; // @[Cat.scala 30:58:@72236.4]
  assign x680_1_number = _T_533 ? 32'h0 : _T_535; // @[Math.scala 454:20:@72237.4]
  assign _GEN_1 = {{4'd0}, x680_1_number}; // @[Math.scala 461:32:@72242.4]
  assign _T_540 = _GEN_1 << 4; // @[Math.scala 461:32:@72242.4]
  assign _GEN_2 = {{6'd0}, x680_1_number}; // @[Math.scala 461:32:@72247.4]
  assign _T_543 = _GEN_2 << 6; // @[Math.scala 461:32:@72247.4]
  assign x685_sum_number = x685_sum_1_io_result; // @[Math.scala 154:22:@72281.4 Math.scala 155:14:@72282.4]
  assign _T_563 = x685_sum_number[31]; // @[FixedPoint.scala 50:25:@72286.4]
  assign _T_567 = _T_563 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@72288.4]
  assign _T_568 = x685_sum_number[31:4]; // @[FixedPoint.scala 18:52:@72289.4]
  assign _T_574 = _T_568 == 28'hfffffff; // @[Math.scala 451:55:@72291.4]
  assign _T_575 = x685_sum_number[3:0]; // @[FixedPoint.scala 18:52:@72292.4]
  assign _T_581 = _T_575 != 4'h0; // @[Math.scala 451:110:@72294.4]
  assign _T_582 = _T_574 & _T_581; // @[Math.scala 451:94:@72295.4]
  assign _T_584 = {_T_567,_T_568}; // @[Cat.scala 30:58:@72297.4]
  assign x686_1_number = _T_582 ? 32'h0 : _T_584; // @[Math.scala 454:20:@72298.4]
  assign _GEN_3 = {{4'd0}, x686_1_number}; // @[Math.scala 461:32:@72303.4]
  assign _GEN_4 = {{6'd0}, x686_1_number}; // @[Math.scala 461:32:@72315.4]
  assign _T_596 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@72321.4 package.scala 96:25:@72322.4]
  assign x755_1_number = _T_596[31:0]; // @[Math.scala 459:22:@72314.4 Math.scala 461:14:@72323.4]
  assign x802_x691_sum_D1_number = RetimeWrapper_3_io_out; // @[package.scala 96:25:@72361.4 package.scala 96:25:@72362.4]
  assign x692_tuple = {1'h0,x755_1_number,x802_x691_sum_D1_number}; // @[Cat.scala 30:58:@72366.4]
  assign _T_626 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@72385.4 package.scala 96:25:@72386.4]
  assign _T_628 = io_rr ? _T_626 : 1'h0; // @[implicits.scala 56:10:@72387.4]
  assign x803_x693_D4 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@72375.4 package.scala 96:25:@72376.4]
  assign _T_629 = _T_628 & x803_x693_D4; // @[sm_x698_inr_UnitPipe.scala 116:121:@72388.4]
  assign _T_633 = ~ io_sigsIn_break; // @[sm_x698_inr_UnitPipe.scala 123:116:@72395.4]
  assign _T_639 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@72404.4 package.scala 96:25:@72405.4]
  assign _T_641 = io_rr ? _T_639 : 1'h0; // @[implicits.scala 56:10:@72406.4]
  assign _T_642 = _T_633 & _T_641; // @[sm_x698_inr_UnitPipe.scala 123:133:@72407.4]
  assign _T_644 = _T_642 & _T_633; // @[sm_x698_inr_UnitPipe.scala 123:230:@72409.4]
  assign _T_654 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@72424.4 package.scala 96:25:@72425.4]
  assign _T_656 = io_rr ? _T_654 : 1'h0; // @[implicits.scala 56:10:@72426.4]
  assign _T_657 = _T_633 & _T_656; // @[sm_x698_inr_UnitPipe.scala 128:133:@72427.4]
  assign _T_659 = _T_657 & _T_633; // @[sm_x698_inr_UnitPipe.scala 128:230:@72429.4]
  assign _T_669 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@72444.4 package.scala 96:25:@72445.4]
  assign _T_671 = io_rr ? _T_669 : 1'h0; // @[implicits.scala 56:10:@72446.4]
  assign _T_672 = _T_633 & _T_671; // @[sm_x698_inr_UnitPipe.scala 133:133:@72447.4]
  assign _T_674 = _T_672 & _T_633; // @[sm_x698_inr_UnitPipe.scala 133:230:@72449.4]
  assign _T_591 = RetimeWrapper_io_out; // @[package.scala 96:25:@72309.4 package.scala 96:25:@72310.4]
  assign io_in_x677_reg_wPort_0_data_0 = x684_sum_1_io_result; // @[MemInterfaceType.scala 90:56:@72432.4]
  assign io_in_x677_reg_wPort_0_reset = io_in_x677_reg_reset; // @[MemInterfaceType.scala 91:23:@72433.4]
  assign io_in_x677_reg_wPort_0_en_0 = _T_659 & io_sigsIn_backpressure; // @[MemInterfaceType.scala 93:57:@72434.4]
  assign io_in_x677_reg_reset = 1'h0;
  assign io_in_x678_reg_wPort_0_data_0 = _T_591[31:0]; // @[MemInterfaceType.scala 90:56:@72452.4]
  assign io_in_x678_reg_wPort_0_reset = io_in_x678_reg_reset; // @[MemInterfaceType.scala 91:23:@72453.4]
  assign io_in_x678_reg_wPort_0_en_0 = _T_674 & io_sigsIn_backpressure; // @[MemInterfaceType.scala 93:57:@72454.4]
  assign io_in_x678_reg_reset = 1'h0;
  assign io_in_x669_valid = _T_629 & io_sigsIn_backpressure; // @[sm_x698_inr_UnitPipe.scala 116:18:@72390.4]
  assign io_in_x669_bits_addr = x692_tuple[63:0]; // @[sm_x698_inr_UnitPipe.scala 117:22:@72392.4]
  assign io_in_x669_bits_size = x692_tuple[95:64]; // @[sm_x698_inr_UnitPipe.scala 118:22:@72394.4]
  assign io_in_x676_reg_wPort_0_data_0 = x683_sub_1_io_result; // @[MemInterfaceType.scala 90:56:@72412.4]
  assign io_in_x676_reg_wPort_0_reset = io_in_x676_reg_reset; // @[MemInterfaceType.scala 91:23:@72413.4]
  assign io_in_x676_reg_wPort_0_en_0 = _T_644 & io_sigsIn_backpressure; // @[MemInterfaceType.scala 93:57:@72414.4]
  assign io_in_x676_reg_reset = 1'h0;
  assign x753_sum_1_clock = clock; // @[:@72215.4]
  assign x753_sum_1_reset = reset; // @[:@72216.4]
  assign x753_sum_1_io_a = _T_508[31:0]; // @[Math.scala 151:17:@72217.4]
  assign x753_sum_1_io_b = io_in_b674_number; // @[Math.scala 152:17:@72218.4]
  assign x753_sum_1_io_flow = io_in_x669_ready; // @[Math.scala 153:20:@72219.4]
  assign x683_sub_1_clock = clock; // @[:@72252.4]
  assign x683_sub_1_reset = reset; // @[:@72253.4]
  assign x683_sub_1_io_a = x753_sum_1_io_result; // @[Math.scala 192:17:@72254.4]
  assign x683_sub_1_io_b = _T_540[31:0]; // @[Math.scala 193:17:@72255.4]
  assign x683_sub_1_io_flow = io_in_x669_ready; // @[Math.scala 194:20:@72256.4]
  assign x684_sum_1_clock = clock; // @[:@72264.4]
  assign x684_sum_1_reset = reset; // @[:@72265.4]
  assign x684_sum_1_io_a = x683_sub_1_io_result; // @[Math.scala 151:17:@72266.4]
  assign x684_sum_1_io_b = 32'h3; // @[Math.scala 152:17:@72267.4]
  assign x684_sum_1_io_flow = io_in_x669_ready; // @[Math.scala 153:20:@72268.4]
  assign x685_sum_1_clock = clock; // @[:@72276.4]
  assign x685_sum_1_reset = reset; // @[:@72277.4]
  assign x685_sum_1_io_a = x683_sub_1_io_result; // @[Math.scala 151:17:@72278.4]
  assign x685_sum_1_io_b = 32'h12; // @[Math.scala 152:17:@72279.4]
  assign x685_sum_1_io_flow = io_in_x669_ready; // @[Math.scala 153:20:@72280.4]
  assign RetimeWrapper_clock = clock; // @[:@72305.4]
  assign RetimeWrapper_reset = reset; // @[:@72306.4]
  assign RetimeWrapper_io_flow = io_in_x669_ready; // @[package.scala 95:18:@72308.4]
  assign RetimeWrapper_io_in = _GEN_3 << 4; // @[package.scala 94:16:@72307.4]
  assign RetimeWrapper_1_clock = clock; // @[:@72317.4]
  assign RetimeWrapper_1_reset = reset; // @[:@72318.4]
  assign RetimeWrapper_1_io_flow = io_in_x669_ready; // @[package.scala 95:18:@72320.4]
  assign RetimeWrapper_1_io_in = _GEN_4 << 6; // @[package.scala 94:16:@72319.4]
  assign x689_1_io_b = _T_543[31:0]; // @[Math.scala 721:17:@72329.4]
  assign RetimeWrapper_2_clock = clock; // @[:@72337.4]
  assign RetimeWrapper_2_reset = reset; // @[:@72338.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@72340.4]
  assign RetimeWrapper_2_io_in = io_in_x470_out_host_number; // @[package.scala 94:16:@72339.4]
  assign x691_sum_1_clock = clock; // @[:@72346.4]
  assign x691_sum_1_reset = reset; // @[:@72347.4]
  assign x691_sum_1_io_a = x689_1_io_result; // @[Math.scala 151:17:@72348.4]
  assign x691_sum_1_io_b = RetimeWrapper_2_io_out; // @[Math.scala 152:17:@72349.4]
  assign x691_sum_1_io_flow = io_in_x669_ready; // @[Math.scala 153:20:@72350.4]
  assign RetimeWrapper_3_clock = clock; // @[:@72357.4]
  assign RetimeWrapper_3_reset = reset; // @[:@72358.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@72360.4]
  assign RetimeWrapper_3_io_in = x691_sum_1_io_result; // @[package.scala 94:16:@72359.4]
  assign RetimeWrapper_4_clock = clock; // @[:@72371.4]
  assign RetimeWrapper_4_reset = reset; // @[:@72372.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@72374.4]
  assign RetimeWrapper_4_io_in = 1'h1; // @[package.scala 94:16:@72373.4]
  assign RetimeWrapper_5_clock = clock; // @[:@72381.4]
  assign RetimeWrapper_5_reset = reset; // @[:@72382.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@72384.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@72383.4]
  assign RetimeWrapper_6_clock = clock; // @[:@72400.4]
  assign RetimeWrapper_6_reset = reset; // @[:@72401.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@72403.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@72402.4]
  assign RetimeWrapper_7_clock = clock; // @[:@72420.4]
  assign RetimeWrapper_7_reset = reset; // @[:@72421.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@72423.4]
  assign RetimeWrapper_7_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@72422.4]
  assign RetimeWrapper_8_clock = clock; // @[:@72440.4]
  assign RetimeWrapper_8_reset = reset; // @[:@72441.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@72443.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@72442.4]
endmodule
module x717_inr_Foreach_kernelx717_inr_Foreach_concrete1( // @[:@73821.2]
  input         clock, // @[:@73822.4]
  input         reset, // @[:@73823.4]
  input  [31:0] io_in_x677_reg_rPort_0_output_0, // @[:@73824.4]
  input         io_in_x670_ready, // @[:@73824.4]
  output        io_in_x670_valid, // @[:@73824.4]
  output [31:0] io_in_x670_bits_wdata_0, // @[:@73824.4]
  output        io_in_x670_bits_wstrb, // @[:@73824.4]
  input  [31:0] io_in_b674_number, // @[:@73824.4]
  output [8:0]  io_in_x539_out_sram_0_rPort_0_ofs_0, // @[:@73824.4]
  output        io_in_x539_out_sram_0_rPort_0_en_0, // @[:@73824.4]
  output        io_in_x539_out_sram_0_rPort_0_backpressure, // @[:@73824.4]
  input  [31:0] io_in_x539_out_sram_0_rPort_0_output_0, // @[:@73824.4]
  input  [31:0] io_in_x676_reg_rPort_0_output_0, // @[:@73824.4]
  input         io_sigsIn_backpressure, // @[:@73824.4]
  input         io_sigsIn_datapathEn, // @[:@73824.4]
  input         io_sigsIn_break, // @[:@73824.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@73824.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@73824.4]
  input         io_rr // @[:@73824.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@73877.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@73877.4]
  wire  x709_sub_1_clock; // @[Math.scala 191:24:@73930.4]
  wire  x709_sub_1_reset; // @[Math.scala 191:24:@73930.4]
  wire [31:0] x709_sub_1_io_a; // @[Math.scala 191:24:@73930.4]
  wire [31:0] x709_sub_1_io_b; // @[Math.scala 191:24:@73930.4]
  wire  x709_sub_1_io_flow; // @[Math.scala 191:24:@73930.4]
  wire [31:0] x709_sub_1_io_result; // @[Math.scala 191:24:@73930.4]
  wire  x757_sum_1_clock; // @[Math.scala 150:24:@73945.4]
  wire  x757_sum_1_reset; // @[Math.scala 150:24:@73945.4]
  wire [31:0] x757_sum_1_io_a; // @[Math.scala 150:24:@73945.4]
  wire [31:0] x757_sum_1_io_b; // @[Math.scala 150:24:@73945.4]
  wire  x757_sum_1_io_flow; // @[Math.scala 150:24:@73945.4]
  wire [31:0] x757_sum_1_io_result; // @[Math.scala 150:24:@73945.4]
  wire  x712_sum_1_clock; // @[Math.scala 150:24:@73955.4]
  wire  x712_sum_1_reset; // @[Math.scala 150:24:@73955.4]
  wire [31:0] x712_sum_1_io_a; // @[Math.scala 150:24:@73955.4]
  wire [31:0] x712_sum_1_io_b; // @[Math.scala 150:24:@73955.4]
  wire  x712_sum_1_io_flow; // @[Math.scala 150:24:@73955.4]
  wire [31:0] x712_sum_1_io_result; // @[Math.scala 150:24:@73955.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@73966.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@73966.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@73966.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@73966.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@73966.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@73976.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@73976.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@73976.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@73976.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@73976.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@73988.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@73988.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@73988.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@73988.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@73988.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@74000.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@74000.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@74000.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@74000.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@74000.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@74021.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@74021.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@74021.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@74021.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@74021.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@74034.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@74034.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@74034.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@74034.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@74034.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@74044.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@74044.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@74044.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@74044.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@74044.4]
  wire  _T_523; // @[sm_x717_inr_Foreach.scala 80:119:@73889.4]
  wire [31:0] _T_535; // @[Math.scala 493:37:@73903.4]
  wire [31:0] b702_number; // @[Math.scala 723:22:@73882.4 Math.scala 724:14:@73883.4]
  wire [31:0] _T_536; // @[Math.scala 493:51:@73904.4]
  wire  x705; // @[Math.scala 493:44:@73905.4]
  wire [31:0] _T_555; // @[Math.scala 476:50:@73923.4]
  wire  x707; // @[Math.scala 476:44:@73924.4]
  wire [32:0] _GEN_0; // @[Math.scala 461:32:@73941.4]
  wire [32:0] _T_564; // @[Math.scala 461:32:@73941.4]
  wire  _T_594; // @[package.scala 96:25:@73993.4 package.scala 96:25:@73994.4]
  wire  _T_596; // @[implicits.scala 56:10:@73995.4]
  wire  _T_598; // @[sm_x717_inr_Foreach.scala 112:111:@73997.4]
  wire  _T_603; // @[package.scala 96:25:@74005.4 package.scala 96:25:@74006.4]
  wire  _T_605; // @[implicits.scala 56:10:@74007.4]
  wire  _T_606; // @[sm_x717_inr_Foreach.scala 112:131:@74008.4]
  wire  x805_x708_D2; // @[package.scala 96:25:@73981.4 package.scala 96:25:@73982.4]
  wire  _T_607; // @[sm_x717_inr_Foreach.scala 112:228:@74009.4]
  wire  x804_b703_D2; // @[package.scala 96:25:@73971.4 package.scala 96:25:@73972.4]
  wire  x806_x708_D4; // @[package.scala 96:25:@74026.4 package.scala 96:25:@74027.4]
  wire [32:0] x715_tuple; // @[Cat.scala 30:58:@74030.4]
  wire  _T_626; // @[package.scala 96:25:@74049.4 package.scala 96:25:@74050.4]
  wire  _T_628; // @[implicits.scala 56:10:@74051.4]
  wire  x807_b703_D4; // @[package.scala 96:25:@74039.4 package.scala 96:25:@74040.4]
  wire  _T_629; // @[sm_x717_inr_Foreach.scala 123:121:@74052.4]
  wire [31:0] x712_sum_number; // @[Math.scala 154:22:@73961.4 Math.scala 155:14:@73962.4]
  _ _ ( // @[Math.scala 720:24:@73877.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x485_sub x709_sub_1 ( // @[Math.scala 191:24:@73930.4]
    .clock(x709_sub_1_clock),
    .reset(x709_sub_1_reset),
    .io_a(x709_sub_1_io_a),
    .io_b(x709_sub_1_io_b),
    .io_flow(x709_sub_1_io_flow),
    .io_result(x709_sub_1_io_result)
  );
  x739_sum x757_sum_1 ( // @[Math.scala 150:24:@73945.4]
    .clock(x757_sum_1_clock),
    .reset(x757_sum_1_reset),
    .io_a(x757_sum_1_io_a),
    .io_b(x757_sum_1_io_b),
    .io_flow(x757_sum_1_io_flow),
    .io_result(x757_sum_1_io_result)
  );
  x739_sum x712_sum_1 ( // @[Math.scala 150:24:@73955.4]
    .clock(x712_sum_1_clock),
    .reset(x712_sum_1_reset),
    .io_a(x712_sum_1_io_a),
    .io_b(x712_sum_1_io_b),
    .io_flow(x712_sum_1_io_flow),
    .io_result(x712_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@73966.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@73976.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@73988.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@74000.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@74021.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_5 ( // @[package.scala 93:22:@74034.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_6 ( // @[package.scala 93:22:@74044.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  assign _T_523 = ~ io_sigsIn_break; // @[sm_x717_inr_Foreach.scala 80:119:@73889.4]
  assign _T_535 = $signed(io_in_x676_reg_rPort_0_output_0); // @[Math.scala 493:37:@73903.4]
  assign b702_number = __io_result; // @[Math.scala 723:22:@73882.4 Math.scala 724:14:@73883.4]
  assign _T_536 = $signed(b702_number); // @[Math.scala 493:51:@73904.4]
  assign x705 = $signed(_T_535) <= $signed(_T_536); // @[Math.scala 493:44:@73905.4]
  assign _T_555 = $signed(io_in_x677_reg_rPort_0_output_0); // @[Math.scala 476:50:@73923.4]
  assign x707 = $signed(_T_536) < $signed(_T_555); // @[Math.scala 476:44:@73924.4]
  assign _GEN_0 = {{1'd0}, io_in_b674_number}; // @[Math.scala 461:32:@73941.4]
  assign _T_564 = _GEN_0 << 1; // @[Math.scala 461:32:@73941.4]
  assign _T_594 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@73993.4 package.scala 96:25:@73994.4]
  assign _T_596 = io_rr ? _T_594 : 1'h0; // @[implicits.scala 56:10:@73995.4]
  assign _T_598 = _T_596 & _T_523; // @[sm_x717_inr_Foreach.scala 112:111:@73997.4]
  assign _T_603 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@74005.4 package.scala 96:25:@74006.4]
  assign _T_605 = io_rr ? _T_603 : 1'h0; // @[implicits.scala 56:10:@74007.4]
  assign _T_606 = _T_598 & _T_605; // @[sm_x717_inr_Foreach.scala 112:131:@74008.4]
  assign x805_x708_D2 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@73981.4 package.scala 96:25:@73982.4]
  assign _T_607 = _T_606 & x805_x708_D2; // @[sm_x717_inr_Foreach.scala 112:228:@74009.4]
  assign x804_b703_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@73971.4 package.scala 96:25:@73972.4]
  assign x806_x708_D4 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@74026.4 package.scala 96:25:@74027.4]
  assign x715_tuple = {x806_x708_D4,io_in_x539_out_sram_0_rPort_0_output_0}; // @[Cat.scala 30:58:@74030.4]
  assign _T_626 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@74049.4 package.scala 96:25:@74050.4]
  assign _T_628 = io_rr ? _T_626 : 1'h0; // @[implicits.scala 56:10:@74051.4]
  assign x807_b703_D4 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@74039.4 package.scala 96:25:@74040.4]
  assign _T_629 = _T_628 & x807_b703_D4; // @[sm_x717_inr_Foreach.scala 123:121:@74052.4]
  assign x712_sum_number = x712_sum_1_io_result; // @[Math.scala 154:22:@73961.4 Math.scala 155:14:@73962.4]
  assign io_in_x670_valid = _T_629 & io_sigsIn_backpressure; // @[sm_x717_inr_Foreach.scala 123:18:@74054.4]
  assign io_in_x670_bits_wdata_0 = x715_tuple[31:0]; // @[sm_x717_inr_Foreach.scala 124:26:@74056.4]
  assign io_in_x670_bits_wstrb = x715_tuple[32]; // @[sm_x717_inr_Foreach.scala 125:23:@74058.4]
  assign io_in_x539_out_sram_0_rPort_0_ofs_0 = x712_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@74013.4]
  assign io_in_x539_out_sram_0_rPort_0_en_0 = _T_607 & x804_b703_D2; // @[MemInterfaceType.scala 110:79:@74015.4]
  assign io_in_x539_out_sram_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@74014.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@73880.4]
  assign x709_sub_1_clock = clock; // @[:@73931.4]
  assign x709_sub_1_reset = reset; // @[:@73932.4]
  assign x709_sub_1_io_a = __io_result; // @[Math.scala 192:17:@73933.4]
  assign x709_sub_1_io_b = io_in_x676_reg_rPort_0_output_0; // @[Math.scala 193:17:@73934.4]
  assign x709_sub_1_io_flow = io_in_x670_ready; // @[Math.scala 194:20:@73935.4]
  assign x757_sum_1_clock = clock; // @[:@73946.4]
  assign x757_sum_1_reset = reset; // @[:@73947.4]
  assign x757_sum_1_io_a = _T_564[31:0]; // @[Math.scala 151:17:@73948.4]
  assign x757_sum_1_io_b = io_in_b674_number; // @[Math.scala 152:17:@73949.4]
  assign x757_sum_1_io_flow = io_in_x670_ready; // @[Math.scala 153:20:@73950.4]
  assign x712_sum_1_clock = clock; // @[:@73956.4]
  assign x712_sum_1_reset = reset; // @[:@73957.4]
  assign x712_sum_1_io_a = x757_sum_1_io_result; // @[Math.scala 151:17:@73958.4]
  assign x712_sum_1_io_b = x709_sub_1_io_result; // @[Math.scala 152:17:@73959.4]
  assign x712_sum_1_io_flow = io_in_x670_ready; // @[Math.scala 153:20:@73960.4]
  assign RetimeWrapper_clock = clock; // @[:@73967.4]
  assign RetimeWrapper_reset = reset; // @[:@73968.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@73970.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@73969.4]
  assign RetimeWrapper_1_clock = clock; // @[:@73977.4]
  assign RetimeWrapper_1_reset = reset; // @[:@73978.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@73980.4]
  assign RetimeWrapper_1_io_in = x705 & x707; // @[package.scala 94:16:@73979.4]
  assign RetimeWrapper_2_clock = clock; // @[:@73989.4]
  assign RetimeWrapper_2_reset = reset; // @[:@73990.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@73992.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@73991.4]
  assign RetimeWrapper_3_clock = clock; // @[:@74001.4]
  assign RetimeWrapper_3_reset = reset; // @[:@74002.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@74004.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@74003.4]
  assign RetimeWrapper_4_clock = clock; // @[:@74022.4]
  assign RetimeWrapper_4_reset = reset; // @[:@74023.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@74025.4]
  assign RetimeWrapper_4_io_in = x705 & x707; // @[package.scala 94:16:@74024.4]
  assign RetimeWrapper_5_clock = clock; // @[:@74035.4]
  assign RetimeWrapper_5_reset = reset; // @[:@74036.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@74038.4]
  assign RetimeWrapper_5_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@74037.4]
  assign RetimeWrapper_6_clock = clock; // @[:@74045.4]
  assign RetimeWrapper_6_reset = reset; // @[:@74046.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@74048.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@74047.4]
endmodule
module x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1( // @[:@74060.2]
  input         clock, // @[:@74061.4]
  input         reset, // @[:@74062.4]
  input         io_in_x670_ready, // @[:@74063.4]
  output        io_in_x670_valid, // @[:@74063.4]
  output [31:0] io_in_x670_bits_wdata_0, // @[:@74063.4]
  output        io_in_x670_bits_wstrb, // @[:@74063.4]
  input         io_in_x669_ready, // @[:@74063.4]
  output        io_in_x669_valid, // @[:@74063.4]
  output [63:0] io_in_x669_bits_addr, // @[:@74063.4]
  output [31:0] io_in_x669_bits_size, // @[:@74063.4]
  input  [31:0] io_in_b674_number, // @[:@74063.4]
  input  [63:0] io_in_x470_out_host_number, // @[:@74063.4]
  output [8:0]  io_in_x539_out_sram_0_rPort_0_ofs_0, // @[:@74063.4]
  output        io_in_x539_out_sram_0_rPort_0_en_0, // @[:@74063.4]
  output        io_in_x539_out_sram_0_rPort_0_backpressure, // @[:@74063.4]
  input  [31:0] io_in_x539_out_sram_0_rPort_0_output_0, // @[:@74063.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@74063.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@74063.4]
  input         io_sigsIn_smChildAcks_0, // @[:@74063.4]
  input         io_sigsIn_smChildAcks_1, // @[:@74063.4]
  output        io_sigsOut_smDoneIn_0, // @[:@74063.4]
  output        io_sigsOut_smDoneIn_1, // @[:@74063.4]
  output        io_sigsOut_smMaskIn_1, // @[:@74063.4]
  input         io_rr // @[:@74063.4]
);
  wire  x676_reg_clock; // @[m_x676_reg.scala 27:22:@74088.4]
  wire  x676_reg_reset; // @[m_x676_reg.scala 27:22:@74088.4]
  wire [31:0] x676_reg_io_rPort_0_output_0; // @[m_x676_reg.scala 27:22:@74088.4]
  wire [31:0] x676_reg_io_wPort_0_data_0; // @[m_x676_reg.scala 27:22:@74088.4]
  wire  x676_reg_io_wPort_0_reset; // @[m_x676_reg.scala 27:22:@74088.4]
  wire  x676_reg_io_wPort_0_en_0; // @[m_x676_reg.scala 27:22:@74088.4]
  wire  x677_reg_clock; // @[m_x677_reg.scala 27:22:@74105.4]
  wire  x677_reg_reset; // @[m_x677_reg.scala 27:22:@74105.4]
  wire [31:0] x677_reg_io_rPort_0_output_0; // @[m_x677_reg.scala 27:22:@74105.4]
  wire [31:0] x677_reg_io_wPort_0_data_0; // @[m_x677_reg.scala 27:22:@74105.4]
  wire  x677_reg_io_wPort_0_reset; // @[m_x677_reg.scala 27:22:@74105.4]
  wire  x677_reg_io_wPort_0_en_0; // @[m_x677_reg.scala 27:22:@74105.4]
  wire  x678_reg_clock; // @[m_x678_reg.scala 27:22:@74122.4]
  wire  x678_reg_reset; // @[m_x678_reg.scala 27:22:@74122.4]
  wire [31:0] x678_reg_io_rPort_0_output_0; // @[m_x678_reg.scala 27:22:@74122.4]
  wire [31:0] x678_reg_io_wPort_0_data_0; // @[m_x678_reg.scala 27:22:@74122.4]
  wire  x678_reg_io_wPort_0_reset; // @[m_x678_reg.scala 27:22:@74122.4]
  wire  x678_reg_io_wPort_0_en_0; // @[m_x678_reg.scala 27:22:@74122.4]
  wire  x698_inr_UnitPipe_sm_clock; // @[sm_x698_inr_UnitPipe.scala 34:18:@74175.4]
  wire  x698_inr_UnitPipe_sm_reset; // @[sm_x698_inr_UnitPipe.scala 34:18:@74175.4]
  wire  x698_inr_UnitPipe_sm_io_enable; // @[sm_x698_inr_UnitPipe.scala 34:18:@74175.4]
  wire  x698_inr_UnitPipe_sm_io_done; // @[sm_x698_inr_UnitPipe.scala 34:18:@74175.4]
  wire  x698_inr_UnitPipe_sm_io_doneLatch; // @[sm_x698_inr_UnitPipe.scala 34:18:@74175.4]
  wire  x698_inr_UnitPipe_sm_io_rst; // @[sm_x698_inr_UnitPipe.scala 34:18:@74175.4]
  wire  x698_inr_UnitPipe_sm_io_ctrDone; // @[sm_x698_inr_UnitPipe.scala 34:18:@74175.4]
  wire  x698_inr_UnitPipe_sm_io_datapathEn; // @[sm_x698_inr_UnitPipe.scala 34:18:@74175.4]
  wire  x698_inr_UnitPipe_sm_io_ctrInc; // @[sm_x698_inr_UnitPipe.scala 34:18:@74175.4]
  wire  x698_inr_UnitPipe_sm_io_ctrRst; // @[sm_x698_inr_UnitPipe.scala 34:18:@74175.4]
  wire  x698_inr_UnitPipe_sm_io_parentAck; // @[sm_x698_inr_UnitPipe.scala 34:18:@74175.4]
  wire  x698_inr_UnitPipe_sm_io_backpressure; // @[sm_x698_inr_UnitPipe.scala 34:18:@74175.4]
  wire  x698_inr_UnitPipe_sm_io_break; // @[sm_x698_inr_UnitPipe.scala 34:18:@74175.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@74233.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@74233.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@74233.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@74233.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@74233.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@74241.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@74241.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@74241.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@74241.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@74241.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_clock; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_reset; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire [31:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_data_0; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_reset; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_en_0; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_reset; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire [31:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_data_0; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_reset; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_en_0; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_reset; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_ready; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_valid; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire [63:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_bits_addr; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire [31:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_bits_size; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire [31:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_b674_number; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire [63:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x470_out_host_number; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire [31:0] x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_data_0; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_reset; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_en_0; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_reset; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_break; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_rr; // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
  wire  x701_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@74414.4]
  wire  x701_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@74414.4]
  wire [31:0] x701_ctrchain_io_setup_stops_0; // @[SpatialBlocks.scala 37:22:@74414.4]
  wire  x701_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@74414.4]
  wire  x701_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@74414.4]
  wire [31:0] x701_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@74414.4]
  wire  x701_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@74414.4]
  wire  x701_ctrchain_io_output_noop; // @[SpatialBlocks.scala 37:22:@74414.4]
  wire  x701_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@74414.4]
  wire  x717_inr_Foreach_sm_clock; // @[sm_x717_inr_Foreach.scala 34:18:@74469.4]
  wire  x717_inr_Foreach_sm_reset; // @[sm_x717_inr_Foreach.scala 34:18:@74469.4]
  wire  x717_inr_Foreach_sm_io_enable; // @[sm_x717_inr_Foreach.scala 34:18:@74469.4]
  wire  x717_inr_Foreach_sm_io_done; // @[sm_x717_inr_Foreach.scala 34:18:@74469.4]
  wire  x717_inr_Foreach_sm_io_doneLatch; // @[sm_x717_inr_Foreach.scala 34:18:@74469.4]
  wire  x717_inr_Foreach_sm_io_ctrDone; // @[sm_x717_inr_Foreach.scala 34:18:@74469.4]
  wire  x717_inr_Foreach_sm_io_datapathEn; // @[sm_x717_inr_Foreach.scala 34:18:@74469.4]
  wire  x717_inr_Foreach_sm_io_ctrInc; // @[sm_x717_inr_Foreach.scala 34:18:@74469.4]
  wire  x717_inr_Foreach_sm_io_ctrRst; // @[sm_x717_inr_Foreach.scala 34:18:@74469.4]
  wire  x717_inr_Foreach_sm_io_parentAck; // @[sm_x717_inr_Foreach.scala 34:18:@74469.4]
  wire  x717_inr_Foreach_sm_io_backpressure; // @[sm_x717_inr_Foreach.scala 34:18:@74469.4]
  wire  x717_inr_Foreach_sm_io_break; // @[sm_x717_inr_Foreach.scala 34:18:@74469.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@74498.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@74498.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@74498.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@74498.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@74498.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@74538.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@74538.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@74538.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@74538.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@74538.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@74546.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@74546.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@74546.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@74546.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@74546.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_clock; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_reset; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire [31:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x677_reg_rPort_0_output_0; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_ready; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_valid; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire [31:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_bits_wdata_0; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_bits_wstrb; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire [31:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_b674_number; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire [8:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_en_0; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire [31:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_output_0; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire [31:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x676_reg_rPort_0_output_0; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire [31:0] x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_rr; // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
  wire  _T_330; // @[package.scala 100:49:@74203.4]
  reg  _T_333; // @[package.scala 48:56:@74204.4]
  reg [31:0] _RAND_0;
  wire  _T_348; // @[package.scala 96:25:@74238.4 package.scala 96:25:@74239.4]
  wire  _T_354; // @[package.scala 96:25:@74246.4 package.scala 96:25:@74247.4]
  wire  _T_357; // @[SpatialBlocks.scala 137:99:@74249.4]
  wire [31:0] x737_rd_x678_number; // @[sm_x718_outr_UnitPipe.scala 92:30:@74400.4 sm_x718_outr_UnitPipe.scala 97:202:@74413.4]
  wire  _T_445; // @[package.scala 96:25:@74503.4 package.scala 96:25:@74504.4]
  wire  x717_inr_Foreach_mySignalsIn_mask; // @[sm_x718_outr_UnitPipe.scala 108:32:@74514.4]
  wire  _T_461; // @[package.scala 96:25:@74543.4 package.scala 96:25:@74544.4]
  wire  _T_467; // @[package.scala 96:25:@74551.4 package.scala 96:25:@74552.4]
  wire  _T_470; // @[SpatialBlocks.scala 137:99:@74554.4]
  wire  _T_472; // @[SpatialBlocks.scala 156:36:@74563.4]
  wire  _T_473; // @[SpatialBlocks.scala 156:78:@74564.4]
  x505_reg x676_reg ( // @[m_x676_reg.scala 27:22:@74088.4]
    .clock(x676_reg_clock),
    .reset(x676_reg_reset),
    .io_rPort_0_output_0(x676_reg_io_rPort_0_output_0),
    .io_wPort_0_data_0(x676_reg_io_wPort_0_data_0),
    .io_wPort_0_reset(x676_reg_io_wPort_0_reset),
    .io_wPort_0_en_0(x676_reg_io_wPort_0_en_0)
  );
  x505_reg x677_reg ( // @[m_x677_reg.scala 27:22:@74105.4]
    .clock(x677_reg_clock),
    .reset(x677_reg_reset),
    .io_rPort_0_output_0(x677_reg_io_rPort_0_output_0),
    .io_wPort_0_data_0(x677_reg_io_wPort_0_data_0),
    .io_wPort_0_reset(x677_reg_io_wPort_0_reset),
    .io_wPort_0_en_0(x677_reg_io_wPort_0_en_0)
  );
  x505_reg x678_reg ( // @[m_x678_reg.scala 27:22:@74122.4]
    .clock(x678_reg_clock),
    .reset(x678_reg_reset),
    .io_rPort_0_output_0(x678_reg_io_rPort_0_output_0),
    .io_wPort_0_data_0(x678_reg_io_wPort_0_data_0),
    .io_wPort_0_reset(x678_reg_io_wPort_0_reset),
    .io_wPort_0_en_0(x678_reg_io_wPort_0_en_0)
  );
  x499_inr_Foreach_sm x698_inr_UnitPipe_sm ( // @[sm_x698_inr_UnitPipe.scala 34:18:@74175.4]
    .clock(x698_inr_UnitPipe_sm_clock),
    .reset(x698_inr_UnitPipe_sm_reset),
    .io_enable(x698_inr_UnitPipe_sm_io_enable),
    .io_done(x698_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x698_inr_UnitPipe_sm_io_doneLatch),
    .io_rst(x698_inr_UnitPipe_sm_io_rst),
    .io_ctrDone(x698_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x698_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x698_inr_UnitPipe_sm_io_ctrInc),
    .io_ctrRst(x698_inr_UnitPipe_sm_io_ctrRst),
    .io_parentAck(x698_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x698_inr_UnitPipe_sm_io_backpressure),
    .io_break(x698_inr_UnitPipe_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@74233.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@74241.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1 x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1 ( // @[sm_x698_inr_UnitPipe.scala 135:24:@74270.4]
    .clock(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_clock),
    .reset(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_reset),
    .io_in_x677_reg_wPort_0_data_0(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_data_0),
    .io_in_x677_reg_wPort_0_reset(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_reset),
    .io_in_x677_reg_wPort_0_en_0(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_en_0),
    .io_in_x677_reg_reset(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_reset),
    .io_in_x678_reg_wPort_0_data_0(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_data_0),
    .io_in_x678_reg_wPort_0_reset(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_reset),
    .io_in_x678_reg_wPort_0_en_0(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_en_0),
    .io_in_x678_reg_reset(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_reset),
    .io_in_x669_ready(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_ready),
    .io_in_x669_valid(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_valid),
    .io_in_x669_bits_addr(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_bits_addr),
    .io_in_x669_bits_size(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_bits_size),
    .io_in_b674_number(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_b674_number),
    .io_in_x470_out_host_number(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x470_out_host_number),
    .io_in_x676_reg_wPort_0_data_0(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_data_0),
    .io_in_x676_reg_wPort_0_reset(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_reset),
    .io_in_x676_reg_wPort_0_en_0(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_en_0),
    .io_in_x676_reg_reset(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_reset),
    .io_sigsIn_backpressure(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_break),
    .io_rr(x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_rr)
  );
  x519_ctrchain x701_ctrchain ( // @[SpatialBlocks.scala 37:22:@74414.4]
    .clock(x701_ctrchain_clock),
    .reset(x701_ctrchain_reset),
    .io_setup_stops_0(x701_ctrchain_io_setup_stops_0),
    .io_input_reset(x701_ctrchain_io_input_reset),
    .io_input_enable(x701_ctrchain_io_input_enable),
    .io_output_counts_0(x701_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x701_ctrchain_io_output_oobs_0),
    .io_output_noop(x701_ctrchain_io_output_noop),
    .io_output_done(x701_ctrchain_io_output_done)
  );
  x652_inr_Foreach_sm x717_inr_Foreach_sm ( // @[sm_x717_inr_Foreach.scala 34:18:@74469.4]
    .clock(x717_inr_Foreach_sm_clock),
    .reset(x717_inr_Foreach_sm_reset),
    .io_enable(x717_inr_Foreach_sm_io_enable),
    .io_done(x717_inr_Foreach_sm_io_done),
    .io_doneLatch(x717_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x717_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x717_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x717_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x717_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x717_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x717_inr_Foreach_sm_io_backpressure),
    .io_break(x717_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@74498.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@74538.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@74546.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x717_inr_Foreach_kernelx717_inr_Foreach_concrete1 x717_inr_Foreach_kernelx717_inr_Foreach_concrete1 ( // @[sm_x717_inr_Foreach.scala 127:24:@74580.4]
    .clock(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_clock),
    .reset(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_reset),
    .io_in_x677_reg_rPort_0_output_0(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x677_reg_rPort_0_output_0),
    .io_in_x670_ready(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_ready),
    .io_in_x670_valid(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_valid),
    .io_in_x670_bits_wdata_0(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_bits_wdata_0),
    .io_in_x670_bits_wstrb(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_bits_wstrb),
    .io_in_b674_number(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_b674_number),
    .io_in_x539_out_sram_0_rPort_0_ofs_0(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0),
    .io_in_x539_out_sram_0_rPort_0_en_0(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_en_0),
    .io_in_x539_out_sram_0_rPort_0_backpressure(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure),
    .io_in_x539_out_sram_0_rPort_0_output_0(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_output_0),
    .io_in_x676_reg_rPort_0_output_0(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x676_reg_rPort_0_output_0),
    .io_sigsIn_backpressure(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_rr)
  );
  assign _T_330 = x698_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@74203.4]
  assign _T_348 = RetimeWrapper_io_out; // @[package.scala 96:25:@74238.4 package.scala 96:25:@74239.4]
  assign _T_354 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@74246.4 package.scala 96:25:@74247.4]
  assign _T_357 = ~ _T_354; // @[SpatialBlocks.scala 137:99:@74249.4]
  assign x737_rd_x678_number = x678_reg_io_rPort_0_output_0; // @[sm_x718_outr_UnitPipe.scala 92:30:@74400.4 sm_x718_outr_UnitPipe.scala 97:202:@74413.4]
  assign _T_445 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@74503.4 package.scala 96:25:@74504.4]
  assign x717_inr_Foreach_mySignalsIn_mask = ~ x701_ctrchain_io_output_noop; // @[sm_x718_outr_UnitPipe.scala 108:32:@74514.4]
  assign _T_461 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@74543.4 package.scala 96:25:@74544.4]
  assign _T_467 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@74551.4 package.scala 96:25:@74552.4]
  assign _T_470 = ~ _T_467; // @[SpatialBlocks.scala 137:99:@74554.4]
  assign _T_472 = x717_inr_Foreach_sm_io_datapathEn & x717_inr_Foreach_mySignalsIn_mask; // @[SpatialBlocks.scala 156:36:@74563.4]
  assign _T_473 = ~ x717_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 156:78:@74564.4]
  assign io_in_x670_valid = x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_valid; // @[sm_x717_inr_Foreach.scala 57:23:@74662.4]
  assign io_in_x670_bits_wdata_0 = x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_bits_wdata_0; // @[sm_x717_inr_Foreach.scala 57:23:@74661.4]
  assign io_in_x670_bits_wstrb = x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_bits_wstrb; // @[sm_x717_inr_Foreach.scala 57:23:@74660.4]
  assign io_in_x669_valid = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_valid; // @[sm_x698_inr_UnitPipe.scala 60:23:@74362.4]
  assign io_in_x669_bits_addr = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_bits_addr; // @[sm_x698_inr_UnitPipe.scala 60:23:@74361.4]
  assign io_in_x669_bits_size = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_bits_size; // @[sm_x698_inr_UnitPipe.scala 60:23:@74360.4]
  assign io_in_x539_out_sram_0_rPort_0_ofs_0 = x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@74668.4]
  assign io_in_x539_out_sram_0_rPort_0_en_0 = x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@74667.4]
  assign io_in_x539_out_sram_0_rPort_0_backpressure = x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@74666.4]
  assign io_sigsOut_smDoneIn_0 = x698_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 155:56:@74256.4]
  assign io_sigsOut_smDoneIn_1 = x717_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@74561.4]
  assign io_sigsOut_smMaskIn_1 = ~ x701_ctrchain_io_output_noop; // @[SpatialBlocks.scala 155:86:@74562.4]
  assign x676_reg_clock = clock; // @[:@74089.4]
  assign x676_reg_reset = reset; // @[:@74090.4]
  assign x676_reg_io_wPort_0_data_0 = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@74370.4]
  assign x676_reg_io_wPort_0_reset = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_reset; // @[MemInterfaceType.scala 67:44:@74369.4]
  assign x676_reg_io_wPort_0_en_0 = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x676_reg_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@74366.4]
  assign x677_reg_clock = clock; // @[:@74106.4]
  assign x677_reg_reset = reset; // @[:@74107.4]
  assign x677_reg_io_wPort_0_data_0 = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@74350.4]
  assign x677_reg_io_wPort_0_reset = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_reset; // @[MemInterfaceType.scala 67:44:@74349.4]
  assign x677_reg_io_wPort_0_en_0 = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x677_reg_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@74346.4]
  assign x678_reg_clock = clock; // @[:@74123.4]
  assign x678_reg_reset = reset; // @[:@74124.4]
  assign x678_reg_io_wPort_0_data_0 = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@74357.4]
  assign x678_reg_io_wPort_0_reset = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_reset; // @[MemInterfaceType.scala 67:44:@74356.4]
  assign x678_reg_io_wPort_0_en_0 = x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x678_reg_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@74353.4]
  assign x698_inr_UnitPipe_sm_clock = clock; // @[:@74176.4]
  assign x698_inr_UnitPipe_sm_reset = reset; // @[:@74177.4]
  assign x698_inr_UnitPipe_sm_io_enable = _T_348 & _T_357; // @[SpatialBlocks.scala 139:18:@74253.4]
  assign x698_inr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 133:15:@74228.4]
  assign x698_inr_UnitPipe_sm_io_ctrDone = x698_inr_UnitPipe_sm_io_ctrInc & _T_333; // @[sm_x718_outr_UnitPipe.scala 84:39:@74207.4]
  assign x698_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@74255.4]
  assign x698_inr_UnitPipe_sm_io_backpressure = io_in_x669_ready | x698_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 132:24:@74227.4]
  assign x698_inr_UnitPipe_sm_io_break = 1'h0; // @[sm_x718_outr_UnitPipe.scala 88:37:@74214.4]
  assign RetimeWrapper_clock = clock; // @[:@74234.4]
  assign RetimeWrapper_reset = reset; // @[:@74235.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@74237.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@74236.4]
  assign RetimeWrapper_1_clock = clock; // @[:@74242.4]
  assign RetimeWrapper_1_reset = reset; // @[:@74243.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@74245.4]
  assign RetimeWrapper_1_io_in = x698_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@74244.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_clock = clock; // @[:@74271.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_reset = reset; // @[:@74272.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x669_ready = io_in_x669_ready; // @[sm_x698_inr_UnitPipe.scala 60:23:@74363.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_b674_number = io_in_b674_number; // @[sm_x698_inr_UnitPipe.scala 61:23:@74364.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_in_x470_out_host_number = io_in_x470_out_host_number; // @[sm_x698_inr_UnitPipe.scala 62:32:@74365.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x669_ready | x698_inr_UnitPipe_sm_io_doneLatch; // @[sm_x698_inr_UnitPipe.scala 140:22:@74387.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x698_inr_UnitPipe_sm_io_datapathEn; // @[sm_x698_inr_UnitPipe.scala 140:22:@74385.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_sigsIn_break = x698_inr_UnitPipe_sm_io_break; // @[sm_x698_inr_UnitPipe.scala 140:22:@74383.4]
  assign x698_inr_UnitPipe_kernelx698_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x698_inr_UnitPipe.scala 139:18:@74373.4]
  assign x701_ctrchain_clock = clock; // @[:@74415.4]
  assign x701_ctrchain_reset = reset; // @[:@74416.4]
  assign x701_ctrchain_io_setup_stops_0 = $signed(x737_rd_x678_number); // @[SpatialBlocks.scala 40:87:@74430.4]
  assign x701_ctrchain_io_input_reset = x717_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@74579.4]
  assign x701_ctrchain_io_input_enable = x717_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 158:42:@74578.4]
  assign x717_inr_Foreach_sm_clock = clock; // @[:@74470.4]
  assign x717_inr_Foreach_sm_reset = reset; // @[:@74471.4]
  assign x717_inr_Foreach_sm_io_enable = _T_461 & _T_470; // @[SpatialBlocks.scala 139:18:@74558.4]
  assign x717_inr_Foreach_sm_io_ctrDone = io_rr ? _T_445 : 1'h0; // @[sm_x718_outr_UnitPipe.scala 103:38:@74506.4]
  assign x717_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 141:21:@74560.4]
  assign x717_inr_Foreach_sm_io_backpressure = io_in_x670_ready | x717_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 132:24:@74532.4]
  assign x717_inr_Foreach_sm_io_break = 1'h0; // @[sm_x718_outr_UnitPipe.scala 107:36:@74513.4]
  assign RetimeWrapper_2_clock = clock; // @[:@74499.4]
  assign RetimeWrapper_2_reset = reset; // @[:@74500.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@74502.4]
  assign RetimeWrapper_2_io_in = x701_ctrchain_io_output_done; // @[package.scala 94:16:@74501.4]
  assign RetimeWrapper_3_clock = clock; // @[:@74539.4]
  assign RetimeWrapper_3_reset = reset; // @[:@74540.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@74542.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@74541.4]
  assign RetimeWrapper_4_clock = clock; // @[:@74547.4]
  assign RetimeWrapper_4_reset = reset; // @[:@74548.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@74550.4]
  assign RetimeWrapper_4_io_in = x717_inr_Foreach_sm_io_done; // @[package.scala 94:16:@74549.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_clock = clock; // @[:@74581.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_reset = reset; // @[:@74582.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x677_reg_rPort_0_output_0 = x677_reg_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@74655.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x670_ready = io_in_x670_ready; // @[sm_x717_inr_Foreach.scala 57:23:@74663.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_b674_number = io_in_b674_number; // @[sm_x717_inr_Foreach.scala 58:23:@74664.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_output_0 = io_in_x539_out_sram_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@74665.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_in_x676_reg_rPort_0_output_0 = x676_reg_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@74670.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x670_ready | x717_inr_Foreach_sm_io_doneLatch; // @[sm_x717_inr_Foreach.scala 132:22:@74689.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_472 & _T_473; // @[sm_x717_inr_Foreach.scala 132:22:@74687.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_break = x717_inr_Foreach_sm_io_break; // @[sm_x717_inr_Foreach.scala 132:22:@74685.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x701_ctrchain_io_output_counts_0; // @[sm_x717_inr_Foreach.scala 132:22:@74680.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x701_ctrchain_io_output_oobs_0; // @[sm_x717_inr_Foreach.scala 132:22:@74679.4]
  assign x717_inr_Foreach_kernelx717_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x717_inr_Foreach.scala 131:18:@74675.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_333 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_333 <= 1'h0;
    end else begin
      _T_333 <= _T_330;
    end
  end
endmodule
module x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1( // @[:@75035.2]
  output  io_in_x671_ready, // @[:@75038.4]
  input   io_sigsIn_datapathEn // @[:@75038.4]
);
  assign io_in_x671_ready = io_sigsIn_datapathEn; // @[sm_x722_inr_UnitPipe.scala 62:18:@75050.4]
endmodule
module x723_outr_Foreach_kernelx723_outr_Foreach_concrete1( // @[:@75053.2]
  input         clock, // @[:@75054.4]
  input         reset, // @[:@75055.4]
  input         io_in_x670_ready, // @[:@75056.4]
  output        io_in_x670_valid, // @[:@75056.4]
  output [31:0] io_in_x670_bits_wdata_0, // @[:@75056.4]
  output        io_in_x670_bits_wstrb, // @[:@75056.4]
  input         io_in_x669_ready, // @[:@75056.4]
  output        io_in_x669_valid, // @[:@75056.4]
  output [63:0] io_in_x669_bits_addr, // @[:@75056.4]
  output [31:0] io_in_x669_bits_size, // @[:@75056.4]
  input  [63:0] io_in_x470_out_host_number, // @[:@75056.4]
  output [8:0]  io_in_x539_out_sram_0_rPort_0_ofs_0, // @[:@75056.4]
  output        io_in_x539_out_sram_0_rPort_0_en_0, // @[:@75056.4]
  output        io_in_x539_out_sram_0_rPort_0_backpressure, // @[:@75056.4]
  input  [31:0] io_in_x539_out_sram_0_rPort_0_output_0, // @[:@75056.4]
  output        io_in_x671_ready, // @[:@75056.4]
  input         io_in_x671_valid, // @[:@75056.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@75056.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@75056.4]
  input         io_sigsIn_smChildAcks_0, // @[:@75056.4]
  input         io_sigsIn_smChildAcks_1, // @[:@75056.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@75056.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@75056.4]
  output        io_sigsOut_smDoneIn_0, // @[:@75056.4]
  output        io_sigsOut_smDoneIn_1, // @[:@75056.4]
  output        io_sigsOut_smMaskIn_0, // @[:@75056.4]
  output        io_sigsOut_smMaskIn_1, // @[:@75056.4]
  input         io_rr // @[:@75056.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@75085.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@75085.4]
  wire  x718_outr_UnitPipe_sm_clock; // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
  wire  x718_outr_UnitPipe_sm_reset; // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
  wire  x718_outr_UnitPipe_sm_io_enable; // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
  wire  x718_outr_UnitPipe_sm_io_done; // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
  wire  x718_outr_UnitPipe_sm_io_ctrDone; // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
  wire  x718_outr_UnitPipe_sm_io_ctrInc; // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
  wire  x718_outr_UnitPipe_sm_io_ctrRst; // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
  wire  x718_outr_UnitPipe_sm_io_parentAck; // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
  wire  x718_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
  wire  x718_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
  wire  x718_outr_UnitPipe_sm_io_maskIn_0; // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
  wire  x718_outr_UnitPipe_sm_io_maskIn_1; // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
  wire  x718_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
  wire  x718_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
  wire  x718_outr_UnitPipe_sm_io_childAck_0; // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
  wire  x718_outr_UnitPipe_sm_io_childAck_1; // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@75203.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@75203.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@75203.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@75203.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@75203.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@75211.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@75211.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@75211.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@75211.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@75211.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_clock; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_reset; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_ready; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_valid; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire [31:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_bits_wdata_0; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_bits_wstrb; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_ready; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_valid; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire [63:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_bits_addr; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire [31:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_bits_size; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire [31:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_b674_number; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire [63:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x470_out_host_number; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire [8:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_en_0; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire [31:0] x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_output_0; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smMaskIn_1; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_rr; // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
  wire  x722_inr_UnitPipe_sm_clock; // @[sm_x722_inr_UnitPipe.scala 33:18:@75384.4]
  wire  x722_inr_UnitPipe_sm_reset; // @[sm_x722_inr_UnitPipe.scala 33:18:@75384.4]
  wire  x722_inr_UnitPipe_sm_io_enable; // @[sm_x722_inr_UnitPipe.scala 33:18:@75384.4]
  wire  x722_inr_UnitPipe_sm_io_done; // @[sm_x722_inr_UnitPipe.scala 33:18:@75384.4]
  wire  x722_inr_UnitPipe_sm_io_doneLatch; // @[sm_x722_inr_UnitPipe.scala 33:18:@75384.4]
  wire  x722_inr_UnitPipe_sm_io_ctrDone; // @[sm_x722_inr_UnitPipe.scala 33:18:@75384.4]
  wire  x722_inr_UnitPipe_sm_io_datapathEn; // @[sm_x722_inr_UnitPipe.scala 33:18:@75384.4]
  wire  x722_inr_UnitPipe_sm_io_ctrInc; // @[sm_x722_inr_UnitPipe.scala 33:18:@75384.4]
  wire  x722_inr_UnitPipe_sm_io_parentAck; // @[sm_x722_inr_UnitPipe.scala 33:18:@75384.4]
  wire  x722_inr_UnitPipe_sm_io_backpressure; // @[sm_x722_inr_UnitPipe.scala 33:18:@75384.4]
  wire  x722_inr_UnitPipe_sm_io_break; // @[sm_x722_inr_UnitPipe.scala 33:18:@75384.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@75442.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@75442.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@75442.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@75442.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@75442.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@75450.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@75450.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@75450.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@75450.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@75450.4]
  wire  x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_x671_ready; // @[sm_x722_inr_UnitPipe.scala 65:24:@75479.4]
  wire  x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x722_inr_UnitPipe.scala 65:24:@75479.4]
  wire  b675; // @[sm_x723_outr_Foreach.scala 77:18:@75093.4]
  wire  _T_342; // @[package.scala 100:49:@75168.4]
  reg  _T_345; // @[package.scala 48:56:@75169.4]
  reg [31:0] _RAND_0;
  wire  _T_360; // @[package.scala 96:25:@75208.4 package.scala 96:25:@75209.4]
  wire  _T_366; // @[package.scala 96:25:@75216.4 package.scala 96:25:@75217.4]
  wire  _T_369; // @[SpatialBlocks.scala 137:99:@75219.4]
  wire  _T_437; // @[package.scala 100:49:@75412.4]
  reg  _T_440; // @[package.scala 48:56:@75413.4]
  reg [31:0] _RAND_1;
  wire  x722_inr_UnitPipe_mySignalsIn_forwardpressure; // @[sm_x723_outr_Foreach.scala 90:69:@75420.4]
  wire  _T_454; // @[package.scala 96:25:@75447.4 package.scala 96:25:@75448.4]
  wire  _T_460; // @[package.scala 96:25:@75455.4 package.scala 96:25:@75456.4]
  wire  _T_463; // @[SpatialBlocks.scala 137:99:@75458.4]
  wire  x722_inr_UnitPipe_mySignalsIn_baseEn; // @[SpatialBlocks.scala 137:96:@75459.4]
  _ _ ( // @[Math.scala 720:24:@75085.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  x537_outr_Foreach_sm x718_outr_UnitPipe_sm ( // @[sm_x718_outr_UnitPipe.scala 36:18:@75135.4]
    .clock(x718_outr_UnitPipe_sm_clock),
    .reset(x718_outr_UnitPipe_sm_reset),
    .io_enable(x718_outr_UnitPipe_sm_io_enable),
    .io_done(x718_outr_UnitPipe_sm_io_done),
    .io_ctrDone(x718_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x718_outr_UnitPipe_sm_io_ctrInc),
    .io_ctrRst(x718_outr_UnitPipe_sm_io_ctrRst),
    .io_parentAck(x718_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x718_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x718_outr_UnitPipe_sm_io_doneIn_1),
    .io_maskIn_0(x718_outr_UnitPipe_sm_io_maskIn_0),
    .io_maskIn_1(x718_outr_UnitPipe_sm_io_maskIn_1),
    .io_enableOut_0(x718_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x718_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x718_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x718_outr_UnitPipe_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@75203.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@75211.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1 x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1 ( // @[sm_x718_outr_UnitPipe.scala 112:24:@75240.4]
    .clock(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_clock),
    .reset(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_reset),
    .io_in_x670_ready(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_ready),
    .io_in_x670_valid(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_valid),
    .io_in_x670_bits_wdata_0(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_bits_wdata_0),
    .io_in_x670_bits_wstrb(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_bits_wstrb),
    .io_in_x669_ready(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_ready),
    .io_in_x669_valid(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_valid),
    .io_in_x669_bits_addr(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_bits_addr),
    .io_in_x669_bits_size(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_bits_size),
    .io_in_b674_number(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_b674_number),
    .io_in_x470_out_host_number(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x470_out_host_number),
    .io_in_x539_out_sram_0_rPort_0_ofs_0(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0),
    .io_in_x539_out_sram_0_rPort_0_en_0(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_en_0),
    .io_in_x539_out_sram_0_rPort_0_backpressure(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure),
    .io_in_x539_out_sram_0_rPort_0_output_0(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_output_0),
    .io_sigsIn_smEnableOuts_0(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smMaskIn_1(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smMaskIn_1),
    .io_rr(x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_rr)
  );
  x516_inr_UnitPipe_sm x722_inr_UnitPipe_sm ( // @[sm_x722_inr_UnitPipe.scala 33:18:@75384.4]
    .clock(x722_inr_UnitPipe_sm_clock),
    .reset(x722_inr_UnitPipe_sm_reset),
    .io_enable(x722_inr_UnitPipe_sm_io_enable),
    .io_done(x722_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x722_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x722_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x722_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x722_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x722_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x722_inr_UnitPipe_sm_io_backpressure),
    .io_break(x722_inr_UnitPipe_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@75442.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@75450.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1 x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1 ( // @[sm_x722_inr_UnitPipe.scala 65:24:@75479.4]
    .io_in_x671_ready(x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_x671_ready),
    .io_sigsIn_datapathEn(x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign b675 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x723_outr_Foreach.scala 77:18:@75093.4]
  assign _T_342 = x718_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@75168.4]
  assign _T_360 = RetimeWrapper_io_out; // @[package.scala 96:25:@75208.4 package.scala 96:25:@75209.4]
  assign _T_366 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@75216.4 package.scala 96:25:@75217.4]
  assign _T_369 = ~ _T_366; // @[SpatialBlocks.scala 137:99:@75219.4]
  assign _T_437 = x722_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@75412.4]
  assign x722_inr_UnitPipe_mySignalsIn_forwardpressure = io_in_x671_valid | x722_inr_UnitPipe_sm_io_doneLatch; // @[sm_x723_outr_Foreach.scala 90:69:@75420.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@75447.4 package.scala 96:25:@75448.4]
  assign _T_460 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@75455.4 package.scala 96:25:@75456.4]
  assign _T_463 = ~ _T_460; // @[SpatialBlocks.scala 137:99:@75458.4]
  assign x722_inr_UnitPipe_mySignalsIn_baseEn = _T_454 & _T_463; // @[SpatialBlocks.scala 137:96:@75459.4]
  assign io_in_x670_valid = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_valid; // @[sm_x718_outr_UnitPipe.scala 60:23:@75302.4]
  assign io_in_x670_bits_wdata_0 = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_bits_wdata_0; // @[sm_x718_outr_UnitPipe.scala 60:23:@75301.4]
  assign io_in_x670_bits_wstrb = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_bits_wstrb; // @[sm_x718_outr_UnitPipe.scala 60:23:@75300.4]
  assign io_in_x669_valid = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_valid; // @[sm_x718_outr_UnitPipe.scala 61:23:@75306.4]
  assign io_in_x669_bits_addr = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_bits_addr; // @[sm_x718_outr_UnitPipe.scala 61:23:@75305.4]
  assign io_in_x669_bits_size = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_bits_size; // @[sm_x718_outr_UnitPipe.scala 61:23:@75304.4]
  assign io_in_x539_out_sram_0_rPort_0_ofs_0 = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@75314.4]
  assign io_in_x539_out_sram_0_rPort_0_en_0 = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@75313.4]
  assign io_in_x539_out_sram_0_rPort_0_backpressure = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@75312.4]
  assign io_in_x671_ready = x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_in_x671_ready; // @[sm_x722_inr_UnitPipe.scala 50:23:@75517.4]
  assign io_sigsOut_smDoneIn_0 = x718_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 155:56:@75226.4]
  assign io_sigsOut_smDoneIn_1 = x722_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 155:56:@75465.4]
  assign io_sigsOut_smMaskIn_0 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[SpatialBlocks.scala 155:86:@75227.4]
  assign io_sigsOut_smMaskIn_1 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[SpatialBlocks.scala 155:86:@75466.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@75088.4]
  assign x718_outr_UnitPipe_sm_clock = clock; // @[:@75136.4]
  assign x718_outr_UnitPipe_sm_reset = reset; // @[:@75137.4]
  assign x718_outr_UnitPipe_sm_io_enable = _T_360 & _T_369; // @[SpatialBlocks.scala 139:18:@75223.4]
  assign x718_outr_UnitPipe_sm_io_ctrDone = x718_outr_UnitPipe_sm_io_ctrInc & _T_345; // @[sm_x723_outr_Foreach.scala 79:40:@75172.4]
  assign x718_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@75225.4]
  assign x718_outr_UnitPipe_sm_io_doneIn_0 = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@75193.4]
  assign x718_outr_UnitPipe_sm_io_doneIn_1 = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:72:@75194.4]
  assign x718_outr_UnitPipe_sm_io_maskIn_0 = 1'h1; // @[SpatialBlocks.scala 131:72:@75195.4]
  assign x718_outr_UnitPipe_sm_io_maskIn_1 = x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsOut_smMaskIn_1; // @[SpatialBlocks.scala 131:72:@75196.4]
  assign RetimeWrapper_clock = clock; // @[:@75204.4]
  assign RetimeWrapper_reset = reset; // @[:@75205.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@75207.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@75206.4]
  assign RetimeWrapper_1_clock = clock; // @[:@75212.4]
  assign RetimeWrapper_1_reset = reset; // @[:@75213.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@75215.4]
  assign RetimeWrapper_1_io_in = x718_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@75214.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_clock = clock; // @[:@75241.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_reset = reset; // @[:@75242.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x670_ready = io_in_x670_ready; // @[sm_x718_outr_UnitPipe.scala 60:23:@75303.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x669_ready = io_in_x669_ready; // @[sm_x718_outr_UnitPipe.scala 61:23:@75307.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_b674_number = __io_result; // @[sm_x718_outr_UnitPipe.scala 62:23:@75308.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x470_out_host_number = io_in_x470_out_host_number; // @[sm_x718_outr_UnitPipe.scala 64:32:@75310.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_in_x539_out_sram_0_rPort_0_output_0 = io_in_x539_out_sram_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@75311.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x718_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x718_outr_UnitPipe.scala 117:22:@75326.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x718_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x718_outr_UnitPipe.scala 117:22:@75327.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x718_outr_UnitPipe_sm_io_childAck_0; // @[sm_x718_outr_UnitPipe.scala 117:22:@75322.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x718_outr_UnitPipe_sm_io_childAck_1; // @[sm_x718_outr_UnitPipe.scala 117:22:@75323.4]
  assign x718_outr_UnitPipe_kernelx718_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x718_outr_UnitPipe.scala 116:18:@75316.4]
  assign x722_inr_UnitPipe_sm_clock = clock; // @[:@75385.4]
  assign x722_inr_UnitPipe_sm_reset = reset; // @[:@75386.4]
  assign x722_inr_UnitPipe_sm_io_enable = x722_inr_UnitPipe_mySignalsIn_baseEn & x722_inr_UnitPipe_mySignalsIn_forwardpressure; // @[SpatialBlocks.scala 139:18:@75462.4]
  assign x722_inr_UnitPipe_sm_io_ctrDone = x722_inr_UnitPipe_sm_io_ctrInc & _T_440; // @[sm_x723_outr_Foreach.scala 88:39:@75416.4]
  assign x722_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 141:21:@75464.4]
  assign x722_inr_UnitPipe_sm_io_backpressure = 1'h1; // @[SpatialBlocks.scala 132:24:@75436.4]
  assign x722_inr_UnitPipe_sm_io_break = 1'h0; // @[sm_x723_outr_Foreach.scala 92:37:@75423.4]
  assign RetimeWrapper_2_clock = clock; // @[:@75443.4]
  assign RetimeWrapper_2_reset = reset; // @[:@75444.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@75446.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@75445.4]
  assign RetimeWrapper_3_clock = clock; // @[:@75451.4]
  assign RetimeWrapper_3_reset = reset; // @[:@75452.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@75454.4]
  assign RetimeWrapper_3_io_in = x722_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@75453.4]
  assign x722_inr_UnitPipe_kernelx722_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x722_inr_UnitPipe_sm_io_datapathEn & b675; // @[sm_x722_inr_UnitPipe.scala 70:22:@75530.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_345 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_440 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_345 <= 1'h0;
    end else begin
      _T_345 <= _T_342;
    end
    if (reset) begin
      _T_440 <= 1'h0;
    end else begin
      _T_440 <= _T_437;
    end
  end
endmodule
module x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1( // @[:@75546.2]
  input         clock, // @[:@75547.4]
  input         reset, // @[:@75548.4]
  input         io_in_x670_ready, // @[:@75549.4]
  output        io_in_x670_valid, // @[:@75549.4]
  output [31:0] io_in_x670_bits_wdata_0, // @[:@75549.4]
  output        io_in_x670_bits_wstrb, // @[:@75549.4]
  input         io_in_x669_ready, // @[:@75549.4]
  output        io_in_x669_valid, // @[:@75549.4]
  output [63:0] io_in_x669_bits_addr, // @[:@75549.4]
  output [31:0] io_in_x669_bits_size, // @[:@75549.4]
  input  [63:0] io_in_x470_out_host_number, // @[:@75549.4]
  output [8:0]  io_in_x539_out_sram_0_rPort_0_ofs_0, // @[:@75549.4]
  output        io_in_x539_out_sram_0_rPort_0_en_0, // @[:@75549.4]
  output        io_in_x539_out_sram_0_rPort_0_backpressure, // @[:@75549.4]
  input  [31:0] io_in_x539_out_sram_0_rPort_0_output_0, // @[:@75549.4]
  output        io_in_x671_ready, // @[:@75549.4]
  input         io_in_x671_valid, // @[:@75549.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@75549.4]
  input         io_sigsIn_smChildAcks_0, // @[:@75549.4]
  output        io_sigsOut_smDoneIn_0, // @[:@75549.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@75549.4]
  input         io_rr // @[:@75549.4]
);
  wire  x673_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@75572.4]
  wire  x673_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@75572.4]
  wire  x673_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@75572.4]
  wire  x673_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@75572.4]
  wire [8:0] x673_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@75572.4]
  wire  x673_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@75572.4]
  wire  x673_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@75572.4]
  wire  x723_outr_Foreach_sm_clock; // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
  wire  x723_outr_Foreach_sm_reset; // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
  wire  x723_outr_Foreach_sm_io_enable; // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
  wire  x723_outr_Foreach_sm_io_done; // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
  wire  x723_outr_Foreach_sm_io_ctrDone; // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
  wire  x723_outr_Foreach_sm_io_ctrInc; // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
  wire  x723_outr_Foreach_sm_io_ctrRst; // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
  wire  x723_outr_Foreach_sm_io_parentAck; // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
  wire  x723_outr_Foreach_sm_io_doneIn_0; // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
  wire  x723_outr_Foreach_sm_io_doneIn_1; // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
  wire  x723_outr_Foreach_sm_io_maskIn_0; // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
  wire  x723_outr_Foreach_sm_io_maskIn_1; // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
  wire  x723_outr_Foreach_sm_io_enableOut_0; // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
  wire  x723_outr_Foreach_sm_io_enableOut_1; // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
  wire  x723_outr_Foreach_sm_io_childAck_0; // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
  wire  x723_outr_Foreach_sm_io_childAck_1; // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@75664.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@75664.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@75664.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@75664.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@75664.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@75709.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@75709.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@75709.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@75709.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@75709.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@75717.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@75717.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@75717.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@75717.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@75717.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_clock; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_reset; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_ready; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_valid; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire [31:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_bits_wdata_0; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_bits_wstrb; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_ready; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_valid; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_bits_addr; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire [31:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_bits_size; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire [63:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x470_out_host_number; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire [8:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_en_0; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire [31:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_output_0; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x671_ready; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x671_valid; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire [31:0] x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_rr; // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
  wire  _T_339; // @[package.scala 96:25:@75669.4 package.scala 96:25:@75670.4]
  wire  _T_356; // @[package.scala 96:25:@75714.4 package.scala 96:25:@75715.4]
  wire  _T_362; // @[package.scala 96:25:@75722.4 package.scala 96:25:@75723.4]
  wire  _T_365; // @[SpatialBlocks.scala 137:99:@75725.4]
  x478_ctrchain x673_ctrchain ( // @[SpatialBlocks.scala 37:22:@75572.4]
    .clock(x673_ctrchain_clock),
    .reset(x673_ctrchain_reset),
    .io_input_reset(x673_ctrchain_io_input_reset),
    .io_input_enable(x673_ctrchain_io_input_enable),
    .io_output_counts_0(x673_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x673_ctrchain_io_output_oobs_0),
    .io_output_done(x673_ctrchain_io_output_done)
  );
  x537_outr_Foreach_sm x723_outr_Foreach_sm ( // @[sm_x723_outr_Foreach.scala 36:18:@75630.4]
    .clock(x723_outr_Foreach_sm_clock),
    .reset(x723_outr_Foreach_sm_reset),
    .io_enable(x723_outr_Foreach_sm_io_enable),
    .io_done(x723_outr_Foreach_sm_io_done),
    .io_ctrDone(x723_outr_Foreach_sm_io_ctrDone),
    .io_ctrInc(x723_outr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x723_outr_Foreach_sm_io_ctrRst),
    .io_parentAck(x723_outr_Foreach_sm_io_parentAck),
    .io_doneIn_0(x723_outr_Foreach_sm_io_doneIn_0),
    .io_doneIn_1(x723_outr_Foreach_sm_io_doneIn_1),
    .io_maskIn_0(x723_outr_Foreach_sm_io_maskIn_0),
    .io_maskIn_1(x723_outr_Foreach_sm_io_maskIn_1),
    .io_enableOut_0(x723_outr_Foreach_sm_io_enableOut_0),
    .io_enableOut_1(x723_outr_Foreach_sm_io_enableOut_1),
    .io_childAck_0(x723_outr_Foreach_sm_io_childAck_0),
    .io_childAck_1(x723_outr_Foreach_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@75664.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@75709.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@75717.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x723_outr_Foreach_kernelx723_outr_Foreach_concrete1 x723_outr_Foreach_kernelx723_outr_Foreach_concrete1 ( // @[sm_x723_outr_Foreach.scala 97:24:@75752.4]
    .clock(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_clock),
    .reset(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_reset),
    .io_in_x670_ready(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_ready),
    .io_in_x670_valid(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_valid),
    .io_in_x670_bits_wdata_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_bits_wdata_0),
    .io_in_x670_bits_wstrb(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_bits_wstrb),
    .io_in_x669_ready(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_ready),
    .io_in_x669_valid(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_valid),
    .io_in_x669_bits_addr(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_bits_addr),
    .io_in_x669_bits_size(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_bits_size),
    .io_in_x470_out_host_number(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x470_out_host_number),
    .io_in_x539_out_sram_0_rPort_0_ofs_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0),
    .io_in_x539_out_sram_0_rPort_0_en_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_en_0),
    .io_in_x539_out_sram_0_rPort_0_backpressure(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure),
    .io_in_x539_out_sram_0_rPort_0_output_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_output_0),
    .io_in_x671_ready(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x671_ready),
    .io_in_x671_valid(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x671_valid),
    .io_sigsIn_smEnableOuts_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsOut_smDoneIn_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smMaskIn_0(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0),
    .io_sigsOut_smMaskIn_1(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1),
    .io_rr(x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_rr)
  );
  assign _T_339 = RetimeWrapper_io_out; // @[package.scala 96:25:@75669.4 package.scala 96:25:@75670.4]
  assign _T_356 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@75714.4 package.scala 96:25:@75715.4]
  assign _T_362 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@75722.4 package.scala 96:25:@75723.4]
  assign _T_365 = ~ _T_362; // @[SpatialBlocks.scala 137:99:@75725.4]
  assign io_in_x670_valid = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_valid; // @[sm_x723_outr_Foreach.scala 58:23:@75815.4]
  assign io_in_x670_bits_wdata_0 = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_bits_wdata_0; // @[sm_x723_outr_Foreach.scala 58:23:@75814.4]
  assign io_in_x670_bits_wstrb = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_bits_wstrb; // @[sm_x723_outr_Foreach.scala 58:23:@75813.4]
  assign io_in_x669_valid = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_valid; // @[sm_x723_outr_Foreach.scala 59:23:@75819.4]
  assign io_in_x669_bits_addr = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_bits_addr; // @[sm_x723_outr_Foreach.scala 59:23:@75818.4]
  assign io_in_x669_bits_size = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_bits_size; // @[sm_x723_outr_Foreach.scala 59:23:@75817.4]
  assign io_in_x539_out_sram_0_rPort_0_ofs_0 = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@75825.4]
  assign io_in_x539_out_sram_0_rPort_0_en_0 = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@75824.4]
  assign io_in_x539_out_sram_0_rPort_0_backpressure = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@75823.4]
  assign io_in_x671_ready = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x671_ready; // @[sm_x723_outr_Foreach.scala 62:23:@75829.4]
  assign io_sigsOut_smDoneIn_0 = x723_outr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@75732.4]
  assign io_sigsOut_smCtrCopyDone_0 = x723_outr_Foreach_sm_io_done; // @[SpatialBlocks.scala 170:140:@75751.4]
  assign x673_ctrchain_clock = clock; // @[:@75573.4]
  assign x673_ctrchain_reset = reset; // @[:@75574.4]
  assign x673_ctrchain_io_input_reset = x723_outr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@75750.4]
  assign x673_ctrchain_io_input_enable = x723_outr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 158:42:@75749.4]
  assign x723_outr_Foreach_sm_clock = clock; // @[:@75631.4]
  assign x723_outr_Foreach_sm_reset = reset; // @[:@75632.4]
  assign x723_outr_Foreach_sm_io_enable = _T_356 & _T_365; // @[SpatialBlocks.scala 139:18:@75729.4]
  assign x723_outr_Foreach_sm_io_ctrDone = io_rr ? _T_339 : 1'h0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 81:39:@75672.4]
  assign x723_outr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@75731.4]
  assign x723_outr_Foreach_sm_io_doneIn_0 = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@75699.4]
  assign x723_outr_Foreach_sm_io_doneIn_1 = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:72:@75700.4]
  assign x723_outr_Foreach_sm_io_maskIn_0 = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0; // @[SpatialBlocks.scala 131:72:@75701.4]
  assign x723_outr_Foreach_sm_io_maskIn_1 = x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1; // @[SpatialBlocks.scala 131:72:@75702.4]
  assign RetimeWrapper_clock = clock; // @[:@75665.4]
  assign RetimeWrapper_reset = reset; // @[:@75666.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@75668.4]
  assign RetimeWrapper_io_in = x673_ctrchain_io_output_done; // @[package.scala 94:16:@75667.4]
  assign RetimeWrapper_1_clock = clock; // @[:@75710.4]
  assign RetimeWrapper_1_reset = reset; // @[:@75711.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@75713.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@75712.4]
  assign RetimeWrapper_2_clock = clock; // @[:@75718.4]
  assign RetimeWrapper_2_reset = reset; // @[:@75719.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@75721.4]
  assign RetimeWrapper_2_io_in = x723_outr_Foreach_sm_io_done; // @[package.scala 94:16:@75720.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_clock = clock; // @[:@75753.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_reset = reset; // @[:@75754.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x670_ready = io_in_x670_ready; // @[sm_x723_outr_Foreach.scala 58:23:@75816.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x669_ready = io_in_x669_ready; // @[sm_x723_outr_Foreach.scala 59:23:@75820.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x470_out_host_number = io_in_x470_out_host_number; // @[sm_x723_outr_Foreach.scala 60:32:@75821.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x539_out_sram_0_rPort_0_output_0 = io_in_x539_out_sram_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@75822.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_in_x671_valid = io_in_x671_valid; // @[sm_x723_outr_Foreach.scala 62:23:@75828.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0 = x723_outr_Foreach_sm_io_enableOut_0; // @[sm_x723_outr_Foreach.scala 102:22:@75840.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1 = x723_outr_Foreach_sm_io_enableOut_1; // @[sm_x723_outr_Foreach.scala 102:22:@75841.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0 = x723_outr_Foreach_sm_io_childAck_0; // @[sm_x723_outr_Foreach.scala 102:22:@75836.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1 = x723_outr_Foreach_sm_io_childAck_1; // @[sm_x723_outr_Foreach.scala 102:22:@75837.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{23{x673_ctrchain_io_output_counts_0[8]}},x673_ctrchain_io_output_counts_0}; // @[sm_x723_outr_Foreach.scala 102:22:@75835.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x673_ctrchain_io_output_oobs_0; // @[sm_x723_outr_Foreach.scala 102:22:@75834.4]
  assign x723_outr_Foreach_kernelx723_outr_Foreach_concrete1_io_rr = io_rr; // @[sm_x723_outr_Foreach.scala 101:18:@75830.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@75863.2]
  input         clock, // @[:@75864.4]
  input         reset, // @[:@75865.4]
  input  [63:0] io_in_x468_A_dram_number, // @[:@75866.4]
  input         io_in_x670_ready, // @[:@75866.4]
  output        io_in_x670_valid, // @[:@75866.4]
  output [31:0] io_in_x670_bits_wdata_0, // @[:@75866.4]
  output        io_in_x670_bits_wstrb, // @[:@75866.4]
  input         io_in_x669_ready, // @[:@75866.4]
  output        io_in_x669_valid, // @[:@75866.4]
  output [63:0] io_in_x669_bits_addr, // @[:@75866.4]
  output [31:0] io_in_x669_bits_size, // @[:@75866.4]
  output        io_in_x476_ready, // @[:@75866.4]
  input         io_in_x476_valid, // @[:@75866.4]
  input  [31:0] io_in_x476_bits_rdata_0, // @[:@75866.4]
  input  [63:0] io_in_x470_out_host_number, // @[:@75866.4]
  output        io_in_x671_ready, // @[:@75866.4]
  input         io_in_x671_valid, // @[:@75866.4]
  input         io_in_x474_ready, // @[:@75866.4]
  output        io_in_x474_valid, // @[:@75866.4]
  output [63:0] io_in_x474_bits_addr, // @[:@75866.4]
  output [31:0] io_in_x474_bits_size, // @[:@75866.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@75866.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@75866.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@75866.4]
  input         io_sigsIn_smChildAcks_0, // @[:@75866.4]
  input         io_sigsIn_smChildAcks_1, // @[:@75866.4]
  input         io_sigsIn_smChildAcks_2, // @[:@75866.4]
  output        io_sigsOut_smDoneIn_0, // @[:@75866.4]
  output        io_sigsOut_smDoneIn_1, // @[:@75866.4]
  output        io_sigsOut_smDoneIn_2, // @[:@75866.4]
  input         io_rr // @[:@75866.4]
);
  wire  x471_A_sram_0_clock; // @[m_x471_A_sram_0.scala 27:22:@75880.4]
  wire  x471_A_sram_0_reset; // @[m_x471_A_sram_0.scala 27:22:@75880.4]
  wire [8:0] x471_A_sram_0_io_rPort_0_ofs_0; // @[m_x471_A_sram_0.scala 27:22:@75880.4]
  wire  x471_A_sram_0_io_rPort_0_en_0; // @[m_x471_A_sram_0.scala 27:22:@75880.4]
  wire  x471_A_sram_0_io_rPort_0_backpressure; // @[m_x471_A_sram_0.scala 27:22:@75880.4]
  wire [31:0] x471_A_sram_0_io_rPort_0_output_0; // @[m_x471_A_sram_0.scala 27:22:@75880.4]
  wire [8:0] x471_A_sram_0_io_wPort_0_ofs_0; // @[m_x471_A_sram_0.scala 27:22:@75880.4]
  wire [31:0] x471_A_sram_0_io_wPort_0_data_0; // @[m_x471_A_sram_0.scala 27:22:@75880.4]
  wire  x471_A_sram_0_io_wPort_0_en_0; // @[m_x471_A_sram_0.scala 27:22:@75880.4]
  wire  x472_A_sram_1_clock; // @[m_x472_A_sram_1.scala 27:22:@75897.4]
  wire  x472_A_sram_1_reset; // @[m_x472_A_sram_1.scala 27:22:@75897.4]
  wire [8:0] x472_A_sram_1_io_rPort_0_ofs_0; // @[m_x472_A_sram_1.scala 27:22:@75897.4]
  wire  x472_A_sram_1_io_rPort_0_en_0; // @[m_x472_A_sram_1.scala 27:22:@75897.4]
  wire  x472_A_sram_1_io_rPort_0_backpressure; // @[m_x472_A_sram_1.scala 27:22:@75897.4]
  wire [31:0] x472_A_sram_1_io_rPort_0_output_0; // @[m_x472_A_sram_1.scala 27:22:@75897.4]
  wire [8:0] x472_A_sram_1_io_wPort_0_ofs_0; // @[m_x472_A_sram_1.scala 27:22:@75897.4]
  wire [31:0] x472_A_sram_1_io_wPort_0_data_0; // @[m_x472_A_sram_1.scala 27:22:@75897.4]
  wire  x472_A_sram_1_io_wPort_0_en_0; // @[m_x472_A_sram_1.scala 27:22:@75897.4]
  wire  x473_A_sram_2_clock; // @[m_x473_A_sram_2.scala 27:22:@75914.4]
  wire  x473_A_sram_2_reset; // @[m_x473_A_sram_2.scala 27:22:@75914.4]
  wire [8:0] x473_A_sram_2_io_rPort_0_ofs_0; // @[m_x473_A_sram_2.scala 27:22:@75914.4]
  wire  x473_A_sram_2_io_rPort_0_en_0; // @[m_x473_A_sram_2.scala 27:22:@75914.4]
  wire  x473_A_sram_2_io_rPort_0_backpressure; // @[m_x473_A_sram_2.scala 27:22:@75914.4]
  wire [31:0] x473_A_sram_2_io_rPort_0_output_0; // @[m_x473_A_sram_2.scala 27:22:@75914.4]
  wire [8:0] x473_A_sram_2_io_wPort_0_ofs_0; // @[m_x473_A_sram_2.scala 27:22:@75914.4]
  wire [31:0] x473_A_sram_2_io_wPort_0_data_0; // @[m_x473_A_sram_2.scala 27:22:@75914.4]
  wire  x473_A_sram_2_io_wPort_0_en_0; // @[m_x473_A_sram_2.scala 27:22:@75914.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_clock; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@75979.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_reset; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@75979.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_enable; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@75979.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_done; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@75979.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_parentAck; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@75979.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_doneIn_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@75979.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_doneIn_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@75979.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_enableOut_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@75979.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_enableOut_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@75979.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_childAck_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@75979.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_childAck_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@75979.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@75979.4]
  wire  x538_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@75979.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@76042.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@76042.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@76042.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@76042.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@76042.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@76050.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@76050.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@76050.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@76050.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@76050.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_clock; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_reset; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x468_A_dram_number; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire [8:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire [31:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_data_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_en_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire [8:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire [31:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_data_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_en_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_ready; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_valid; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire [31:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_bits_rdata_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire [8:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire [31:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_data_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_en_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_ready; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_valid; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire [63:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_bits_addr; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire [31:0] x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_bits_size; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_rr; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
  wire  x539_out_sram_0_clock; // @[m_x539_out_sram_0.scala 27:22:@76239.4]
  wire  x539_out_sram_0_reset; // @[m_x539_out_sram_0.scala 27:22:@76239.4]
  wire [8:0] x539_out_sram_0_io_rPort_0_ofs_0; // @[m_x539_out_sram_0.scala 27:22:@76239.4]
  wire  x539_out_sram_0_io_rPort_0_en_0; // @[m_x539_out_sram_0.scala 27:22:@76239.4]
  wire  x539_out_sram_0_io_rPort_0_backpressure; // @[m_x539_out_sram_0.scala 27:22:@76239.4]
  wire [31:0] x539_out_sram_0_io_rPort_0_output_0; // @[m_x539_out_sram_0.scala 27:22:@76239.4]
  wire [8:0] x539_out_sram_0_io_wPort_0_ofs_0; // @[m_x539_out_sram_0.scala 27:22:@76239.4]
  wire [31:0] x539_out_sram_0_io_wPort_0_data_0; // @[m_x539_out_sram_0.scala 27:22:@76239.4]
  wire  x539_out_sram_0_io_wPort_0_en_0; // @[m_x539_out_sram_0.scala 27:22:@76239.4]
  wire  x541_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@76256.4]
  wire  x541_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@76256.4]
  wire  x541_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@76256.4]
  wire  x541_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@76256.4]
  wire [8:0] x541_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@76256.4]
  wire  x541_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@76256.4]
  wire  x541_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@76256.4]
  wire  x668_outr_Foreach_sm_clock; // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
  wire  x668_outr_Foreach_sm_reset; // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
  wire  x668_outr_Foreach_sm_io_enable; // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
  wire  x668_outr_Foreach_sm_io_done; // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
  wire  x668_outr_Foreach_sm_io_ctrDone; // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
  wire  x668_outr_Foreach_sm_io_ctrInc; // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
  wire  x668_outr_Foreach_sm_io_ctrRst; // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
  wire  x668_outr_Foreach_sm_io_parentAck; // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
  wire  x668_outr_Foreach_sm_io_doneIn_0; // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
  wire  x668_outr_Foreach_sm_io_doneIn_1; // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
  wire  x668_outr_Foreach_sm_io_maskIn_0; // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
  wire  x668_outr_Foreach_sm_io_maskIn_1; // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
  wire  x668_outr_Foreach_sm_io_enableOut_0; // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
  wire  x668_outr_Foreach_sm_io_enableOut_1; // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
  wire  x668_outr_Foreach_sm_io_childAck_0; // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
  wire  x668_outr_Foreach_sm_io_childAck_1; // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@76348.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@76348.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@76348.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@76348.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@76348.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@76393.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@76393.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@76393.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@76393.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@76393.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@76401.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@76401.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@76401.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@76401.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@76401.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_clock; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_reset; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire [8:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_en_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire [31:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_output_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire [8:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_en_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire [31:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_output_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire [8:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_ofs_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_en_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire [31:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_output_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire [8:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_ofs_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire [31:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_data_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_en_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire [31:0] x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_rr; // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_clock; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@76613.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_reset; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@76613.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_io_enable; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@76613.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_io_done; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@76613.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_io_parentAck; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@76613.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_io_doneIn_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@76613.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_io_enableOut_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@76613.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_io_childAck_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@76613.4]
  wire  x724_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@76613.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@76666.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@76666.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@76666.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@76666.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@76666.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@76674.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@76674.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@76674.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@76674.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@76674.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_clock; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_reset; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_ready; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_valid; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire [31:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_bits_wdata_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_bits_wstrb; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_ready; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_valid; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_bits_addr; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire [31:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_bits_size; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire [63:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x470_out_host_number; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire [8:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_en_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire [31:0] x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_output_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x671_ready; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x671_valid; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_rr; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
  wire  _T_263; // @[package.scala 96:25:@76047.4 package.scala 96:25:@76048.4]
  wire  _T_269; // @[package.scala 96:25:@76055.4 package.scala 96:25:@76056.4]
  wire  _T_272; // @[SpatialBlocks.scala 137:99:@76058.4]
  wire  _T_345; // @[package.scala 96:25:@76353.4 package.scala 96:25:@76354.4]
  wire  _T_362; // @[package.scala 96:25:@76398.4 package.scala 96:25:@76399.4]
  wire  _T_368; // @[package.scala 96:25:@76406.4 package.scala 96:25:@76407.4]
  wire  _T_371; // @[SpatialBlocks.scala 137:99:@76409.4]
  wire  _T_454; // @[package.scala 96:25:@76671.4 package.scala 96:25:@76672.4]
  wire  _T_460; // @[package.scala 96:25:@76679.4 package.scala 96:25:@76680.4]
  wire  _T_463; // @[SpatialBlocks.scala 137:99:@76682.4]
  x471_A_sram_0 x471_A_sram_0 ( // @[m_x471_A_sram_0.scala 27:22:@75880.4]
    .clock(x471_A_sram_0_clock),
    .reset(x471_A_sram_0_reset),
    .io_rPort_0_ofs_0(x471_A_sram_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x471_A_sram_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x471_A_sram_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x471_A_sram_0_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(x471_A_sram_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x471_A_sram_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x471_A_sram_0_io_wPort_0_en_0)
  );
  x471_A_sram_0 x472_A_sram_1 ( // @[m_x472_A_sram_1.scala 27:22:@75897.4]
    .clock(x472_A_sram_1_clock),
    .reset(x472_A_sram_1_reset),
    .io_rPort_0_ofs_0(x472_A_sram_1_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x472_A_sram_1_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x472_A_sram_1_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x472_A_sram_1_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(x472_A_sram_1_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x472_A_sram_1_io_wPort_0_data_0),
    .io_wPort_0_en_0(x472_A_sram_1_io_wPort_0_en_0)
  );
  x471_A_sram_0 x473_A_sram_2 ( // @[m_x473_A_sram_2.scala 27:22:@75914.4]
    .clock(x473_A_sram_2_clock),
    .reset(x473_A_sram_2_reset),
    .io_rPort_0_ofs_0(x473_A_sram_2_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x473_A_sram_2_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x473_A_sram_2_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x473_A_sram_2_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(x473_A_sram_2_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x473_A_sram_2_io_wPort_0_data_0),
    .io_wPort_0_en_0(x473_A_sram_2_io_wPort_0_en_0)
  );
  x538_outr_UnitPipe_DenseTransfer_sm x538_outr_UnitPipe_DenseTransfer_sm ( // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 35:18:@75979.4]
    .clock(x538_outr_UnitPipe_DenseTransfer_sm_clock),
    .reset(x538_outr_UnitPipe_DenseTransfer_sm_reset),
    .io_enable(x538_outr_UnitPipe_DenseTransfer_sm_io_enable),
    .io_done(x538_outr_UnitPipe_DenseTransfer_sm_io_done),
    .io_parentAck(x538_outr_UnitPipe_DenseTransfer_sm_io_parentAck),
    .io_doneIn_0(x538_outr_UnitPipe_DenseTransfer_sm_io_doneIn_0),
    .io_doneIn_1(x538_outr_UnitPipe_DenseTransfer_sm_io_doneIn_1),
    .io_enableOut_0(x538_outr_UnitPipe_DenseTransfer_sm_io_enableOut_0),
    .io_enableOut_1(x538_outr_UnitPipe_DenseTransfer_sm_io_enableOut_1),
    .io_childAck_0(x538_outr_UnitPipe_DenseTransfer_sm_io_childAck_0),
    .io_childAck_1(x538_outr_UnitPipe_DenseTransfer_sm_io_childAck_1),
    .io_ctrCopyDone_0(x538_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x538_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@76042.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@76050.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1 x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1 ( // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 107:24:@76081.4]
    .clock(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_clock),
    .reset(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_reset),
    .io_in_x468_A_dram_number(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x468_A_dram_number),
    .io_in_x472_A_sram_1_wPort_0_ofs_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0),
    .io_in_x472_A_sram_1_wPort_0_data_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_data_0),
    .io_in_x472_A_sram_1_wPort_0_en_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_en_0),
    .io_in_x471_A_sram_0_wPort_0_ofs_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0),
    .io_in_x471_A_sram_0_wPort_0_data_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_data_0),
    .io_in_x471_A_sram_0_wPort_0_en_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_en_0),
    .io_in_x476_ready(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_ready),
    .io_in_x476_valid(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_valid),
    .io_in_x476_bits_rdata_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_bits_rdata_0),
    .io_in_x473_A_sram_2_wPort_0_ofs_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0),
    .io_in_x473_A_sram_2_wPort_0_data_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_data_0),
    .io_in_x473_A_sram_2_wPort_0_en_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_en_0),
    .io_in_x474_ready(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_ready),
    .io_in_x474_valid(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_valid),
    .io_in_x474_bits_addr(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_bits_addr),
    .io_in_x474_bits_size(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_bits_size),
    .io_sigsIn_smEnableOuts_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_rr)
  );
  x471_A_sram_0 x539_out_sram_0 ( // @[m_x539_out_sram_0.scala 27:22:@76239.4]
    .clock(x539_out_sram_0_clock),
    .reset(x539_out_sram_0_reset),
    .io_rPort_0_ofs_0(x539_out_sram_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x539_out_sram_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x539_out_sram_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x539_out_sram_0_io_rPort_0_output_0),
    .io_wPort_0_ofs_0(x539_out_sram_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x539_out_sram_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x539_out_sram_0_io_wPort_0_en_0)
  );
  x478_ctrchain x541_ctrchain ( // @[SpatialBlocks.scala 37:22:@76256.4]
    .clock(x541_ctrchain_clock),
    .reset(x541_ctrchain_reset),
    .io_input_reset(x541_ctrchain_io_input_reset),
    .io_input_enable(x541_ctrchain_io_input_enable),
    .io_output_counts_0(x541_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x541_ctrchain_io_output_oobs_0),
    .io_output_done(x541_ctrchain_io_output_done)
  );
  x668_outr_Foreach_sm x668_outr_Foreach_sm ( // @[sm_x668_outr_Foreach.scala 32:18:@76314.4]
    .clock(x668_outr_Foreach_sm_clock),
    .reset(x668_outr_Foreach_sm_reset),
    .io_enable(x668_outr_Foreach_sm_io_enable),
    .io_done(x668_outr_Foreach_sm_io_done),
    .io_ctrDone(x668_outr_Foreach_sm_io_ctrDone),
    .io_ctrInc(x668_outr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x668_outr_Foreach_sm_io_ctrRst),
    .io_parentAck(x668_outr_Foreach_sm_io_parentAck),
    .io_doneIn_0(x668_outr_Foreach_sm_io_doneIn_0),
    .io_doneIn_1(x668_outr_Foreach_sm_io_doneIn_1),
    .io_maskIn_0(x668_outr_Foreach_sm_io_maskIn_0),
    .io_maskIn_1(x668_outr_Foreach_sm_io_maskIn_1),
    .io_enableOut_0(x668_outr_Foreach_sm_io_enableOut_0),
    .io_enableOut_1(x668_outr_Foreach_sm_io_enableOut_1),
    .io_childAck_0(x668_outr_Foreach_sm_io_childAck_0),
    .io_childAck_1(x668_outr_Foreach_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@76348.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@76393.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@76401.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x668_outr_Foreach_kernelx668_outr_Foreach_concrete1 x668_outr_Foreach_kernelx668_outr_Foreach_concrete1 ( // @[sm_x668_outr_Foreach.scala 113:24:@76435.4]
    .clock(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_clock),
    .reset(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_reset),
    .io_in_x472_A_sram_1_rPort_0_ofs_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0),
    .io_in_x472_A_sram_1_rPort_0_en_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_en_0),
    .io_in_x472_A_sram_1_rPort_0_output_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_output_0),
    .io_in_x471_A_sram_0_rPort_0_ofs_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0),
    .io_in_x471_A_sram_0_rPort_0_en_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_en_0),
    .io_in_x471_A_sram_0_rPort_0_output_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_output_0),
    .io_in_x473_A_sram_2_rPort_0_ofs_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_ofs_0),
    .io_in_x473_A_sram_2_rPort_0_en_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_en_0),
    .io_in_x473_A_sram_2_rPort_0_output_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_output_0),
    .io_in_x539_out_sram_0_wPort_0_ofs_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_ofs_0),
    .io_in_x539_out_sram_0_wPort_0_data_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_data_0),
    .io_in_x539_out_sram_0_wPort_0_en_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_en_0),
    .io_sigsIn_smEnableOuts_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsOut_smDoneIn_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smMaskIn_0(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0),
    .io_sigsOut_smMaskIn_1(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1),
    .io_rr(x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_rr)
  );
  x724_outr_UnitPipe_DenseTransfer_sm x724_outr_UnitPipe_DenseTransfer_sm ( // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 36:18:@76613.4]
    .clock(x724_outr_UnitPipe_DenseTransfer_sm_clock),
    .reset(x724_outr_UnitPipe_DenseTransfer_sm_reset),
    .io_enable(x724_outr_UnitPipe_DenseTransfer_sm_io_enable),
    .io_done(x724_outr_UnitPipe_DenseTransfer_sm_io_done),
    .io_parentAck(x724_outr_UnitPipe_DenseTransfer_sm_io_parentAck),
    .io_doneIn_0(x724_outr_UnitPipe_DenseTransfer_sm_io_doneIn_0),
    .io_enableOut_0(x724_outr_UnitPipe_DenseTransfer_sm_io_enableOut_0),
    .io_childAck_0(x724_outr_UnitPipe_DenseTransfer_sm_io_childAck_0),
    .io_ctrCopyDone_0(x724_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@76666.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@76674.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1 x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1 ( // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 90:24:@76704.4]
    .clock(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_clock),
    .reset(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_reset),
    .io_in_x670_ready(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_ready),
    .io_in_x670_valid(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_valid),
    .io_in_x670_bits_wdata_0(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_bits_wdata_0),
    .io_in_x670_bits_wstrb(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_bits_wstrb),
    .io_in_x669_ready(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_ready),
    .io_in_x669_valid(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_valid),
    .io_in_x669_bits_addr(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_bits_addr),
    .io_in_x669_bits_size(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_bits_size),
    .io_in_x470_out_host_number(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x470_out_host_number),
    .io_in_x539_out_sram_0_rPort_0_ofs_0(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0),
    .io_in_x539_out_sram_0_rPort_0_en_0(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_en_0),
    .io_in_x539_out_sram_0_rPort_0_backpressure(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure),
    .io_in_x539_out_sram_0_rPort_0_output_0(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_output_0),
    .io_in_x671_ready(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x671_ready),
    .io_in_x671_valid(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x671_valid),
    .io_sigsIn_smEnableOuts_0(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_rr)
  );
  assign _T_263 = RetimeWrapper_io_out; // @[package.scala 96:25:@76047.4 package.scala 96:25:@76048.4]
  assign _T_269 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@76055.4 package.scala 96:25:@76056.4]
  assign _T_272 = ~ _T_269; // @[SpatialBlocks.scala 137:99:@76058.4]
  assign _T_345 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@76353.4 package.scala 96:25:@76354.4]
  assign _T_362 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@76398.4 package.scala 96:25:@76399.4]
  assign _T_368 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@76406.4 package.scala 96:25:@76407.4]
  assign _T_371 = ~ _T_368; // @[SpatialBlocks.scala 137:99:@76409.4]
  assign _T_454 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@76671.4 package.scala 96:25:@76672.4]
  assign _T_460 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@76679.4 package.scala 96:25:@76680.4]
  assign _T_463 = ~ _T_460; // @[SpatialBlocks.scala 137:99:@76682.4]
  assign io_in_x670_valid = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_valid; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 58:23:@76762.4]
  assign io_in_x670_bits_wdata_0 = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_bits_wdata_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 58:23:@76761.4]
  assign io_in_x670_bits_wstrb = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_bits_wstrb; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 58:23:@76760.4]
  assign io_in_x669_valid = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_valid; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 59:23:@76766.4]
  assign io_in_x669_bits_addr = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_bits_addr; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 59:23:@76765.4]
  assign io_in_x669_bits_size = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_bits_size; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 59:23:@76764.4]
  assign io_in_x476_ready = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_ready; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 62:23:@76188.4]
  assign io_in_x671_ready = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x671_ready; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 62:23:@76776.4]
  assign io_in_x474_valid = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_valid; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 64:23:@76198.4]
  assign io_in_x474_bits_addr = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_bits_addr; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 64:23:@76197.4]
  assign io_in_x474_bits_size = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_bits_size; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 64:23:@76196.4]
  assign io_sigsOut_smDoneIn_0 = x538_outr_UnitPipe_DenseTransfer_sm_io_done; // @[SpatialBlocks.scala 155:56:@76065.4]
  assign io_sigsOut_smDoneIn_1 = x668_outr_Foreach_sm_io_done; // @[SpatialBlocks.scala 155:56:@76416.4]
  assign io_sigsOut_smDoneIn_2 = x724_outr_UnitPipe_DenseTransfer_sm_io_done; // @[SpatialBlocks.scala 155:56:@76689.4]
  assign x471_A_sram_0_clock = clock; // @[:@75881.4]
  assign x471_A_sram_0_reset = reset; // @[:@75882.4]
  assign x471_A_sram_0_io_rPort_0_ofs_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@76531.4]
  assign x471_A_sram_0_io_rPort_0_en_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@76530.4]
  assign x471_A_sram_0_io_rPort_0_backpressure = 1'h1; // @[MemInterfaceType.scala 66:44:@76529.4]
  assign x471_A_sram_0_io_wPort_0_ofs_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@76184.4]
  assign x471_A_sram_0_io_wPort_0_data_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@76183.4]
  assign x471_A_sram_0_io_wPort_0_en_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x471_A_sram_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@76179.4]
  assign x472_A_sram_1_clock = clock; // @[:@75898.4]
  assign x472_A_sram_1_reset = reset; // @[:@75899.4]
  assign x472_A_sram_1_io_rPort_0_ofs_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@76526.4]
  assign x472_A_sram_1_io_rPort_0_en_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@76525.4]
  assign x472_A_sram_1_io_rPort_0_backpressure = 1'h1; // @[MemInterfaceType.scala 66:44:@76524.4]
  assign x472_A_sram_1_io_wPort_0_ofs_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@76177.4]
  assign x472_A_sram_1_io_wPort_0_data_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@76176.4]
  assign x472_A_sram_1_io_wPort_0_en_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x472_A_sram_1_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@76172.4]
  assign x473_A_sram_2_clock = clock; // @[:@75915.4]
  assign x473_A_sram_2_reset = reset; // @[:@75916.4]
  assign x473_A_sram_2_io_rPort_0_ofs_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@76536.4]
  assign x473_A_sram_2_io_rPort_0_en_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@76535.4]
  assign x473_A_sram_2_io_rPort_0_backpressure = 1'h1; // @[MemInterfaceType.scala 66:44:@76534.4]
  assign x473_A_sram_2_io_wPort_0_ofs_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@76194.4]
  assign x473_A_sram_2_io_wPort_0_data_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@76193.4]
  assign x473_A_sram_2_io_wPort_0_en_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x473_A_sram_2_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@76189.4]
  assign x538_outr_UnitPipe_DenseTransfer_sm_clock = clock; // @[:@75980.4]
  assign x538_outr_UnitPipe_DenseTransfer_sm_reset = reset; // @[:@75981.4]
  assign x538_outr_UnitPipe_DenseTransfer_sm_io_enable = _T_263 & _T_272; // @[SpatialBlocks.scala 139:18:@76062.4]
  assign x538_outr_UnitPipe_DenseTransfer_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 141:21:@76064.4]
  assign x538_outr_UnitPipe_DenseTransfer_sm_io_doneIn_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@76032.4]
  assign x538_outr_UnitPipe_DenseTransfer_sm_io_doneIn_1 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:72:@76033.4]
  assign x538_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_0 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:95:@76079.4]
  assign x538_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_1 = x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:95:@76080.4]
  assign RetimeWrapper_clock = clock; // @[:@76043.4]
  assign RetimeWrapper_reset = reset; // @[:@76044.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@76046.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@76045.4]
  assign RetimeWrapper_1_clock = clock; // @[:@76051.4]
  assign RetimeWrapper_1_reset = reset; // @[:@76052.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@76054.4]
  assign RetimeWrapper_1_io_in = x538_outr_UnitPipe_DenseTransfer_sm_io_done; // @[package.scala 94:16:@76053.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_clock = clock; // @[:@76082.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_reset = reset; // @[:@76083.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x468_A_dram_number = io_in_x468_A_dram_number; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 59:30:@76171.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_valid = io_in_x476_valid; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 62:23:@76187.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x476_bits_rdata_0 = io_in_x476_bits_rdata_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 62:23:@76186.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_in_x474_ready = io_in_x474_ready; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 64:23:@76199.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_0 = x538_outr_UnitPipe_DenseTransfer_sm_io_enableOut_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 112:22:@76215.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_1 = x538_outr_UnitPipe_DenseTransfer_sm_io_enableOut_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 112:22:@76216.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_0 = x538_outr_UnitPipe_DenseTransfer_sm_io_childAck_0; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 112:22:@76211.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_1 = x538_outr_UnitPipe_DenseTransfer_sm_io_childAck_1; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 112:22:@76212.4]
  assign x538_outr_UnitPipe_DenseTransfer_kernelx538_outr_UnitPipe_DenseTransfer_concrete1_io_rr = io_rr; // @[sm_x538_outr_UnitPipe_DenseTransfer.scala 111:18:@76200.4]
  assign x539_out_sram_0_clock = clock; // @[:@76240.4]
  assign x539_out_sram_0_reset = reset; // @[:@76241.4]
  assign x539_out_sram_0_io_rPort_0_ofs_0 = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@76772.4]
  assign x539_out_sram_0_io_rPort_0_en_0 = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@76771.4]
  assign x539_out_sram_0_io_rPort_0_backpressure = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@76770.4]
  assign x539_out_sram_0_io_wPort_0_ofs_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_ofs_0; // @[MemInterfaceType.scala 67:44:@76543.4]
  assign x539_out_sram_0_io_wPort_0_data_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_data_0; // @[MemInterfaceType.scala 67:44:@76542.4]
  assign x539_out_sram_0_io_wPort_0_en_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x539_out_sram_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@76538.4]
  assign x541_ctrchain_clock = clock; // @[:@76257.4]
  assign x541_ctrchain_reset = reset; // @[:@76258.4]
  assign x541_ctrchain_io_input_reset = x668_outr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 158:100:@76434.4]
  assign x541_ctrchain_io_input_enable = x668_outr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 158:42:@76433.4]
  assign x668_outr_Foreach_sm_clock = clock; // @[:@76315.4]
  assign x668_outr_Foreach_sm_reset = reset; // @[:@76316.4]
  assign x668_outr_Foreach_sm_io_enable = _T_362 & _T_371; // @[SpatialBlocks.scala 139:18:@76413.4]
  assign x668_outr_Foreach_sm_io_ctrDone = io_rr ? _T_345 : 1'h0; // @[sm_RootController.scala 101:39:@76356.4]
  assign x668_outr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 141:21:@76415.4]
  assign x668_outr_Foreach_sm_io_doneIn_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@76383.4]
  assign x668_outr_Foreach_sm_io_doneIn_1 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:72:@76384.4]
  assign x668_outr_Foreach_sm_io_maskIn_0 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smMaskIn_0; // @[SpatialBlocks.scala 131:72:@76385.4]
  assign x668_outr_Foreach_sm_io_maskIn_1 = x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsOut_smMaskIn_1; // @[SpatialBlocks.scala 131:72:@76386.4]
  assign RetimeWrapper_2_clock = clock; // @[:@76349.4]
  assign RetimeWrapper_2_reset = reset; // @[:@76350.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@76352.4]
  assign RetimeWrapper_2_io_in = x541_ctrchain_io_output_done; // @[package.scala 94:16:@76351.4]
  assign RetimeWrapper_3_clock = clock; // @[:@76394.4]
  assign RetimeWrapper_3_reset = reset; // @[:@76395.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@76397.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@76396.4]
  assign RetimeWrapper_4_clock = clock; // @[:@76402.4]
  assign RetimeWrapper_4_reset = reset; // @[:@76403.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@76405.4]
  assign RetimeWrapper_4_io_in = x668_outr_Foreach_sm_io_done; // @[package.scala 94:16:@76404.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_clock = clock; // @[:@76436.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_reset = reset; // @[:@76437.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x472_A_sram_1_rPort_0_output_0 = x472_A_sram_1_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@76523.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x471_A_sram_0_rPort_0_output_0 = x471_A_sram_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@76528.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_in_x473_A_sram_2_rPort_0_output_0 = x473_A_sram_2_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@76533.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_0 = x668_outr_Foreach_sm_io_enableOut_0; // @[sm_x668_outr_Foreach.scala 118:22:@76555.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smEnableOuts_1 = x668_outr_Foreach_sm_io_enableOut_1; // @[sm_x668_outr_Foreach.scala 118:22:@76556.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smChildAcks_0 = x668_outr_Foreach_sm_io_childAck_0; // @[sm_x668_outr_Foreach.scala 118:22:@76551.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_smChildAcks_1 = x668_outr_Foreach_sm_io_childAck_1; // @[sm_x668_outr_Foreach.scala 118:22:@76552.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{23{x541_ctrchain_io_output_counts_0[8]}},x541_ctrchain_io_output_counts_0}; // @[sm_x668_outr_Foreach.scala 118:22:@76550.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x541_ctrchain_io_output_oobs_0; // @[sm_x668_outr_Foreach.scala 118:22:@76549.4]
  assign x668_outr_Foreach_kernelx668_outr_Foreach_concrete1_io_rr = io_rr; // @[sm_x668_outr_Foreach.scala 117:18:@76545.4]
  assign x724_outr_UnitPipe_DenseTransfer_sm_clock = clock; // @[:@76614.4]
  assign x724_outr_UnitPipe_DenseTransfer_sm_reset = reset; // @[:@76615.4]
  assign x724_outr_UnitPipe_DenseTransfer_sm_io_enable = _T_454 & _T_463; // @[SpatialBlocks.scala 139:18:@76686.4]
  assign x724_outr_UnitPipe_DenseTransfer_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 141:21:@76688.4]
  assign x724_outr_UnitPipe_DenseTransfer_sm_io_doneIn_0 = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@76658.4]
  assign x724_outr_UnitPipe_DenseTransfer_sm_io_ctrCopyDone_0 = x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:95:@76703.4]
  assign RetimeWrapper_5_clock = clock; // @[:@76667.4]
  assign RetimeWrapper_5_reset = reset; // @[:@76668.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@76670.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@76669.4]
  assign RetimeWrapper_6_clock = clock; // @[:@76675.4]
  assign RetimeWrapper_6_reset = reset; // @[:@76676.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@76678.4]
  assign RetimeWrapper_6_io_in = x724_outr_UnitPipe_DenseTransfer_sm_io_done; // @[package.scala 94:16:@76677.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_clock = clock; // @[:@76705.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_reset = reset; // @[:@76706.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x670_ready = io_in_x670_ready; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 58:23:@76763.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x669_ready = io_in_x669_ready; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 59:23:@76767.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x470_out_host_number = io_in_x470_out_host_number; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 60:32:@76768.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x539_out_sram_0_rPort_0_output_0 = x539_out_sram_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@76769.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_in_x671_valid = io_in_x671_valid; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 62:23:@76775.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smEnableOuts_0 = x724_outr_UnitPipe_DenseTransfer_sm_io_enableOut_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 95:22:@76785.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_sigsIn_smChildAcks_0 = x724_outr_UnitPipe_DenseTransfer_sm_io_childAck_0; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 95:22:@76783.4]
  assign x724_outr_UnitPipe_DenseTransfer_kernelx724_outr_UnitPipe_DenseTransfer_concrete1_io_rr = io_rr; // @[sm_x724_outr_UnitPipe_DenseTransfer.scala 94:18:@76777.4]
endmodule
module AccelUnit( // @[:@76805.2]
  input          clock, // @[:@76806.4]
  input          reset, // @[:@76807.4]
  input          io_enable, // @[:@76808.4]
  output         io_done, // @[:@76808.4]
  input          io_reset, // @[:@76808.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@76808.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@76808.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@76808.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@76808.4]
  output         io_memStreams_loads_0_data_ready, // @[:@76808.4]
  input          io_memStreams_loads_0_data_valid, // @[:@76808.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@76808.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@76808.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@76808.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@76808.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@76808.4]
  input          io_memStreams_stores_0_data_ready, // @[:@76808.4]
  output         io_memStreams_stores_0_data_valid, // @[:@76808.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@76808.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@76808.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@76808.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@76808.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@76808.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@76808.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@76808.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@76808.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@76808.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@76808.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@76808.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@76808.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@76808.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@76808.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@76808.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@76808.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@76808.4]
  input  [63:0]  io_memStreams_gathers_0_data_bits_0, // @[:@76808.4]
  input  [63:0]  io_memStreams_gathers_0_data_bits_1, // @[:@76808.4]
  input  [63:0]  io_memStreams_gathers_0_data_bits_2, // @[:@76808.4]
  input  [63:0]  io_memStreams_gathers_0_data_bits_3, // @[:@76808.4]
  input  [63:0]  io_memStreams_gathers_0_data_bits_4, // @[:@76808.4]
  input  [63:0]  io_memStreams_gathers_0_data_bits_5, // @[:@76808.4]
  input  [63:0]  io_memStreams_gathers_0_data_bits_6, // @[:@76808.4]
  input  [63:0]  io_memStreams_gathers_0_data_bits_7, // @[:@76808.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@76808.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@76808.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@76808.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@76808.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@76808.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@76808.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@76808.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@76808.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@76808.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@76808.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@76808.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@76808.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@76808.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@76808.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@76808.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@76808.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@76808.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@76808.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@76808.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@76808.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@76808.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@76808.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@76808.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@76808.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@76808.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@76808.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@76808.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@76808.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@76808.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@76808.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@76808.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@76808.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@76808.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@76808.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@76808.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@76808.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@76808.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@76808.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@76808.4]
  output         io_heap_0_req_valid, // @[:@76808.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@76808.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@76808.4]
  input          io_heap_0_resp_valid, // @[:@76808.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@76808.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@76808.4]
  input  [63:0]  io_argIns_0, // @[:@76808.4]
  input  [63:0]  io_argIns_1, // @[:@76808.4]
  input          io_argOuts_0_port_ready, // @[:@76808.4]
  output         io_argOuts_0_port_valid, // @[:@76808.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@76808.4]
  input  [63:0]  io_argOuts_0_echo // @[:@76808.4]
);
  wire  SingleCounter_clock; // @[Main.scala 42:32:@76909.4]
  wire  SingleCounter_reset; // @[Main.scala 42:32:@76909.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 42:32:@76909.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 42:32:@76909.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@76927.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@76927.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@76927.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@76927.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@76927.4]
  wire  SRFF_clock; // @[Main.scala 46:28:@76936.4]
  wire  SRFF_reset; // @[Main.scala 46:28:@76936.4]
  wire  SRFF_io_input_set; // @[Main.scala 46:28:@76936.4]
  wire  SRFF_io_input_reset; // @[Main.scala 46:28:@76936.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 46:28:@76936.4]
  wire  SRFF_io_output; // @[Main.scala 46:28:@76936.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@76985.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@76985.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@76985.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@76985.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@76985.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@76985.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@76985.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@76985.4]
  wire  RootController_sm_io_doneIn_1; // @[sm_RootController.scala 36:18:@76985.4]
  wire  RootController_sm_io_doneIn_2; // @[sm_RootController.scala 36:18:@76985.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@76985.4]
  wire  RootController_sm_io_enableOut_1; // @[sm_RootController.scala 36:18:@76985.4]
  wire  RootController_sm_io_enableOut_2; // @[sm_RootController.scala 36:18:@76985.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@76985.4]
  wire  RootController_sm_io_childAck_1; // @[sm_RootController.scala 36:18:@76985.4]
  wire  RootController_sm_io_childAck_2; // @[sm_RootController.scala 36:18:@76985.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@77027.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@77027.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@77027.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@77027.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@77027.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 118:24:@77101.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x468_A_dram_number; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_in_x670_ready; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_in_x670_valid; // @[sm_RootController.scala 118:24:@77101.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x670_bits_wdata_0; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_in_x670_bits_wstrb; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_in_x669_ready; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_in_x669_valid; // @[sm_RootController.scala 118:24:@77101.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x669_bits_addr; // @[sm_RootController.scala 118:24:@77101.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x669_bits_size; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_in_x476_ready; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_in_x476_valid; // @[sm_RootController.scala 118:24:@77101.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x476_bits_rdata_0; // @[sm_RootController.scala 118:24:@77101.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x470_out_host_number; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_in_x671_ready; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_in_x671_valid; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_in_x474_ready; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_in_x474_valid; // @[sm_RootController.scala 118:24:@77101.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x474_bits_addr; // @[sm_RootController.scala 118:24:@77101.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x474_bits_size; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_2; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_2; // @[sm_RootController.scala 118:24:@77101.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 118:24:@77101.4]
  wire  _T_567; // @[package.scala 96:25:@76932.4 package.scala 96:25:@76933.4]
  wire  _T_632; // @[Main.scala 48:50:@77023.4]
  wire  _T_633; // @[Main.scala 48:59:@77024.4]
  wire  _T_647; // @[package.scala 100:49:@77045.4]
  reg  _T_650; // @[package.scala 48:56:@77046.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 42:32:@76909.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@76927.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 46:28:@76936.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@76985.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_doneIn_1(RootController_sm_io_doneIn_1),
    .io_doneIn_2(RootController_sm_io_doneIn_2),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_enableOut_1(RootController_sm_io_enableOut_1),
    .io_enableOut_2(RootController_sm_io_enableOut_2),
    .io_childAck_0(RootController_sm_io_childAck_0),
    .io_childAck_1(RootController_sm_io_childAck_1),
    .io_childAck_2(RootController_sm_io_childAck_2)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@77027.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 118:24:@77101.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x468_A_dram_number(RootController_kernelRootController_concrete1_io_in_x468_A_dram_number),
    .io_in_x670_ready(RootController_kernelRootController_concrete1_io_in_x670_ready),
    .io_in_x670_valid(RootController_kernelRootController_concrete1_io_in_x670_valid),
    .io_in_x670_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x670_bits_wdata_0),
    .io_in_x670_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x670_bits_wstrb),
    .io_in_x669_ready(RootController_kernelRootController_concrete1_io_in_x669_ready),
    .io_in_x669_valid(RootController_kernelRootController_concrete1_io_in_x669_valid),
    .io_in_x669_bits_addr(RootController_kernelRootController_concrete1_io_in_x669_bits_addr),
    .io_in_x669_bits_size(RootController_kernelRootController_concrete1_io_in_x669_bits_size),
    .io_in_x476_ready(RootController_kernelRootController_concrete1_io_in_x476_ready),
    .io_in_x476_valid(RootController_kernelRootController_concrete1_io_in_x476_valid),
    .io_in_x476_bits_rdata_0(RootController_kernelRootController_concrete1_io_in_x476_bits_rdata_0),
    .io_in_x470_out_host_number(RootController_kernelRootController_concrete1_io_in_x470_out_host_number),
    .io_in_x671_ready(RootController_kernelRootController_concrete1_io_in_x671_ready),
    .io_in_x671_valid(RootController_kernelRootController_concrete1_io_in_x671_valid),
    .io_in_x474_ready(RootController_kernelRootController_concrete1_io_in_x474_ready),
    .io_in_x474_valid(RootController_kernelRootController_concrete1_io_in_x474_valid),
    .io_in_x474_bits_addr(RootController_kernelRootController_concrete1_io_in_x474_bits_addr),
    .io_in_x474_bits_size(RootController_kernelRootController_concrete1_io_in_x474_bits_size),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_2),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_567 = RetimeWrapper_io_out; // @[package.scala 96:25:@76932.4 package.scala 96:25:@76933.4]
  assign _T_632 = io_enable & _T_567; // @[Main.scala 48:50:@77023.4]
  assign _T_633 = ~ SRFF_io_output; // @[Main.scala 48:59:@77024.4]
  assign _T_647 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@77045.4]
  assign io_done = SRFF_io_output; // @[Main.scala 55:23:@77044.4]
  assign io_memStreams_loads_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x474_valid; // @[sm_RootController.scala 68:23:@77180.4]
  assign io_memStreams_loads_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x474_bits_addr; // @[sm_RootController.scala 68:23:@77179.4]
  assign io_memStreams_loads_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x474_bits_size; // @[sm_RootController.scala 68:23:@77178.4]
  assign io_memStreams_loads_0_data_ready = RootController_kernelRootController_concrete1_io_in_x476_ready; // @[sm_RootController.scala 65:23:@77173.4]
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x669_valid; // @[sm_RootController.scala 64:23:@77169.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x669_bits_addr; // @[sm_RootController.scala 64:23:@77168.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x669_bits_size; // @[sm_RootController.scala 64:23:@77167.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x670_valid; // @[sm_RootController.scala 63:23:@77165.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x670_bits_wdata_0; // @[sm_RootController.scala 63:23:@77164.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x670_bits_wstrb; // @[sm_RootController.scala 63:23:@77163.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x671_ready; // @[sm_RootController.scala 67:23:@77177.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 64'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = 1'h0;
  assign io_axiStreamsOut_0_TVALID = 1'h0;
  assign io_axiStreamsOut_0_TDATA = 256'h0;
  assign io_axiStreamsOut_0_TSTRB = 32'h0;
  assign io_axiStreamsOut_0_TKEEP = 32'h0;
  assign io_axiStreamsOut_0_TLAST = 1'h0;
  assign io_axiStreamsOut_0_TID = 8'h0;
  assign io_axiStreamsOut_0_TDEST = 8'h0;
  assign io_axiStreamsOut_0_TUSER = 32'h0;
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@76910.4]
  assign SingleCounter_reset = reset; // @[:@76911.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 43:79:@76925.4]
  assign RetimeWrapper_clock = clock; // @[:@76928.4]
  assign RetimeWrapper_reset = reset; // @[:@76929.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@76931.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@76930.4]
  assign SRFF_clock = clock; // @[:@76937.4]
  assign SRFF_reset = reset; // @[:@76938.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 64:29:@77219.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 53:31:@77042.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 54:36:@77043.4]
  assign RootController_sm_clock = clock; // @[:@76986.4]
  assign RootController_sm_reset = reset; // @[:@76987.4]
  assign RootController_sm_io_enable = _T_632 & _T_633; // @[Main.scala 52:33:@77041.4 SpatialBlocks.scala 139:18:@77086.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 133:15:@77080.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_650; // @[Main.scala 56:34:@77049.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:72:@77073.4]
  assign RootController_sm_io_doneIn_1 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:72:@77074.4]
  assign RootController_sm_io_doneIn_2 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:72:@77075.4]
  assign RetimeWrapper_1_clock = clock; // @[:@77028.4]
  assign RetimeWrapper_1_reset = reset; // @[:@77029.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@77031.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@77030.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@77102.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@77103.4]
  assign RootController_kernelRootController_concrete1_io_in_x468_A_dram_number = io_argIns_0; // @[sm_RootController.scala 62:30:@77162.4]
  assign RootController_kernelRootController_concrete1_io_in_x670_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 63:23:@77166.4]
  assign RootController_kernelRootController_concrete1_io_in_x669_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 64:23:@77170.4]
  assign RootController_kernelRootController_concrete1_io_in_x476_valid = io_memStreams_loads_0_data_valid; // @[sm_RootController.scala 65:23:@77172.4]
  assign RootController_kernelRootController_concrete1_io_in_x476_bits_rdata_0 = io_memStreams_loads_0_data_bits_rdata_0; // @[sm_RootController.scala 65:23:@77171.4]
  assign RootController_kernelRootController_concrete1_io_in_x470_out_host_number = io_argIns_1; // @[sm_RootController.scala 66:32:@77174.4]
  assign RootController_kernelRootController_concrete1_io_in_x671_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 67:23:@77176.4]
  assign RootController_kernelRootController_concrete1_io_in_x474_ready = io_memStreams_loads_0_cmd_ready; // @[sm_RootController.scala 68:23:@77181.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 123:22:@77194.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_1 = RootController_sm_io_enableOut_1; // @[sm_RootController.scala 123:22:@77195.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_2 = RootController_sm_io_enableOut_2; // @[sm_RootController.scala 123:22:@77196.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 123:22:@77188.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_1 = RootController_sm_io_childAck_1; // @[sm_RootController.scala 123:22:@77189.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_2 = RootController_sm_io_childAck_2; // @[sm_RootController.scala 123:22:@77190.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 122:18:@77182.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_650 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_650 <= 1'h0;
    end else begin
      _T_650 <= _T_647;
    end
  end
endmodule
module Counter( // @[:@77221.2]
  input        clock, // @[:@77222.4]
  input        reset, // @[:@77223.4]
  input        io_reset, // @[:@77224.4]
  input        io_enable, // @[:@77224.4]
  input  [5:0] io_stride, // @[:@77224.4]
  output [5:0] io_out, // @[:@77224.4]
  output [5:0] io_next // @[:@77224.4]
);
  reg [5:0] count; // @[Counter.scala 15:22:@77226.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_17; // @[Counter.scala 17:24:@77227.4]
  wire [5:0] newCount; // @[Counter.scala 17:24:@77228.4]
  wire [5:0] _GEN_0; // @[Counter.scala 21:26:@77233.6]
  wire [5:0] _GEN_1; // @[Counter.scala 19:18:@77229.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@77227.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@77228.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@77233.6]
  assign _GEN_1 = io_reset ? 6'h0 : _GEN_0; // @[Counter.scala 19:18:@77229.4]
  assign io_out = count; // @[Counter.scala 25:10:@77236.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@77237.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 6'h0;
    end else begin
      if (io_reset) begin
        count <= 6'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_76( // @[:@77273.2]
  input         clock, // @[:@77274.4]
  input         reset, // @[:@77275.4]
  input  [5:0]  io_raddr, // @[:@77276.4]
  input         io_wen, // @[:@77276.4]
  input  [5:0]  io_waddr, // @[:@77276.4]
  input  [63:0] io_wdata_addr, // @[:@77276.4]
  input  [31:0] io_wdata_size, // @[:@77276.4]
  output [63:0] io_rdata_addr, // @[:@77276.4]
  output [31:0] io_rdata_size, // @[:@77276.4]
  input         io_backpressure // @[:@77276.4]
);
  wire [95:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@77278.4]
  wire [95:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@77278.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@77278.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@77278.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@77278.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@77278.4]
  wire [5:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@77278.4]
  wire [5:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@77278.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@77278.4]
  wire [95:0] _T_17; // @[SRAM.scala 175:38:@77292.4]
  wire  _T_20; // @[SRAM.scala 182:49:@77297.4]
  wire  _T_21; // @[SRAM.scala 182:37:@77298.4]
  reg  _T_24; // @[SRAM.scala 182:29:@77299.4]
  reg [31:0] _RAND_0;
  reg [95:0] _T_28; // @[SRAM.scala 183:29:@77302.4]
  reg [95:0] _RAND_1;
  wire [95:0] _T_29; // @[SRAM.scala 184:22:@77304.4]
  SRAMVerilogAWS #(.DWIDTH(96), .WORDS(64), .AWIDTH(6)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@77278.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_17 = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:38:@77292.4]
  assign _T_20 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@77297.4]
  assign _T_21 = io_wen & _T_20; // @[SRAM.scala 182:37:@77298.4]
  assign _T_29 = _T_24 ? _T_28 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:22:@77304.4]
  assign io_rdata_addr = _T_29[95:32]; // @[SRAM.scala 184:16:@77313.4]
  assign io_rdata_size = _T_29[31:0]; // @[SRAM.scala 184:16:@77312.4]
  assign SRAMVerilogAWS_wdata = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:20:@77293.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@77294.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@77290.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@77296.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@77295.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@77291.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@77289.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@77288.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_24 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _T_28 = _RAND_1[95:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_21;
    end
    if (reset) begin
      _T_28 <= 96'h0;
    end else begin
      _T_28 <= _T_17;
    end
  end
endmodule
module FIFO( // @[:@77315.2]
  input         clock, // @[:@77316.4]
  input         reset, // @[:@77317.4]
  output        io_in_ready, // @[:@77318.4]
  input         io_in_valid, // @[:@77318.4]
  input  [63:0] io_in_bits_addr, // @[:@77318.4]
  input  [31:0] io_in_bits_size, // @[:@77318.4]
  input         io_out_ready, // @[:@77318.4]
  output        io_out_valid, // @[:@77318.4]
  output [63:0] io_out_bits_addr, // @[:@77318.4]
  output [31:0] io_out_bits_size // @[:@77318.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@77714.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@77714.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@77714.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@77714.4]
  wire [5:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@77714.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@77714.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@77714.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@77724.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@77724.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@77724.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@77724.4]
  wire [5:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@77724.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@77724.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@77724.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@77739.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@77739.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@77739.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@77739.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@77739.4]
  wire [63:0] SRAM_io_wdata_addr; // @[FIFO.scala 73:19:@77739.4]
  wire [31:0] SRAM_io_wdata_size; // @[FIFO.scala 73:19:@77739.4]
  wire [63:0] SRAM_io_rdata_addr; // @[FIFO.scala 73:19:@77739.4]
  wire [31:0] SRAM_io_rdata_size; // @[FIFO.scala 73:19:@77739.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@77739.4]
  wire  writeEn; // @[FIFO.scala 30:29:@77712.4]
  wire  readEn; // @[FIFO.scala 31:29:@77713.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@77734.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@77735.4]
  wire  _T_824; // @[FIFO.scala 45:27:@77736.4]
  wire  empty; // @[FIFO.scala 45:24:@77737.4]
  wire  full; // @[FIFO.scala 46:23:@77738.4]
  wire  _T_827; // @[FIFO.scala 83:17:@77751.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@77752.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@77714.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@77724.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_76 SRAM ( // @[FIFO.scala 73:19:@77739.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata_addr(SRAM_io_wdata_addr),
    .io_wdata_size(SRAM_io_wdata_size),
    .io_rdata_addr(SRAM_io_rdata_addr),
    .io_rdata_size(SRAM_io_rdata_size),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@77712.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@77713.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@77735.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@77736.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@77737.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@77738.4]
  assign _T_827 = writeEn != readEn; // @[FIFO.scala 83:17:@77751.4]
  assign _GEN_0 = _T_827 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@77752.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@77758.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@77756.4]
  assign io_out_bits_addr = SRAM_io_rdata_addr; // @[FIFO.scala 79:17:@77749.4]
  assign io_out_bits_size = SRAM_io_rdata_size; // @[FIFO.scala 79:17:@77748.4]
  assign enqCounter_clock = clock; // @[:@77715.4]
  assign enqCounter_reset = reset; // @[:@77716.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@77722.4]
  assign enqCounter_io_stride = 6'h1; // @[FIFO.scala 37:24:@77723.4]
  assign deqCounter_clock = clock; // @[:@77725.4]
  assign deqCounter_reset = reset; // @[:@77726.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@77732.4]
  assign deqCounter_io_stride = 6'h1; // @[FIFO.scala 41:24:@77733.4]
  assign SRAM_clock = clock; // @[:@77740.4]
  assign SRAM_reset = reset; // @[:@77741.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@77743.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@77744.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@77745.4]
  assign SRAM_io_wdata_addr = io_in_bits_addr; // @[FIFO.scala 78:16:@77747.4]
  assign SRAM_io_wdata_size = io_in_bits_size; // @[FIFO.scala 78:16:@77746.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@77750.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_827) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module Counter_2( // @[:@77760.2]
  input        clock, // @[:@77761.4]
  input        reset, // @[:@77762.4]
  input        io_reset, // @[:@77763.4]
  input        io_enable, // @[:@77763.4]
  input  [3:0] io_stride, // @[:@77763.4]
  output [3:0] io_out // @[:@77763.4]
);
  reg [3:0] count; // @[Counter.scala 15:22:@77765.4]
  reg [31:0] _RAND_0;
  wire [4:0] _T_17; // @[Counter.scala 17:24:@77766.4]
  wire [3:0] newCount; // @[Counter.scala 17:24:@77767.4]
  wire [3:0] _GEN_0; // @[Counter.scala 21:26:@77772.6]
  wire [3:0] _GEN_1; // @[Counter.scala 19:18:@77768.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@77766.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@77767.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@77772.6]
  assign _GEN_1 = io_reset ? 4'h0 : _GEN_0; // @[Counter.scala 19:18:@77768.4]
  assign io_out = count; // @[Counter.scala 25:10:@77775.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 4'h0;
    end else begin
      if (io_reset) begin
        count <= 4'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module Counter_4( // @[:@77796.2]
  input        clock, // @[:@77797.4]
  input        reset, // @[:@77798.4]
  input        io_reset, // @[:@77799.4]
  input        io_enable, // @[:@77799.4]
  input  [1:0] io_stride, // @[:@77799.4]
  output [1:0] io_out, // @[:@77799.4]
  output [1:0] io_next // @[:@77799.4]
);
  reg [1:0] count; // @[Counter.scala 15:22:@77801.4]
  reg [31:0] _RAND_0;
  wire [2:0] _T_17; // @[Counter.scala 17:24:@77802.4]
  wire [1:0] newCount; // @[Counter.scala 17:24:@77803.4]
  wire [1:0] _GEN_0; // @[Counter.scala 21:26:@77808.6]
  wire [1:0] _GEN_1; // @[Counter.scala 19:18:@77804.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@77802.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@77803.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@77808.6]
  assign _GEN_1 = io_reset ? 2'h0 : _GEN_0; // @[Counter.scala 19:18:@77804.4]
  assign io_out = count; // @[Counter.scala 25:10:@77811.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@77812.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 2'h0;
    end else begin
      if (io_reset) begin
        count <= 2'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_77( // @[:@77848.2]
  input         clock, // @[:@77849.4]
  input         reset, // @[:@77850.4]
  input  [1:0]  io_raddr, // @[:@77851.4]
  input         io_wen, // @[:@77851.4]
  input  [1:0]  io_waddr, // @[:@77851.4]
  input  [31:0] io_wdata, // @[:@77851.4]
  output [31:0] io_rdata, // @[:@77851.4]
  input         io_backpressure // @[:@77851.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@77853.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@77853.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@77853.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@77853.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@77853.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@77853.4]
  wire [1:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@77853.4]
  wire [1:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@77853.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@77853.4]
  wire  _T_19; // @[SRAM.scala 182:49:@77871.4]
  wire  _T_20; // @[SRAM.scala 182:37:@77872.4]
  reg  _T_23; // @[SRAM.scala 182:29:@77873.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@77875.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(4), .AWIDTH(2)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@77853.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@77871.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@77872.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@77880.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@77867.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@77868.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@77865.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@77870.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@77869.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@77866.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@77864.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@77863.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module FIFO_1( // @[:@77882.2]
  input         clock, // @[:@77883.4]
  input         reset, // @[:@77884.4]
  output        io_in_ready, // @[:@77885.4]
  input         io_in_valid, // @[:@77885.4]
  input  [31:0] io_in_bits, // @[:@77885.4]
  input         io_out_ready, // @[:@77885.4]
  output        io_out_valid, // @[:@77885.4]
  output [31:0] io_out_bits // @[:@77885.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@77911.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@77911.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@77911.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@77911.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@77911.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@77911.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@77911.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@77921.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@77921.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@77921.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@77921.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@77921.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@77921.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@77921.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@77936.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@77936.4]
  wire [1:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@77936.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@77936.4]
  wire [1:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@77936.4]
  wire [31:0] SRAM_io_wdata; // @[FIFO.scala 73:19:@77936.4]
  wire [31:0] SRAM_io_rdata; // @[FIFO.scala 73:19:@77936.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@77936.4]
  wire  writeEn; // @[FIFO.scala 30:29:@77909.4]
  wire  readEn; // @[FIFO.scala 31:29:@77910.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@77931.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@77932.4]
  wire  _T_104; // @[FIFO.scala 45:27:@77933.4]
  wire  empty; // @[FIFO.scala 45:24:@77934.4]
  wire  full; // @[FIFO.scala 46:23:@77935.4]
  wire  _T_107; // @[FIFO.scala 83:17:@77946.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@77947.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@77911.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@77921.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_77 SRAM ( // @[FIFO.scala 73:19:@77936.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@77909.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@77910.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@77932.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@77933.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@77934.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@77935.4]
  assign _T_107 = writeEn != readEn; // @[FIFO.scala 83:17:@77946.4]
  assign _GEN_0 = _T_107 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@77947.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@77953.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@77951.4]
  assign io_out_bits = SRAM_io_rdata; // @[FIFO.scala 79:17:@77944.4]
  assign enqCounter_clock = clock; // @[:@77912.4]
  assign enqCounter_reset = reset; // @[:@77913.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@77919.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@77920.4]
  assign deqCounter_clock = clock; // @[:@77922.4]
  assign deqCounter_reset = reset; // @[:@77923.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@77929.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@77930.4]
  assign SRAM_clock = clock; // @[:@77937.4]
  assign SRAM_reset = reset; // @[:@77938.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@77940.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@77941.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@77942.4]
  assign SRAM_io_wdata = io_in_bits; // @[FIFO.scala 78:16:@77943.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@77945.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_107) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec( // @[:@80340.2]
  input         clock, // @[:@80341.4]
  input         reset, // @[:@80342.4]
  output        io_in_ready, // @[:@80343.4]
  input         io_in_valid, // @[:@80343.4]
  input  [31:0] io_in_bits_0, // @[:@80343.4]
  input  [31:0] io_in_bits_1, // @[:@80343.4]
  input  [31:0] io_in_bits_2, // @[:@80343.4]
  input  [31:0] io_in_bits_3, // @[:@80343.4]
  input  [31:0] io_in_bits_4, // @[:@80343.4]
  input  [31:0] io_in_bits_5, // @[:@80343.4]
  input  [31:0] io_in_bits_6, // @[:@80343.4]
  input  [31:0] io_in_bits_7, // @[:@80343.4]
  input  [31:0] io_in_bits_8, // @[:@80343.4]
  input  [31:0] io_in_bits_9, // @[:@80343.4]
  input  [31:0] io_in_bits_10, // @[:@80343.4]
  input  [31:0] io_in_bits_11, // @[:@80343.4]
  input  [31:0] io_in_bits_12, // @[:@80343.4]
  input  [31:0] io_in_bits_13, // @[:@80343.4]
  input  [31:0] io_in_bits_14, // @[:@80343.4]
  input  [31:0] io_in_bits_15, // @[:@80343.4]
  input         io_out_ready, // @[:@80343.4]
  output        io_out_valid, // @[:@80343.4]
  output [31:0] io_out_bits_0, // @[:@80343.4]
  output [31:0] io_out_bits_1, // @[:@80343.4]
  output [31:0] io_out_bits_2, // @[:@80343.4]
  output [31:0] io_out_bits_3, // @[:@80343.4]
  output [31:0] io_out_bits_4, // @[:@80343.4]
  output [31:0] io_out_bits_5, // @[:@80343.4]
  output [31:0] io_out_bits_6, // @[:@80343.4]
  output [31:0] io_out_bits_7, // @[:@80343.4]
  output [31:0] io_out_bits_8, // @[:@80343.4]
  output [31:0] io_out_bits_9, // @[:@80343.4]
  output [31:0] io_out_bits_10, // @[:@80343.4]
  output [31:0] io_out_bits_11, // @[:@80343.4]
  output [31:0] io_out_bits_12, // @[:@80343.4]
  output [31:0] io_out_bits_13, // @[:@80343.4]
  output [31:0] io_out_bits_14, // @[:@80343.4]
  output [31:0] io_out_bits_15, // @[:@80343.4]
  input         io_chainEnq, // @[:@80343.4]
  input         io_chainDeq // @[:@80343.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@80347.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@80347.4]
  wire  enqCounter_io_reset; // @[FIFOVec.scala 24:26:@80347.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@80347.4]
  wire [3:0] enqCounter_io_stride; // @[FIFOVec.scala 24:26:@80347.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@80347.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@80358.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@80358.4]
  wire  deqCounter_io_reset; // @[FIFOVec.scala 28:26:@80358.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@80358.4]
  wire [3:0] deqCounter_io_stride; // @[FIFOVec.scala 28:26:@80358.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@80358.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@80371.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@80371.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@80371.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@80371.4]
  wire [31:0] fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@80371.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@80371.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@80371.4]
  wire [31:0] fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@80371.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@80406.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@80406.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@80406.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@80406.4]
  wire [31:0] fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@80406.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@80406.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@80406.4]
  wire [31:0] fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@80406.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@80441.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@80441.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@80441.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@80441.4]
  wire [31:0] fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@80441.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@80441.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@80441.4]
  wire [31:0] fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@80441.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@80476.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@80476.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@80476.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@80476.4]
  wire [31:0] fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@80476.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@80476.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@80476.4]
  wire [31:0] fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@80476.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@80511.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@80511.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@80511.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@80511.4]
  wire [31:0] fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@80511.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@80511.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@80511.4]
  wire [31:0] fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@80511.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@80546.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@80546.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@80546.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@80546.4]
  wire [31:0] fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@80546.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@80546.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@80546.4]
  wire [31:0] fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@80546.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@80581.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@80581.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@80581.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@80581.4]
  wire [31:0] fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@80581.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@80581.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@80581.4]
  wire [31:0] fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@80581.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@80616.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@80616.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@80616.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@80616.4]
  wire [31:0] fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@80616.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@80616.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@80616.4]
  wire [31:0] fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@80616.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@80651.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@80651.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@80651.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@80651.4]
  wire [31:0] fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@80651.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@80651.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@80651.4]
  wire [31:0] fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@80651.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@80686.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@80686.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@80686.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@80686.4]
  wire [31:0] fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@80686.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@80686.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@80686.4]
  wire [31:0] fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@80686.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@80721.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@80721.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@80721.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@80721.4]
  wire [31:0] fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@80721.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@80721.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@80721.4]
  wire [31:0] fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@80721.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@80756.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@80756.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@80756.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@80756.4]
  wire [31:0] fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@80756.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@80756.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@80756.4]
  wire [31:0] fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@80756.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@80791.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@80791.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@80791.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@80791.4]
  wire [31:0] fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@80791.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@80791.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@80791.4]
  wire [31:0] fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@80791.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@80826.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@80826.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@80826.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@80826.4]
  wire [31:0] fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@80826.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@80826.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@80826.4]
  wire [31:0] fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@80826.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@80861.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@80861.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@80861.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@80861.4]
  wire [31:0] fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@80861.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@80861.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@80861.4]
  wire [31:0] fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@80861.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@80896.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@80896.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@80896.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@80896.4]
  wire [31:0] fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@80896.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@80896.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@80896.4]
  wire [31:0] fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@80896.4]
  wire  readEn; // @[FIFOVec.scala 20:29:@80345.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@80346.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@80369.4]
  wire [15:0] deqDecoder; // @[OneHot.scala 45:35:@80370.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@80396.4]
  wire  _T_151; // @[FIFOVec.scala 42:25:@80397.4]
  wire  _T_154; // @[FIFOVec.scala 44:50:@80402.4]
  wire  _T_156; // @[FIFOVec.scala 44:26:@80403.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@80431.4]
  wire  _T_160; // @[FIFOVec.scala 42:25:@80432.4]
  wire  _T_163; // @[FIFOVec.scala 44:50:@80437.4]
  wire  _T_165; // @[FIFOVec.scala 44:26:@80438.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@80466.4]
  wire  _T_169; // @[FIFOVec.scala 42:25:@80467.4]
  wire  _T_172; // @[FIFOVec.scala 44:50:@80472.4]
  wire  _T_174; // @[FIFOVec.scala 44:26:@80473.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@80501.4]
  wire  _T_178; // @[FIFOVec.scala 42:25:@80502.4]
  wire  _T_181; // @[FIFOVec.scala 44:50:@80507.4]
  wire  _T_183; // @[FIFOVec.scala 44:26:@80508.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@80536.4]
  wire  _T_187; // @[FIFOVec.scala 42:25:@80537.4]
  wire  _T_190; // @[FIFOVec.scala 44:50:@80542.4]
  wire  _T_192; // @[FIFOVec.scala 44:26:@80543.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@80571.4]
  wire  _T_196; // @[FIFOVec.scala 42:25:@80572.4]
  wire  _T_199; // @[FIFOVec.scala 44:50:@80577.4]
  wire  _T_201; // @[FIFOVec.scala 44:26:@80578.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@80606.4]
  wire  _T_205; // @[FIFOVec.scala 42:25:@80607.4]
  wire  _T_208; // @[FIFOVec.scala 44:50:@80612.4]
  wire  _T_210; // @[FIFOVec.scala 44:26:@80613.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@80641.4]
  wire  _T_214; // @[FIFOVec.scala 42:25:@80642.4]
  wire  _T_217; // @[FIFOVec.scala 44:50:@80647.4]
  wire  _T_219; // @[FIFOVec.scala 44:26:@80648.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@80676.4]
  wire  _T_223; // @[FIFOVec.scala 42:25:@80677.4]
  wire  _T_226; // @[FIFOVec.scala 44:50:@80682.4]
  wire  _T_228; // @[FIFOVec.scala 44:26:@80683.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@80711.4]
  wire  _T_232; // @[FIFOVec.scala 42:25:@80712.4]
  wire  _T_235; // @[FIFOVec.scala 44:50:@80717.4]
  wire  _T_237; // @[FIFOVec.scala 44:26:@80718.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@80746.4]
  wire  _T_241; // @[FIFOVec.scala 42:25:@80747.4]
  wire  _T_244; // @[FIFOVec.scala 44:50:@80752.4]
  wire  _T_246; // @[FIFOVec.scala 44:26:@80753.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@80781.4]
  wire  _T_250; // @[FIFOVec.scala 42:25:@80782.4]
  wire  _T_253; // @[FIFOVec.scala 44:50:@80787.4]
  wire  _T_255; // @[FIFOVec.scala 44:26:@80788.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@80816.4]
  wire  _T_259; // @[FIFOVec.scala 42:25:@80817.4]
  wire  _T_262; // @[FIFOVec.scala 44:50:@80822.4]
  wire  _T_264; // @[FIFOVec.scala 44:26:@80823.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@80851.4]
  wire  _T_268; // @[FIFOVec.scala 42:25:@80852.4]
  wire  _T_271; // @[FIFOVec.scala 44:50:@80857.4]
  wire  _T_273; // @[FIFOVec.scala 44:26:@80858.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@80886.4]
  wire  _T_277; // @[FIFOVec.scala 42:25:@80887.4]
  wire  _T_280; // @[FIFOVec.scala 44:50:@80892.4]
  wire  _T_282; // @[FIFOVec.scala 44:26:@80893.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@80921.4]
  wire  _T_286; // @[FIFOVec.scala 42:25:@80922.4]
  wire  _T_289; // @[FIFOVec.scala 44:50:@80927.4]
  wire  _T_291; // @[FIFOVec.scala 44:26:@80928.4]
  wire  _T_316; // @[FIFOVec.scala 49:90:@80948.4]
  wire  _T_317; // @[FIFOVec.scala 49:90:@80949.4]
  wire  _T_318; // @[FIFOVec.scala 49:90:@80950.4]
  wire  _T_319; // @[FIFOVec.scala 49:90:@80951.4]
  wire  _T_320; // @[FIFOVec.scala 49:90:@80952.4]
  wire  _T_321; // @[FIFOVec.scala 49:90:@80953.4]
  wire  _T_322; // @[FIFOVec.scala 49:90:@80954.4]
  wire  _T_323; // @[FIFOVec.scala 49:90:@80955.4]
  wire  _T_324; // @[FIFOVec.scala 49:90:@80956.4]
  wire  _T_325; // @[FIFOVec.scala 49:90:@80957.4]
  wire  _T_326; // @[FIFOVec.scala 49:90:@80958.4]
  wire  _T_327; // @[FIFOVec.scala 49:90:@80959.4]
  wire  _T_328; // @[FIFOVec.scala 49:90:@80960.4]
  wire  _T_329; // @[FIFOVec.scala 49:90:@80961.4]
  wire  _T_330; // @[FIFOVec.scala 49:90:@80962.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80932.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80933.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@80963.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80934.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@80963.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80935.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@80963.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80936.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@80963.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80937.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@80963.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80938.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@80963.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80939.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@80963.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80940.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@80963.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80941.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@80963.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80942.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@80963.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80943.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@80963.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80944.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@80963.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80945.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@80963.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80946.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@80963.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80947.4]
  wire  _GEN_15; // @[FIFOVec.scala 49:21:@80963.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@80982.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@80983.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@80984.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@80985.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@80986.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@80987.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@80988.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@80989.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@80990.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@80991.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@80992.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@80993.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@80994.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@80995.4]
  wire  _T_369; // @[FIFOVec.scala 51:93:@80996.4]
  wire  _T_335_0; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80966.4]
  wire  _T_335_1; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80967.4]
  wire  _GEN_17; // @[FIFOVec.scala 51:22:@80997.4]
  wire  _T_335_2; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80968.4]
  wire  _GEN_18; // @[FIFOVec.scala 51:22:@80997.4]
  wire  _T_335_3; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80969.4]
  wire  _GEN_19; // @[FIFOVec.scala 51:22:@80997.4]
  wire  _T_335_4; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80970.4]
  wire  _GEN_20; // @[FIFOVec.scala 51:22:@80997.4]
  wire  _T_335_5; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80971.4]
  wire  _GEN_21; // @[FIFOVec.scala 51:22:@80997.4]
  wire  _T_335_6; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80972.4]
  wire  _GEN_22; // @[FIFOVec.scala 51:22:@80997.4]
  wire  _T_335_7; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80973.4]
  wire  _GEN_23; // @[FIFOVec.scala 51:22:@80997.4]
  wire  _T_335_8; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80974.4]
  wire  _GEN_24; // @[FIFOVec.scala 51:22:@80997.4]
  wire  _T_335_9; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80975.4]
  wire  _GEN_25; // @[FIFOVec.scala 51:22:@80997.4]
  wire  _T_335_10; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80976.4]
  wire  _GEN_26; // @[FIFOVec.scala 51:22:@80997.4]
  wire  _T_335_11; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80977.4]
  wire  _GEN_27; // @[FIFOVec.scala 51:22:@80997.4]
  wire  _T_335_12; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80978.4]
  wire  _GEN_28; // @[FIFOVec.scala 51:22:@80997.4]
  wire  _T_335_13; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80979.4]
  wire  _GEN_29; // @[FIFOVec.scala 51:22:@80997.4]
  wire  _T_335_14; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80980.4]
  wire  _GEN_30; // @[FIFOVec.scala 51:22:@80997.4]
  wire  _T_335_15; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80981.4]
  wire  _GEN_31; // @[FIFOVec.scala 51:22:@80997.4]
  wire [31:0] _T_374_0; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81000.4]
  wire [31:0] _T_374_1; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81001.4]
  wire [31:0] _GEN_33; // @[FIFOVec.scala 53:42:@81272.4]
  wire [31:0] _T_374_2; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81002.4]
  wire [31:0] _GEN_34; // @[FIFOVec.scala 53:42:@81272.4]
  wire [31:0] _T_374_3; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81003.4]
  wire [31:0] _GEN_35; // @[FIFOVec.scala 53:42:@81272.4]
  wire [31:0] _T_374_4; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81004.4]
  wire [31:0] _GEN_36; // @[FIFOVec.scala 53:42:@81272.4]
  wire [31:0] _T_374_5; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81005.4]
  wire [31:0] _GEN_37; // @[FIFOVec.scala 53:42:@81272.4]
  wire [31:0] _T_374_6; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81006.4]
  wire [31:0] _GEN_38; // @[FIFOVec.scala 53:42:@81272.4]
  wire [31:0] _T_374_7; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81007.4]
  wire [31:0] _GEN_39; // @[FIFOVec.scala 53:42:@81272.4]
  wire [31:0] _T_374_8; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81008.4]
  wire [31:0] _GEN_40; // @[FIFOVec.scala 53:42:@81272.4]
  wire [31:0] _T_374_9; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81009.4]
  wire [31:0] _GEN_41; // @[FIFOVec.scala 53:42:@81272.4]
  wire [31:0] _T_374_10; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81010.4]
  wire [31:0] _GEN_42; // @[FIFOVec.scala 53:42:@81272.4]
  wire [31:0] _T_374_11; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81011.4]
  wire [31:0] _GEN_43; // @[FIFOVec.scala 53:42:@81272.4]
  wire [31:0] _T_374_12; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81012.4]
  wire [31:0] _GEN_44; // @[FIFOVec.scala 53:42:@81272.4]
  wire [31:0] _T_374_13; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81013.4]
  wire [31:0] _GEN_45; // @[FIFOVec.scala 53:42:@81272.4]
  wire [31:0] _T_374_14; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81014.4]
  wire [31:0] _GEN_46; // @[FIFOVec.scala 53:42:@81272.4]
  wire [31:0] _T_374_15; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81015.4]
  wire [31:0] _GEN_47; // @[FIFOVec.scala 53:42:@81272.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@80347.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@80358.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out)
  );
  FIFO_1 fifos_0 ( // @[FIFOVec.scala 40:19:@80371.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_1 fifos_1 ( // @[FIFOVec.scala 40:19:@80406.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_1 fifos_2 ( // @[FIFOVec.scala 40:19:@80441.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_1 fifos_3 ( // @[FIFOVec.scala 40:19:@80476.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_1 fifos_4 ( // @[FIFOVec.scala 40:19:@80511.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_1 fifos_5 ( // @[FIFOVec.scala 40:19:@80546.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_1 fifos_6 ( // @[FIFOVec.scala 40:19:@80581.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_1 fifos_7 ( // @[FIFOVec.scala 40:19:@80616.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_1 fifos_8 ( // @[FIFOVec.scala 40:19:@80651.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_1 fifos_9 ( // @[FIFOVec.scala 40:19:@80686.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_1 fifos_10 ( // @[FIFOVec.scala 40:19:@80721.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_1 fifos_11 ( // @[FIFOVec.scala 40:19:@80756.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_1 fifos_12 ( // @[FIFOVec.scala 40:19:@80791.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_1 fifos_13 ( // @[FIFOVec.scala 40:19:@80826.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_1 fifos_14 ( // @[FIFOVec.scala 40:19:@80861.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_1 fifos_15 ( // @[FIFOVec.scala 40:19:@80896.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign readEn = io_out_valid & io_out_ready; // @[FIFOVec.scala 20:29:@80345.4]
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@80346.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@80369.4]
  assign deqDecoder = 16'h1 << deqCounter_io_out; // @[OneHot.scala 45:35:@80370.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@80396.4]
  assign _T_151 = io_chainEnq ? _T_149 : 1'h1; // @[FIFOVec.scala 42:25:@80397.4]
  assign _T_154 = deqDecoder[0]; // @[FIFOVec.scala 44:50:@80402.4]
  assign _T_156 = io_chainDeq ? _T_154 : 1'h1; // @[FIFOVec.scala 44:26:@80403.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@80431.4]
  assign _T_160 = io_chainEnq ? _T_158 : 1'h1; // @[FIFOVec.scala 42:25:@80432.4]
  assign _T_163 = deqDecoder[1]; // @[FIFOVec.scala 44:50:@80437.4]
  assign _T_165 = io_chainDeq ? _T_163 : 1'h1; // @[FIFOVec.scala 44:26:@80438.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@80466.4]
  assign _T_169 = io_chainEnq ? _T_167 : 1'h1; // @[FIFOVec.scala 42:25:@80467.4]
  assign _T_172 = deqDecoder[2]; // @[FIFOVec.scala 44:50:@80472.4]
  assign _T_174 = io_chainDeq ? _T_172 : 1'h1; // @[FIFOVec.scala 44:26:@80473.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@80501.4]
  assign _T_178 = io_chainEnq ? _T_176 : 1'h1; // @[FIFOVec.scala 42:25:@80502.4]
  assign _T_181 = deqDecoder[3]; // @[FIFOVec.scala 44:50:@80507.4]
  assign _T_183 = io_chainDeq ? _T_181 : 1'h1; // @[FIFOVec.scala 44:26:@80508.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@80536.4]
  assign _T_187 = io_chainEnq ? _T_185 : 1'h1; // @[FIFOVec.scala 42:25:@80537.4]
  assign _T_190 = deqDecoder[4]; // @[FIFOVec.scala 44:50:@80542.4]
  assign _T_192 = io_chainDeq ? _T_190 : 1'h1; // @[FIFOVec.scala 44:26:@80543.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@80571.4]
  assign _T_196 = io_chainEnq ? _T_194 : 1'h1; // @[FIFOVec.scala 42:25:@80572.4]
  assign _T_199 = deqDecoder[5]; // @[FIFOVec.scala 44:50:@80577.4]
  assign _T_201 = io_chainDeq ? _T_199 : 1'h1; // @[FIFOVec.scala 44:26:@80578.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@80606.4]
  assign _T_205 = io_chainEnq ? _T_203 : 1'h1; // @[FIFOVec.scala 42:25:@80607.4]
  assign _T_208 = deqDecoder[6]; // @[FIFOVec.scala 44:50:@80612.4]
  assign _T_210 = io_chainDeq ? _T_208 : 1'h1; // @[FIFOVec.scala 44:26:@80613.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@80641.4]
  assign _T_214 = io_chainEnq ? _T_212 : 1'h1; // @[FIFOVec.scala 42:25:@80642.4]
  assign _T_217 = deqDecoder[7]; // @[FIFOVec.scala 44:50:@80647.4]
  assign _T_219 = io_chainDeq ? _T_217 : 1'h1; // @[FIFOVec.scala 44:26:@80648.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@80676.4]
  assign _T_223 = io_chainEnq ? _T_221 : 1'h1; // @[FIFOVec.scala 42:25:@80677.4]
  assign _T_226 = deqDecoder[8]; // @[FIFOVec.scala 44:50:@80682.4]
  assign _T_228 = io_chainDeq ? _T_226 : 1'h1; // @[FIFOVec.scala 44:26:@80683.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@80711.4]
  assign _T_232 = io_chainEnq ? _T_230 : 1'h1; // @[FIFOVec.scala 42:25:@80712.4]
  assign _T_235 = deqDecoder[9]; // @[FIFOVec.scala 44:50:@80717.4]
  assign _T_237 = io_chainDeq ? _T_235 : 1'h1; // @[FIFOVec.scala 44:26:@80718.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@80746.4]
  assign _T_241 = io_chainEnq ? _T_239 : 1'h1; // @[FIFOVec.scala 42:25:@80747.4]
  assign _T_244 = deqDecoder[10]; // @[FIFOVec.scala 44:50:@80752.4]
  assign _T_246 = io_chainDeq ? _T_244 : 1'h1; // @[FIFOVec.scala 44:26:@80753.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@80781.4]
  assign _T_250 = io_chainEnq ? _T_248 : 1'h1; // @[FIFOVec.scala 42:25:@80782.4]
  assign _T_253 = deqDecoder[11]; // @[FIFOVec.scala 44:50:@80787.4]
  assign _T_255 = io_chainDeq ? _T_253 : 1'h1; // @[FIFOVec.scala 44:26:@80788.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@80816.4]
  assign _T_259 = io_chainEnq ? _T_257 : 1'h1; // @[FIFOVec.scala 42:25:@80817.4]
  assign _T_262 = deqDecoder[12]; // @[FIFOVec.scala 44:50:@80822.4]
  assign _T_264 = io_chainDeq ? _T_262 : 1'h1; // @[FIFOVec.scala 44:26:@80823.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@80851.4]
  assign _T_268 = io_chainEnq ? _T_266 : 1'h1; // @[FIFOVec.scala 42:25:@80852.4]
  assign _T_271 = deqDecoder[13]; // @[FIFOVec.scala 44:50:@80857.4]
  assign _T_273 = io_chainDeq ? _T_271 : 1'h1; // @[FIFOVec.scala 44:26:@80858.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@80886.4]
  assign _T_277 = io_chainEnq ? _T_275 : 1'h1; // @[FIFOVec.scala 42:25:@80887.4]
  assign _T_280 = deqDecoder[14]; // @[FIFOVec.scala 44:50:@80892.4]
  assign _T_282 = io_chainDeq ? _T_280 : 1'h1; // @[FIFOVec.scala 44:26:@80893.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@80921.4]
  assign _T_286 = io_chainEnq ? _T_284 : 1'h1; // @[FIFOVec.scala 42:25:@80922.4]
  assign _T_289 = deqDecoder[15]; // @[FIFOVec.scala 44:50:@80927.4]
  assign _T_291 = io_chainDeq ? _T_289 : 1'h1; // @[FIFOVec.scala 44:26:@80928.4]
  assign _T_316 = fifos_0_io_in_ready & fifos_1_io_in_ready; // @[FIFOVec.scala 49:90:@80948.4]
  assign _T_317 = _T_316 & fifos_2_io_in_ready; // @[FIFOVec.scala 49:90:@80949.4]
  assign _T_318 = _T_317 & fifos_3_io_in_ready; // @[FIFOVec.scala 49:90:@80950.4]
  assign _T_319 = _T_318 & fifos_4_io_in_ready; // @[FIFOVec.scala 49:90:@80951.4]
  assign _T_320 = _T_319 & fifos_5_io_in_ready; // @[FIFOVec.scala 49:90:@80952.4]
  assign _T_321 = _T_320 & fifos_6_io_in_ready; // @[FIFOVec.scala 49:90:@80953.4]
  assign _T_322 = _T_321 & fifos_7_io_in_ready; // @[FIFOVec.scala 49:90:@80954.4]
  assign _T_323 = _T_322 & fifos_8_io_in_ready; // @[FIFOVec.scala 49:90:@80955.4]
  assign _T_324 = _T_323 & fifos_9_io_in_ready; // @[FIFOVec.scala 49:90:@80956.4]
  assign _T_325 = _T_324 & fifos_10_io_in_ready; // @[FIFOVec.scala 49:90:@80957.4]
  assign _T_326 = _T_325 & fifos_11_io_in_ready; // @[FIFOVec.scala 49:90:@80958.4]
  assign _T_327 = _T_326 & fifos_12_io_in_ready; // @[FIFOVec.scala 49:90:@80959.4]
  assign _T_328 = _T_327 & fifos_13_io_in_ready; // @[FIFOVec.scala 49:90:@80960.4]
  assign _T_329 = _T_328 & fifos_14_io_in_ready; // @[FIFOVec.scala 49:90:@80961.4]
  assign _T_330 = _T_329 & fifos_15_io_in_ready; // @[FIFOVec.scala 49:90:@80962.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80932.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80933.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@80963.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80934.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@80963.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80935.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@80963.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80936.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@80963.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80937.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@80963.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80938.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@80963.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80939.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@80963.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80940.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@80963.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80941.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@80963.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80942.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@80963.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80943.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@80963.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80944.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@80963.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80945.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@80963.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80946.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@80963.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@80931.4 FIFOVec.scala 49:42:@80947.4]
  assign _GEN_15 = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:21:@80963.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@80982.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@80983.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@80984.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@80985.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@80986.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@80987.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@80988.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@80989.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@80990.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@80991.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@80992.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@80993.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@80994.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@80995.4]
  assign _T_369 = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:93:@80996.4]
  assign _T_335_0 = fifos_0_io_out_valid; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80966.4]
  assign _T_335_1 = fifos_1_io_out_valid; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80967.4]
  assign _GEN_17 = 4'h1 == deqCounter_io_out ? _T_335_1 : _T_335_0; // @[FIFOVec.scala 51:22:@80997.4]
  assign _T_335_2 = fifos_2_io_out_valid; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80968.4]
  assign _GEN_18 = 4'h2 == deqCounter_io_out ? _T_335_2 : _GEN_17; // @[FIFOVec.scala 51:22:@80997.4]
  assign _T_335_3 = fifos_3_io_out_valid; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80969.4]
  assign _GEN_19 = 4'h3 == deqCounter_io_out ? _T_335_3 : _GEN_18; // @[FIFOVec.scala 51:22:@80997.4]
  assign _T_335_4 = fifos_4_io_out_valid; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80970.4]
  assign _GEN_20 = 4'h4 == deqCounter_io_out ? _T_335_4 : _GEN_19; // @[FIFOVec.scala 51:22:@80997.4]
  assign _T_335_5 = fifos_5_io_out_valid; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80971.4]
  assign _GEN_21 = 4'h5 == deqCounter_io_out ? _T_335_5 : _GEN_20; // @[FIFOVec.scala 51:22:@80997.4]
  assign _T_335_6 = fifos_6_io_out_valid; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80972.4]
  assign _GEN_22 = 4'h6 == deqCounter_io_out ? _T_335_6 : _GEN_21; // @[FIFOVec.scala 51:22:@80997.4]
  assign _T_335_7 = fifos_7_io_out_valid; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80973.4]
  assign _GEN_23 = 4'h7 == deqCounter_io_out ? _T_335_7 : _GEN_22; // @[FIFOVec.scala 51:22:@80997.4]
  assign _T_335_8 = fifos_8_io_out_valid; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80974.4]
  assign _GEN_24 = 4'h8 == deqCounter_io_out ? _T_335_8 : _GEN_23; // @[FIFOVec.scala 51:22:@80997.4]
  assign _T_335_9 = fifos_9_io_out_valid; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80975.4]
  assign _GEN_25 = 4'h9 == deqCounter_io_out ? _T_335_9 : _GEN_24; // @[FIFOVec.scala 51:22:@80997.4]
  assign _T_335_10 = fifos_10_io_out_valid; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80976.4]
  assign _GEN_26 = 4'ha == deqCounter_io_out ? _T_335_10 : _GEN_25; // @[FIFOVec.scala 51:22:@80997.4]
  assign _T_335_11 = fifos_11_io_out_valid; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80977.4]
  assign _GEN_27 = 4'hb == deqCounter_io_out ? _T_335_11 : _GEN_26; // @[FIFOVec.scala 51:22:@80997.4]
  assign _T_335_12 = fifos_12_io_out_valid; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80978.4]
  assign _GEN_28 = 4'hc == deqCounter_io_out ? _T_335_12 : _GEN_27; // @[FIFOVec.scala 51:22:@80997.4]
  assign _T_335_13 = fifos_13_io_out_valid; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80979.4]
  assign _GEN_29 = 4'hd == deqCounter_io_out ? _T_335_13 : _GEN_28; // @[FIFOVec.scala 51:22:@80997.4]
  assign _T_335_14 = fifos_14_io_out_valid; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80980.4]
  assign _GEN_30 = 4'he == deqCounter_io_out ? _T_335_14 : _GEN_29; // @[FIFOVec.scala 51:22:@80997.4]
  assign _T_335_15 = fifos_15_io_out_valid; // @[FIFOVec.scala 51:43:@80965.4 FIFOVec.scala 51:43:@80981.4]
  assign _GEN_31 = 4'hf == deqCounter_io_out ? _T_335_15 : _GEN_30; // @[FIFOVec.scala 51:22:@80997.4]
  assign _T_374_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81000.4]
  assign _T_374_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81001.4]
  assign _GEN_33 = 4'h1 == deqCounter_io_out ? _T_374_1 : _T_374_0; // @[FIFOVec.scala 53:42:@81272.4]
  assign _T_374_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81002.4]
  assign _GEN_34 = 4'h2 == deqCounter_io_out ? _T_374_2 : _GEN_33; // @[FIFOVec.scala 53:42:@81272.4]
  assign _T_374_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81003.4]
  assign _GEN_35 = 4'h3 == deqCounter_io_out ? _T_374_3 : _GEN_34; // @[FIFOVec.scala 53:42:@81272.4]
  assign _T_374_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81004.4]
  assign _GEN_36 = 4'h4 == deqCounter_io_out ? _T_374_4 : _GEN_35; // @[FIFOVec.scala 53:42:@81272.4]
  assign _T_374_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81005.4]
  assign _GEN_37 = 4'h5 == deqCounter_io_out ? _T_374_5 : _GEN_36; // @[FIFOVec.scala 53:42:@81272.4]
  assign _T_374_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81006.4]
  assign _GEN_38 = 4'h6 == deqCounter_io_out ? _T_374_6 : _GEN_37; // @[FIFOVec.scala 53:42:@81272.4]
  assign _T_374_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81007.4]
  assign _GEN_39 = 4'h7 == deqCounter_io_out ? _T_374_7 : _GEN_38; // @[FIFOVec.scala 53:42:@81272.4]
  assign _T_374_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81008.4]
  assign _GEN_40 = 4'h8 == deqCounter_io_out ? _T_374_8 : _GEN_39; // @[FIFOVec.scala 53:42:@81272.4]
  assign _T_374_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81009.4]
  assign _GEN_41 = 4'h9 == deqCounter_io_out ? _T_374_9 : _GEN_40; // @[FIFOVec.scala 53:42:@81272.4]
  assign _T_374_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81010.4]
  assign _GEN_42 = 4'ha == deqCounter_io_out ? _T_374_10 : _GEN_41; // @[FIFOVec.scala 53:42:@81272.4]
  assign _T_374_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81011.4]
  assign _GEN_43 = 4'hb == deqCounter_io_out ? _T_374_11 : _GEN_42; // @[FIFOVec.scala 53:42:@81272.4]
  assign _T_374_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81012.4]
  assign _GEN_44 = 4'hc == deqCounter_io_out ? _T_374_12 : _GEN_43; // @[FIFOVec.scala 53:42:@81272.4]
  assign _T_374_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81013.4]
  assign _GEN_45 = 4'hd == deqCounter_io_out ? _T_374_13 : _GEN_44; // @[FIFOVec.scala 53:42:@81272.4]
  assign _T_374_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81014.4]
  assign _GEN_46 = 4'he == deqCounter_io_out ? _T_374_14 : _GEN_45; // @[FIFOVec.scala 53:42:@81272.4]
  assign _T_374_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:65:@80999.4 FIFOVec.scala 53:65:@81015.4]
  assign _GEN_47 = 4'hf == deqCounter_io_out ? _T_374_15 : _GEN_46; // @[FIFOVec.scala 53:42:@81272.4]
  assign io_in_ready = io_chainEnq ? _GEN_15 : _T_330; // @[FIFOVec.scala 49:15:@80964.4]
  assign io_out_valid = io_chainDeq ? _GEN_31 : _T_369; // @[FIFOVec.scala 51:16:@80998.4]
  assign io_out_bits_0 = io_chainDeq ? _GEN_47 : _T_374_0; // @[FIFOVec.scala 53:15:@81306.4]
  assign io_out_bits_1 = io_chainDeq ? _GEN_47 : _T_374_1; // @[FIFOVec.scala 53:15:@81307.4]
  assign io_out_bits_2 = io_chainDeq ? _GEN_47 : _T_374_2; // @[FIFOVec.scala 53:15:@81308.4]
  assign io_out_bits_3 = io_chainDeq ? _GEN_47 : _T_374_3; // @[FIFOVec.scala 53:15:@81309.4]
  assign io_out_bits_4 = io_chainDeq ? _GEN_47 : _T_374_4; // @[FIFOVec.scala 53:15:@81310.4]
  assign io_out_bits_5 = io_chainDeq ? _GEN_47 : _T_374_5; // @[FIFOVec.scala 53:15:@81311.4]
  assign io_out_bits_6 = io_chainDeq ? _GEN_47 : _T_374_6; // @[FIFOVec.scala 53:15:@81312.4]
  assign io_out_bits_7 = io_chainDeq ? _GEN_47 : _T_374_7; // @[FIFOVec.scala 53:15:@81313.4]
  assign io_out_bits_8 = io_chainDeq ? _GEN_47 : _T_374_8; // @[FIFOVec.scala 53:15:@81314.4]
  assign io_out_bits_9 = io_chainDeq ? _GEN_47 : _T_374_9; // @[FIFOVec.scala 53:15:@81315.4]
  assign io_out_bits_10 = io_chainDeq ? _GEN_47 : _T_374_10; // @[FIFOVec.scala 53:15:@81316.4]
  assign io_out_bits_11 = io_chainDeq ? _GEN_47 : _T_374_11; // @[FIFOVec.scala 53:15:@81317.4]
  assign io_out_bits_12 = io_chainDeq ? _GEN_47 : _T_374_12; // @[FIFOVec.scala 53:15:@81318.4]
  assign io_out_bits_13 = io_chainDeq ? _GEN_47 : _T_374_13; // @[FIFOVec.scala 53:15:@81319.4]
  assign io_out_bits_14 = io_chainDeq ? _GEN_47 : _T_374_14; // @[FIFOVec.scala 53:15:@81320.4]
  assign io_out_bits_15 = io_chainDeq ? _GEN_47 : _T_374_15; // @[FIFOVec.scala 53:15:@81321.4]
  assign enqCounter_clock = clock; // @[:@80348.4]
  assign enqCounter_reset = reset; // @[:@80349.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = writeEn & io_chainEnq; // @[FIFOVec.scala 26:24:@80356.4]
  assign enqCounter_io_stride = 4'h1; // @[FIFOVec.scala 27:24:@80357.4]
  assign deqCounter_clock = clock; // @[:@80359.4]
  assign deqCounter_reset = reset; // @[:@80360.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = readEn & io_chainDeq; // @[FIFOVec.scala 30:24:@80367.4]
  assign deqCounter_io_stride = 4'h1; // @[FIFOVec.scala 31:24:@80368.4]
  assign fifos_0_clock = clock; // @[:@80372.4]
  assign fifos_0_reset = reset; // @[:@80373.4]
  assign fifos_0_io_in_valid = _T_151 & writeEn; // @[FIFOVec.scala 42:19:@80399.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@80401.4]
  assign fifos_0_io_out_ready = _T_156 & readEn; // @[FIFOVec.scala 44:20:@80405.4]
  assign fifos_1_clock = clock; // @[:@80407.4]
  assign fifos_1_reset = reset; // @[:@80408.4]
  assign fifos_1_io_in_valid = _T_160 & writeEn; // @[FIFOVec.scala 42:19:@80434.4]
  assign fifos_1_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_1; // @[FIFOVec.scala 43:18:@80436.4]
  assign fifos_1_io_out_ready = _T_165 & readEn; // @[FIFOVec.scala 44:20:@80440.4]
  assign fifos_2_clock = clock; // @[:@80442.4]
  assign fifos_2_reset = reset; // @[:@80443.4]
  assign fifos_2_io_in_valid = _T_169 & writeEn; // @[FIFOVec.scala 42:19:@80469.4]
  assign fifos_2_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_2; // @[FIFOVec.scala 43:18:@80471.4]
  assign fifos_2_io_out_ready = _T_174 & readEn; // @[FIFOVec.scala 44:20:@80475.4]
  assign fifos_3_clock = clock; // @[:@80477.4]
  assign fifos_3_reset = reset; // @[:@80478.4]
  assign fifos_3_io_in_valid = _T_178 & writeEn; // @[FIFOVec.scala 42:19:@80504.4]
  assign fifos_3_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_3; // @[FIFOVec.scala 43:18:@80506.4]
  assign fifos_3_io_out_ready = _T_183 & readEn; // @[FIFOVec.scala 44:20:@80510.4]
  assign fifos_4_clock = clock; // @[:@80512.4]
  assign fifos_4_reset = reset; // @[:@80513.4]
  assign fifos_4_io_in_valid = _T_187 & writeEn; // @[FIFOVec.scala 42:19:@80539.4]
  assign fifos_4_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_4; // @[FIFOVec.scala 43:18:@80541.4]
  assign fifos_4_io_out_ready = _T_192 & readEn; // @[FIFOVec.scala 44:20:@80545.4]
  assign fifos_5_clock = clock; // @[:@80547.4]
  assign fifos_5_reset = reset; // @[:@80548.4]
  assign fifos_5_io_in_valid = _T_196 & writeEn; // @[FIFOVec.scala 42:19:@80574.4]
  assign fifos_5_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_5; // @[FIFOVec.scala 43:18:@80576.4]
  assign fifos_5_io_out_ready = _T_201 & readEn; // @[FIFOVec.scala 44:20:@80580.4]
  assign fifos_6_clock = clock; // @[:@80582.4]
  assign fifos_6_reset = reset; // @[:@80583.4]
  assign fifos_6_io_in_valid = _T_205 & writeEn; // @[FIFOVec.scala 42:19:@80609.4]
  assign fifos_6_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_6; // @[FIFOVec.scala 43:18:@80611.4]
  assign fifos_6_io_out_ready = _T_210 & readEn; // @[FIFOVec.scala 44:20:@80615.4]
  assign fifos_7_clock = clock; // @[:@80617.4]
  assign fifos_7_reset = reset; // @[:@80618.4]
  assign fifos_7_io_in_valid = _T_214 & writeEn; // @[FIFOVec.scala 42:19:@80644.4]
  assign fifos_7_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_7; // @[FIFOVec.scala 43:18:@80646.4]
  assign fifos_7_io_out_ready = _T_219 & readEn; // @[FIFOVec.scala 44:20:@80650.4]
  assign fifos_8_clock = clock; // @[:@80652.4]
  assign fifos_8_reset = reset; // @[:@80653.4]
  assign fifos_8_io_in_valid = _T_223 & writeEn; // @[FIFOVec.scala 42:19:@80679.4]
  assign fifos_8_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_8; // @[FIFOVec.scala 43:18:@80681.4]
  assign fifos_8_io_out_ready = _T_228 & readEn; // @[FIFOVec.scala 44:20:@80685.4]
  assign fifos_9_clock = clock; // @[:@80687.4]
  assign fifos_9_reset = reset; // @[:@80688.4]
  assign fifos_9_io_in_valid = _T_232 & writeEn; // @[FIFOVec.scala 42:19:@80714.4]
  assign fifos_9_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_9; // @[FIFOVec.scala 43:18:@80716.4]
  assign fifos_9_io_out_ready = _T_237 & readEn; // @[FIFOVec.scala 44:20:@80720.4]
  assign fifos_10_clock = clock; // @[:@80722.4]
  assign fifos_10_reset = reset; // @[:@80723.4]
  assign fifos_10_io_in_valid = _T_241 & writeEn; // @[FIFOVec.scala 42:19:@80749.4]
  assign fifos_10_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_10; // @[FIFOVec.scala 43:18:@80751.4]
  assign fifos_10_io_out_ready = _T_246 & readEn; // @[FIFOVec.scala 44:20:@80755.4]
  assign fifos_11_clock = clock; // @[:@80757.4]
  assign fifos_11_reset = reset; // @[:@80758.4]
  assign fifos_11_io_in_valid = _T_250 & writeEn; // @[FIFOVec.scala 42:19:@80784.4]
  assign fifos_11_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_11; // @[FIFOVec.scala 43:18:@80786.4]
  assign fifos_11_io_out_ready = _T_255 & readEn; // @[FIFOVec.scala 44:20:@80790.4]
  assign fifos_12_clock = clock; // @[:@80792.4]
  assign fifos_12_reset = reset; // @[:@80793.4]
  assign fifos_12_io_in_valid = _T_259 & writeEn; // @[FIFOVec.scala 42:19:@80819.4]
  assign fifos_12_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_12; // @[FIFOVec.scala 43:18:@80821.4]
  assign fifos_12_io_out_ready = _T_264 & readEn; // @[FIFOVec.scala 44:20:@80825.4]
  assign fifos_13_clock = clock; // @[:@80827.4]
  assign fifos_13_reset = reset; // @[:@80828.4]
  assign fifos_13_io_in_valid = _T_268 & writeEn; // @[FIFOVec.scala 42:19:@80854.4]
  assign fifos_13_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_13; // @[FIFOVec.scala 43:18:@80856.4]
  assign fifos_13_io_out_ready = _T_273 & readEn; // @[FIFOVec.scala 44:20:@80860.4]
  assign fifos_14_clock = clock; // @[:@80862.4]
  assign fifos_14_reset = reset; // @[:@80863.4]
  assign fifos_14_io_in_valid = _T_277 & writeEn; // @[FIFOVec.scala 42:19:@80889.4]
  assign fifos_14_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_14; // @[FIFOVec.scala 43:18:@80891.4]
  assign fifos_14_io_out_ready = _T_282 & readEn; // @[FIFOVec.scala 44:20:@80895.4]
  assign fifos_15_clock = clock; // @[:@80897.4]
  assign fifos_15_reset = reset; // @[:@80898.4]
  assign fifos_15_io_in_valid = _T_286 & writeEn; // @[FIFOVec.scala 42:19:@80924.4]
  assign fifos_15_io_in_bits = io_chainEnq ? io_in_bits_0 : io_in_bits_15; // @[FIFOVec.scala 43:18:@80926.4]
  assign fifos_15_io_out_ready = _T_291 & readEn; // @[FIFOVec.scala 44:20:@80930.4]
endmodule
module SRAM_93( // @[:@81411.2]
  input        clock, // @[:@81412.4]
  input  [5:0] io_raddr, // @[:@81414.4]
  input        io_wen, // @[:@81414.4]
  input  [5:0] io_waddr // @[:@81414.4]
);
  wire [7:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@81416.4]
  wire [7:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@81416.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@81416.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@81416.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@81416.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@81416.4]
  wire [5:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@81416.4]
  wire [5:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@81416.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@81416.4]
  SRAMVerilogAWS #(.DWIDTH(8), .WORDS(64), .AWIDTH(6)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@81416.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign SRAMVerilogAWS_wdata = 8'h0; // @[SRAM.scala 175:20:@81430.4]
  assign SRAMVerilogAWS_backpressure = 1'h1; // @[SRAM.scala 176:27:@81431.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@81428.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@81433.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@81432.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@81429.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@81427.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@81426.4]
endmodule
module FIFO_17( // @[:@81445.2]
  input   clock, // @[:@81446.4]
  input   reset, // @[:@81447.4]
  output  io_in_ready, // @[:@81448.4]
  input   io_in_valid // @[:@81448.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@81714.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@81714.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@81714.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@81714.4]
  wire [5:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@81714.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@81714.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@81714.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@81724.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@81724.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@81724.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@81724.4]
  wire [5:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@81724.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@81724.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@81724.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@81739.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@81739.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@81739.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@81739.4]
  wire  writeEn; // @[FIFO.scala 30:29:@81712.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@81734.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@81735.4]
  wire  full; // @[FIFO.scala 46:23:@81738.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@81750.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@81714.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@81724.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_93 SRAM ( // @[FIFO.scala 73:19:@81739.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@81712.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@81735.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@81738.4]
  assign _GEN_0 = writeEn ? writeEn : maybeFull; // @[FIFO.scala 83:29:@81750.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@81756.4]
  assign enqCounter_clock = clock; // @[:@81715.4]
  assign enqCounter_reset = reset; // @[:@81716.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@81722.4]
  assign enqCounter_io_stride = 6'h1; // @[FIFO.scala 37:24:@81723.4]
  assign deqCounter_clock = clock; // @[:@81725.4]
  assign deqCounter_reset = reset; // @[:@81726.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = 1'h0; // @[FIFO.scala 40:24:@81732.4]
  assign deqCounter_io_stride = 6'h1; // @[FIFO.scala 41:24:@81733.4]
  assign SRAM_clock = clock; // @[:@81740.4]
  assign SRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 75:16:@81743.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@81744.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@81745.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (writeEn) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_1( // @[:@81758.2]
  input   clock, // @[:@81759.4]
  input   reset, // @[:@81760.4]
  output  io_in_ready, // @[:@81761.4]
  input   io_in_valid // @[:@81761.4]
);
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@81789.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@81789.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@81789.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@81789.4]
  FIFO_17 fifos_0 ( // @[FIFOVec.scala 40:19:@81789.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid)
  );
  assign io_in_ready = fifos_0_io_in_ready; // @[FIFOVec.scala 49:15:@82067.4]
  assign fifos_0_clock = clock; // @[:@81790.4]
  assign fifos_0_reset = reset; // @[:@81791.4]
  assign fifos_0_io_in_valid = io_in_valid & io_in_ready; // @[FIFOVec.scala 42:19:@82057.4]
endmodule
module FIFOWidthConvert( // @[:@82081.2]
  input         clock, // @[:@82082.4]
  input         reset, // @[:@82083.4]
  output        io_in_ready, // @[:@82084.4]
  input         io_in_valid, // @[:@82084.4]
  input  [63:0] io_in_bits_data_0, // @[:@82084.4]
  input  [63:0] io_in_bits_data_1, // @[:@82084.4]
  input  [63:0] io_in_bits_data_2, // @[:@82084.4]
  input  [63:0] io_in_bits_data_3, // @[:@82084.4]
  input  [63:0] io_in_bits_data_4, // @[:@82084.4]
  input  [63:0] io_in_bits_data_5, // @[:@82084.4]
  input  [63:0] io_in_bits_data_6, // @[:@82084.4]
  input  [63:0] io_in_bits_data_7, // @[:@82084.4]
  input         io_out_ready, // @[:@82084.4]
  output        io_out_valid, // @[:@82084.4]
  output [31:0] io_out_bits_data_0 // @[:@82084.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_in_bits_1; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_in_bits_2; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_in_bits_3; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_in_bits_4; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_in_bits_5; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_in_bits_6; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_in_bits_7; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_in_bits_8; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_in_bits_9; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_in_bits_10; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_in_bits_11; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_in_bits_12; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_in_bits_13; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_in_bits_14; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_in_bits_15; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_out_bits_1; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_out_bits_2; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_out_bits_3; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_out_bits_4; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_out_bits_5; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_out_bits_6; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_out_bits_7; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_out_bits_8; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_out_bits_9; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_out_bits_10; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_out_bits_11; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_out_bits_12; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_out_bits_13; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_out_bits_14; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire [31:0] FIFOVec_io_out_bits_15; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire  FIFOVec_io_chainEnq; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire  FIFOVec_io_chainDeq; // @[FIFOWidthConvert.scala 82:22:@82086.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 83:26:@82127.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 83:26:@82127.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 83:26:@82127.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 83:26:@82127.4]
  wire [511:0] _T_53; // @[Cat.scala 30:58:@82150.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 82:22:@82086.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_in_bits_1(FIFOVec_io_in_bits_1),
    .io_in_bits_2(FIFOVec_io_in_bits_2),
    .io_in_bits_3(FIFOVec_io_in_bits_3),
    .io_in_bits_4(FIFOVec_io_in_bits_4),
    .io_in_bits_5(FIFOVec_io_in_bits_5),
    .io_in_bits_6(FIFOVec_io_in_bits_6),
    .io_in_bits_7(FIFOVec_io_in_bits_7),
    .io_in_bits_8(FIFOVec_io_in_bits_8),
    .io_in_bits_9(FIFOVec_io_in_bits_9),
    .io_in_bits_10(FIFOVec_io_in_bits_10),
    .io_in_bits_11(FIFOVec_io_in_bits_11),
    .io_in_bits_12(FIFOVec_io_in_bits_12),
    .io_in_bits_13(FIFOVec_io_in_bits_13),
    .io_in_bits_14(FIFOVec_io_in_bits_14),
    .io_in_bits_15(FIFOVec_io_in_bits_15),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0),
    .io_out_bits_1(FIFOVec_io_out_bits_1),
    .io_out_bits_2(FIFOVec_io_out_bits_2),
    .io_out_bits_3(FIFOVec_io_out_bits_3),
    .io_out_bits_4(FIFOVec_io_out_bits_4),
    .io_out_bits_5(FIFOVec_io_out_bits_5),
    .io_out_bits_6(FIFOVec_io_out_bits_6),
    .io_out_bits_7(FIFOVec_io_out_bits_7),
    .io_out_bits_8(FIFOVec_io_out_bits_8),
    .io_out_bits_9(FIFOVec_io_out_bits_9),
    .io_out_bits_10(FIFOVec_io_out_bits_10),
    .io_out_bits_11(FIFOVec_io_out_bits_11),
    .io_out_bits_12(FIFOVec_io_out_bits_12),
    .io_out_bits_13(FIFOVec_io_out_bits_13),
    .io_out_bits_14(FIFOVec_io_out_bits_14),
    .io_out_bits_15(FIFOVec_io_out_bits_15),
    .io_chainEnq(FIFOVec_io_chainEnq),
    .io_chainDeq(FIFOVec_io_chainDeq)
  );
  FIFOVec_1 FIFOVec_1 ( // @[FIFOWidthConvert.scala 83:26:@82127.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid)
  );
  assign _T_53 = {io_in_bits_data_7,io_in_bits_data_6,io_in_bits_data_5,io_in_bits_data_4,io_in_bits_data_3,io_in_bits_data_2,io_in_bits_data_1,io_in_bits_data_0}; // @[Cat.scala 30:58:@82150.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 88:17:@82142.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 89:18:@82143.4]
  assign io_out_bits_data_0 = FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 96:22:@82208.4]
  assign FIFOVec_clock = clock; // @[:@82087.4]
  assign FIFOVec_reset = reset; // @[:@82088.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 92:22:@82200.4]
  assign FIFOVec_io_in_bits_0 = _T_53[31:0]; // @[FIFOWidthConvert.scala 91:21:@82184.4]
  assign FIFOVec_io_in_bits_1 = _T_53[63:32]; // @[FIFOWidthConvert.scala 91:21:@82185.4]
  assign FIFOVec_io_in_bits_2 = _T_53[95:64]; // @[FIFOWidthConvert.scala 91:21:@82186.4]
  assign FIFOVec_io_in_bits_3 = _T_53[127:96]; // @[FIFOWidthConvert.scala 91:21:@82187.4]
  assign FIFOVec_io_in_bits_4 = _T_53[159:128]; // @[FIFOWidthConvert.scala 91:21:@82188.4]
  assign FIFOVec_io_in_bits_5 = _T_53[191:160]; // @[FIFOWidthConvert.scala 91:21:@82189.4]
  assign FIFOVec_io_in_bits_6 = _T_53[223:192]; // @[FIFOWidthConvert.scala 91:21:@82190.4]
  assign FIFOVec_io_in_bits_7 = _T_53[255:224]; // @[FIFOWidthConvert.scala 91:21:@82191.4]
  assign FIFOVec_io_in_bits_8 = _T_53[287:256]; // @[FIFOWidthConvert.scala 91:21:@82192.4]
  assign FIFOVec_io_in_bits_9 = _T_53[319:288]; // @[FIFOWidthConvert.scala 91:21:@82193.4]
  assign FIFOVec_io_in_bits_10 = _T_53[351:320]; // @[FIFOWidthConvert.scala 91:21:@82194.4]
  assign FIFOVec_io_in_bits_11 = _T_53[383:352]; // @[FIFOWidthConvert.scala 91:21:@82195.4]
  assign FIFOVec_io_in_bits_12 = _T_53[415:384]; // @[FIFOWidthConvert.scala 91:21:@82196.4]
  assign FIFOVec_io_in_bits_13 = _T_53[447:416]; // @[FIFOWidthConvert.scala 91:21:@82197.4]
  assign FIFOVec_io_in_bits_14 = _T_53[479:448]; // @[FIFOWidthConvert.scala 91:21:@82198.4]
  assign FIFOVec_io_in_bits_15 = _T_53[511:480]; // @[FIFOWidthConvert.scala 91:21:@82199.4]
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 98:23:@82222.4]
  assign FIFOVec_io_chainEnq = 1'h0; // @[FIFOWidthConvert.scala 84:22:@82138.4]
  assign FIFOVec_io_chainDeq = 1'h1; // @[FIFOWidthConvert.scala 85:22:@82139.4]
  assign FIFOVec_1_clock = clock; // @[:@82128.4]
  assign FIFOVec_1_reset = reset; // @[:@82129.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 94:26:@82202.4]
endmodule
module StreamControllerLoad( // @[:@82224.2]
  input         clock, // @[:@82225.4]
  input         reset, // @[:@82226.4]
  input         io_dram_cmd_ready, // @[:@82227.4]
  output        io_dram_cmd_valid, // @[:@82227.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@82227.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@82227.4]
  output        io_dram_rresp_ready, // @[:@82227.4]
  input         io_dram_rresp_valid, // @[:@82227.4]
  input  [63:0] io_dram_rresp_bits_rdata_0, // @[:@82227.4]
  input  [63:0] io_dram_rresp_bits_rdata_1, // @[:@82227.4]
  input  [63:0] io_dram_rresp_bits_rdata_2, // @[:@82227.4]
  input  [63:0] io_dram_rresp_bits_rdata_3, // @[:@82227.4]
  input  [63:0] io_dram_rresp_bits_rdata_4, // @[:@82227.4]
  input  [63:0] io_dram_rresp_bits_rdata_5, // @[:@82227.4]
  input  [63:0] io_dram_rresp_bits_rdata_6, // @[:@82227.4]
  input  [63:0] io_dram_rresp_bits_rdata_7, // @[:@82227.4]
  output        io_load_cmd_ready, // @[:@82227.4]
  input         io_load_cmd_valid, // @[:@82227.4]
  input  [63:0] io_load_cmd_bits_addr, // @[:@82227.4]
  input  [31:0] io_load_cmd_bits_size, // @[:@82227.4]
  input         io_load_data_ready, // @[:@82227.4]
  output        io_load_data_valid, // @[:@82227.4]
  output [31:0] io_load_data_bits_rdata_0 // @[:@82227.4]
);
  wire  cmd_clock; // @[StreamController.scala 38:19:@82332.4]
  wire  cmd_reset; // @[StreamController.scala 38:19:@82332.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 38:19:@82332.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 38:19:@82332.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 38:19:@82332.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 38:19:@82332.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 38:19:@82332.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 38:19:@82332.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 38:19:@82332.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 38:19:@82332.4]
  wire  rdata_clock; // @[StreamController.scala 51:21:@82738.4]
  wire  rdata_reset; // @[StreamController.scala 51:21:@82738.4]
  wire  rdata_io_in_ready; // @[StreamController.scala 51:21:@82738.4]
  wire  rdata_io_in_valid; // @[StreamController.scala 51:21:@82738.4]
  wire [63:0] rdata_io_in_bits_data_0; // @[StreamController.scala 51:21:@82738.4]
  wire [63:0] rdata_io_in_bits_data_1; // @[StreamController.scala 51:21:@82738.4]
  wire [63:0] rdata_io_in_bits_data_2; // @[StreamController.scala 51:21:@82738.4]
  wire [63:0] rdata_io_in_bits_data_3; // @[StreamController.scala 51:21:@82738.4]
  wire [63:0] rdata_io_in_bits_data_4; // @[StreamController.scala 51:21:@82738.4]
  wire [63:0] rdata_io_in_bits_data_5; // @[StreamController.scala 51:21:@82738.4]
  wire [63:0] rdata_io_in_bits_data_6; // @[StreamController.scala 51:21:@82738.4]
  wire [63:0] rdata_io_in_bits_data_7; // @[StreamController.scala 51:21:@82738.4]
  wire  rdata_io_out_ready; // @[StreamController.scala 51:21:@82738.4]
  wire  rdata_io_out_valid; // @[StreamController.scala 51:21:@82738.4]
  wire [31:0] rdata_io_out_bits_data_0; // @[StreamController.scala 51:21:@82738.4]
  wire [25:0] _T_95; // @[StreamController.scala 21:10:@82735.4]
  FIFO cmd ( // @[StreamController.scala 38:19:@82332.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert rdata ( // @[StreamController.scala 51:21:@82738.4]
    .clock(rdata_clock),
    .reset(rdata_reset),
    .io_in_ready(rdata_io_in_ready),
    .io_in_valid(rdata_io_in_valid),
    .io_in_bits_data_0(rdata_io_in_bits_data_0),
    .io_in_bits_data_1(rdata_io_in_bits_data_1),
    .io_in_bits_data_2(rdata_io_in_bits_data_2),
    .io_in_bits_data_3(rdata_io_in_bits_data_3),
    .io_in_bits_data_4(rdata_io_in_bits_data_4),
    .io_in_bits_data_5(rdata_io_in_bits_data_5),
    .io_in_bits_data_6(rdata_io_in_bits_data_6),
    .io_in_bits_data_7(rdata_io_in_bits_data_7),
    .io_out_ready(rdata_io_out_ready),
    .io_out_valid(rdata_io_out_valid),
    .io_out_bits_data_0(rdata_io_out_bits_data_0)
  );
  assign _T_95 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@82735.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 44:21:@82732.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 46:25:@82733.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_95}; // @[StreamController.scala 48:25:@82736.4]
  assign io_dram_rresp_ready = rdata_io_in_ready; // @[StreamController.scala 55:23:@82765.4]
  assign io_load_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 42:21:@82730.4]
  assign io_load_data_valid = rdata_io_out_valid; // @[StreamController.scala 57:22:@82766.4]
  assign io_load_data_bits_rdata_0 = rdata_io_out_bits_data_0; // @[StreamController.scala 58:27:@82767.4]
  assign cmd_clock = clock; // @[:@82333.4]
  assign cmd_reset = reset; // @[:@82334.4]
  assign cmd_io_in_valid = io_load_cmd_valid; // @[StreamController.scala 40:19:@82727.4]
  assign cmd_io_in_bits_addr = io_load_cmd_bits_addr; // @[StreamController.scala 41:18:@82729.4]
  assign cmd_io_in_bits_size = io_load_cmd_bits_size; // @[StreamController.scala 41:18:@82728.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 43:20:@82731.4]
  assign rdata_clock = clock; // @[:@82739.4]
  assign rdata_reset = reset; // @[:@82740.4]
  assign rdata_io_in_valid = io_dram_rresp_valid; // @[StreamController.scala 54:21:@82764.4]
  assign rdata_io_in_bits_data_0 = io_dram_rresp_bits_rdata_0; // @[StreamController.scala 53:25:@82756.4]
  assign rdata_io_in_bits_data_1 = io_dram_rresp_bits_rdata_1; // @[StreamController.scala 53:25:@82757.4]
  assign rdata_io_in_bits_data_2 = io_dram_rresp_bits_rdata_2; // @[StreamController.scala 53:25:@82758.4]
  assign rdata_io_in_bits_data_3 = io_dram_rresp_bits_rdata_3; // @[StreamController.scala 53:25:@82759.4]
  assign rdata_io_in_bits_data_4 = io_dram_rresp_bits_rdata_4; // @[StreamController.scala 53:25:@82760.4]
  assign rdata_io_in_bits_data_5 = io_dram_rresp_bits_rdata_5; // @[StreamController.scala 53:25:@82761.4]
  assign rdata_io_in_bits_data_6 = io_dram_rresp_bits_rdata_6; // @[StreamController.scala 53:25:@82762.4]
  assign rdata_io_in_bits_data_7 = io_dram_rresp_bits_rdata_7; // @[StreamController.scala 53:25:@82763.4]
  assign rdata_io_out_ready = io_load_data_ready; // @[StreamController.scala 59:22:@82768.4]
endmodule
module FFRAM( // @[:@86944.2]
  input        clock, // @[:@86945.4]
  input        reset, // @[:@86946.4]
  input  [1:0] io_raddr, // @[:@86947.4]
  input        io_wen, // @[:@86947.4]
  input  [1:0] io_waddr, // @[:@86947.4]
  input        io_wdata, // @[:@86947.4]
  output       io_rdata, // @[:@86947.4]
  input        io_banks_0_wdata_valid, // @[:@86947.4]
  input        io_banks_0_wdata_bits, // @[:@86947.4]
  input        io_banks_1_wdata_valid, // @[:@86947.4]
  input        io_banks_1_wdata_bits, // @[:@86947.4]
  input        io_banks_2_wdata_valid, // @[:@86947.4]
  input        io_banks_2_wdata_bits, // @[:@86947.4]
  input        io_banks_3_wdata_valid, // @[:@86947.4]
  input        io_banks_3_wdata_bits // @[:@86947.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@86951.4]
  reg [31:0] _RAND_0;
  wire  _T_88; // @[SRAM.scala 148:37:@86952.4]
  wire  _T_89; // @[SRAM.scala 148:25:@86953.4]
  wire  _T_90; // @[SRAM.scala 148:15:@86954.4]
  wire  _T_91; // @[SRAM.scala 149:15:@86956.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@86955.4]
  reg  regs_1; // @[SRAM.scala 145:20:@86962.4]
  reg [31:0] _RAND_1;
  wire  _T_97; // @[SRAM.scala 148:37:@86963.4]
  wire  _T_98; // @[SRAM.scala 148:25:@86964.4]
  wire  _T_99; // @[SRAM.scala 148:15:@86965.4]
  wire  _T_100; // @[SRAM.scala 149:15:@86967.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@86966.4]
  reg  regs_2; // @[SRAM.scala 145:20:@86973.4]
  reg [31:0] _RAND_2;
  wire  _T_106; // @[SRAM.scala 148:37:@86974.4]
  wire  _T_107; // @[SRAM.scala 148:25:@86975.4]
  wire  _T_108; // @[SRAM.scala 148:15:@86976.4]
  wire  _T_109; // @[SRAM.scala 149:15:@86978.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@86977.4]
  reg  regs_3; // @[SRAM.scala 145:20:@86984.4]
  reg [31:0] _RAND_3;
  wire  _T_115; // @[SRAM.scala 148:37:@86985.4]
  wire  _T_116; // @[SRAM.scala 148:25:@86986.4]
  wire  _T_117; // @[SRAM.scala 148:15:@86987.4]
  wire  _T_118; // @[SRAM.scala 149:15:@86989.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@86988.4]
  wire  _GEN_5; // @[SRAM.scala 155:12:@86998.4]
  wire  _GEN_6; // @[SRAM.scala 155:12:@86998.4]
  assign _T_88 = io_waddr == 2'h0; // @[SRAM.scala 148:37:@86952.4]
  assign _T_89 = io_wen & _T_88; // @[SRAM.scala 148:25:@86953.4]
  assign _T_90 = io_banks_0_wdata_valid | _T_89; // @[SRAM.scala 148:15:@86954.4]
  assign _T_91 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@86956.6]
  assign _GEN_0 = _T_90 ? _T_91 : regs_0; // @[SRAM.scala 148:48:@86955.4]
  assign _T_97 = io_waddr == 2'h1; // @[SRAM.scala 148:37:@86963.4]
  assign _T_98 = io_wen & _T_97; // @[SRAM.scala 148:25:@86964.4]
  assign _T_99 = io_banks_1_wdata_valid | _T_98; // @[SRAM.scala 148:15:@86965.4]
  assign _T_100 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@86967.6]
  assign _GEN_1 = _T_99 ? _T_100 : regs_1; // @[SRAM.scala 148:48:@86966.4]
  assign _T_106 = io_waddr == 2'h2; // @[SRAM.scala 148:37:@86974.4]
  assign _T_107 = io_wen & _T_106; // @[SRAM.scala 148:25:@86975.4]
  assign _T_108 = io_banks_2_wdata_valid | _T_107; // @[SRAM.scala 148:15:@86976.4]
  assign _T_109 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@86978.6]
  assign _GEN_2 = _T_108 ? _T_109 : regs_2; // @[SRAM.scala 148:48:@86977.4]
  assign _T_115 = io_waddr == 2'h3; // @[SRAM.scala 148:37:@86985.4]
  assign _T_116 = io_wen & _T_115; // @[SRAM.scala 148:25:@86986.4]
  assign _T_117 = io_banks_3_wdata_valid | _T_116; // @[SRAM.scala 148:15:@86987.4]
  assign _T_118 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@86989.6]
  assign _GEN_3 = _T_117 ? _T_118 : regs_3; // @[SRAM.scala 148:48:@86988.4]
  assign _GEN_5 = 2'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@86998.4]
  assign _GEN_6 = 2'h2 == io_raddr ? regs_2 : _GEN_5; // @[SRAM.scala 155:12:@86998.4]
  assign io_rdata = 2'h3 == io_raddr ? regs_3 : _GEN_6; // @[SRAM.scala 155:12:@86998.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_90) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_99) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_108) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_117) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_35( // @[:@87000.2]
  input   clock, // @[:@87001.4]
  input   reset, // @[:@87002.4]
  output  io_in_ready, // @[:@87003.4]
  input   io_in_valid, // @[:@87003.4]
  input   io_in_bits, // @[:@87003.4]
  input   io_out_ready, // @[:@87003.4]
  output  io_out_valid, // @[:@87003.4]
  output  io_out_bits // @[:@87003.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@87029.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@87029.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@87029.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@87029.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@87029.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@87029.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@87029.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@87039.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@87039.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@87039.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@87039.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@87039.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@87039.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@87039.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@87054.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@87054.4]
  wire [1:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@87054.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@87054.4]
  wire [1:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@87054.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@87054.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@87054.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@87054.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@87054.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@87054.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@87054.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@87054.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@87054.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@87054.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@87054.4]
  wire  writeEn; // @[FIFO.scala 30:29:@87027.4]
  wire  readEn; // @[FIFO.scala 31:29:@87028.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@87049.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@87050.4]
  wire  _T_104; // @[FIFO.scala 45:27:@87051.4]
  wire  empty; // @[FIFO.scala 45:24:@87052.4]
  wire  full; // @[FIFO.scala 46:23:@87053.4]
  wire  _T_157; // @[FIFO.scala 83:17:@87140.4]
  wire  _GEN_4; // @[FIFO.scala 83:29:@87141.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@87029.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@87039.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM FFRAM ( // @[FIFO.scala 49:19:@87054.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@87027.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@87028.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@87050.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@87051.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@87052.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@87053.4]
  assign _T_157 = writeEn != readEn; // @[FIFO.scala 83:17:@87140.4]
  assign _GEN_4 = _T_157 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@87141.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@87147.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@87145.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@87079.4]
  assign enqCounter_clock = clock; // @[:@87030.4]
  assign enqCounter_reset = reset; // @[:@87031.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@87037.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@87038.4]
  assign deqCounter_clock = clock; // @[:@87040.4]
  assign deqCounter_reset = reset; // @[:@87041.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@87047.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@87048.4]
  assign FFRAM_clock = clock; // @[:@87055.4]
  assign FFRAM_reset = reset; // @[:@87056.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@87075.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@87076.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@87077.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@87078.4]
  assign FFRAM_io_banks_0_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@87081.4]
  assign FFRAM_io_banks_0_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@87080.4]
  assign FFRAM_io_banks_1_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@87084.4]
  assign FFRAM_io_banks_1_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@87083.4]
  assign FFRAM_io_banks_2_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@87087.4]
  assign FFRAM_io_banks_2_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@87086.4]
  assign FFRAM_io_banks_3_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@87090.4]
  assign FFRAM_io_banks_3_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@87089.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_157) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_3( // @[:@90764.2]
  input   clock, // @[:@90765.4]
  input   reset, // @[:@90766.4]
  output  io_in_ready, // @[:@90767.4]
  input   io_in_valid, // @[:@90767.4]
  input   io_in_bits_0, // @[:@90767.4]
  input   io_out_ready, // @[:@90767.4]
  output  io_out_valid, // @[:@90767.4]
  output  io_out_bits_0, // @[:@90767.4]
  output  io_out_bits_1, // @[:@90767.4]
  output  io_out_bits_2, // @[:@90767.4]
  output  io_out_bits_3, // @[:@90767.4]
  output  io_out_bits_4, // @[:@90767.4]
  output  io_out_bits_5, // @[:@90767.4]
  output  io_out_bits_6, // @[:@90767.4]
  output  io_out_bits_7, // @[:@90767.4]
  output  io_out_bits_8, // @[:@90767.4]
  output  io_out_bits_9, // @[:@90767.4]
  output  io_out_bits_10, // @[:@90767.4]
  output  io_out_bits_11, // @[:@90767.4]
  output  io_out_bits_12, // @[:@90767.4]
  output  io_out_bits_13, // @[:@90767.4]
  output  io_out_bits_14, // @[:@90767.4]
  output  io_out_bits_15 // @[:@90767.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@90771.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@90771.4]
  wire  enqCounter_io_reset; // @[FIFOVec.scala 24:26:@90771.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@90771.4]
  wire [3:0] enqCounter_io_stride; // @[FIFOVec.scala 24:26:@90771.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@90771.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@90782.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@90782.4]
  wire  deqCounter_io_reset; // @[FIFOVec.scala 28:26:@90782.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@90782.4]
  wire [3:0] deqCounter_io_stride; // @[FIFOVec.scala 28:26:@90782.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@90782.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@90795.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@90795.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@90795.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@90795.4]
  wire  fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@90795.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@90795.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@90795.4]
  wire  fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@90795.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@90830.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@90830.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@90830.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@90830.4]
  wire  fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@90830.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@90830.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@90830.4]
  wire  fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@90830.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@90865.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@90865.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@90865.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@90865.4]
  wire  fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@90865.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@90865.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@90865.4]
  wire  fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@90865.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@90900.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@90900.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@90900.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@90900.4]
  wire  fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@90900.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@90900.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@90900.4]
  wire  fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@90900.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@90935.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@90935.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@90935.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@90935.4]
  wire  fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@90935.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@90935.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@90935.4]
  wire  fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@90935.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@90970.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@90970.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@90970.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@90970.4]
  wire  fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@90970.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@90970.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@90970.4]
  wire  fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@90970.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@91005.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@91005.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@91005.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@91005.4]
  wire  fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@91005.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@91005.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@91005.4]
  wire  fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@91005.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@91040.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@91040.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@91040.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@91040.4]
  wire  fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@91040.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@91040.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@91040.4]
  wire  fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@91040.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@91075.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@91075.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@91075.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@91075.4]
  wire  fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@91075.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@91075.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@91075.4]
  wire  fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@91075.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@91110.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@91110.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@91110.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@91110.4]
  wire  fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@91110.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@91110.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@91110.4]
  wire  fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@91110.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@91145.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@91145.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@91145.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@91145.4]
  wire  fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@91145.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@91145.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@91145.4]
  wire  fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@91145.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@91180.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@91180.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@91180.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@91180.4]
  wire  fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@91180.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@91180.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@91180.4]
  wire  fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@91180.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@91215.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@91215.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@91215.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@91215.4]
  wire  fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@91215.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@91215.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@91215.4]
  wire  fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@91215.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@91250.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@91250.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@91250.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@91250.4]
  wire  fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@91250.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@91250.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@91250.4]
  wire  fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@91250.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@91285.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@91285.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@91285.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@91285.4]
  wire  fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@91285.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@91285.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@91285.4]
  wire  fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@91285.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@91320.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@91320.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@91320.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@91320.4]
  wire  fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@91320.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@91320.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@91320.4]
  wire  fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@91320.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@90770.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@90793.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@90820.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@90855.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@90890.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@90925.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@90960.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@90995.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@91030.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@91065.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@91100.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@91135.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@91170.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@91205.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@91240.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@91275.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@91310.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@91345.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91356.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91357.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@91387.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91358.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@91387.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91359.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@91387.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91360.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@91387.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91361.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@91387.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91362.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@91387.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91363.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@91387.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91364.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@91387.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91365.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@91387.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91366.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@91387.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91367.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@91387.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91368.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@91387.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91369.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@91387.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91370.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@91387.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91371.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@91406.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@91407.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@91408.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@91409.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@91410.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@91411.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@91412.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@91413.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@91414.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@91415.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@91416.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@91417.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@91418.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@91419.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@90771.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@90782.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out)
  );
  FIFO_35 fifos_0 ( // @[FIFOVec.scala 40:19:@90795.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_35 fifos_1 ( // @[FIFOVec.scala 40:19:@90830.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_35 fifos_2 ( // @[FIFOVec.scala 40:19:@90865.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_35 fifos_3 ( // @[FIFOVec.scala 40:19:@90900.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_35 fifos_4 ( // @[FIFOVec.scala 40:19:@90935.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_35 fifos_5 ( // @[FIFOVec.scala 40:19:@90970.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_35 fifos_6 ( // @[FIFOVec.scala 40:19:@91005.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_35 fifos_7 ( // @[FIFOVec.scala 40:19:@91040.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_35 fifos_8 ( // @[FIFOVec.scala 40:19:@91075.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_35 fifos_9 ( // @[FIFOVec.scala 40:19:@91110.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_35 fifos_10 ( // @[FIFOVec.scala 40:19:@91145.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_35 fifos_11 ( // @[FIFOVec.scala 40:19:@91180.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_35 fifos_12 ( // @[FIFOVec.scala 40:19:@91215.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_35 fifos_13 ( // @[FIFOVec.scala 40:19:@91250.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_35 fifos_14 ( // @[FIFOVec.scala 40:19:@91285.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_35 fifos_15 ( // @[FIFOVec.scala 40:19:@91320.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@90770.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@90793.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@90820.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@90855.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@90890.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@90925.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@90960.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@90995.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@91030.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@91065.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@91100.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@91135.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@91170.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@91205.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@91240.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@91275.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@91310.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@91345.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91356.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91357.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@91387.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91358.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@91387.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91359.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@91387.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91360.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@91387.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91361.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@91387.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91362.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@91387.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91363.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@91387.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91364.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@91387.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91365.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@91387.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91366.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@91387.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91367.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@91387.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91368.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@91387.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91369.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@91387.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91370.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@91387.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@91355.4 FIFOVec.scala 49:42:@91371.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@91406.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@91407.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@91408.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@91409.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@91410.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@91411.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@91412.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@91413.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@91414.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@91415.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@91416.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@91417.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@91418.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@91419.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@91388.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@91422.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@91730.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@91731.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@91732.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@91733.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@91734.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@91735.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@91736.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@91737.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@91738.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@91739.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@91740.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@91741.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@91742.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@91743.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@91744.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@91745.4]
  assign enqCounter_clock = clock; // @[:@90772.4]
  assign enqCounter_reset = reset; // @[:@90773.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@90780.4]
  assign enqCounter_io_stride = 4'h1; // @[FIFOVec.scala 27:24:@90781.4]
  assign deqCounter_clock = clock; // @[:@90783.4]
  assign deqCounter_reset = reset; // @[:@90784.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@90791.4]
  assign deqCounter_io_stride = 4'h1; // @[FIFOVec.scala 31:24:@90792.4]
  assign fifos_0_clock = clock; // @[:@90796.4]
  assign fifos_0_reset = reset; // @[:@90797.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@90823.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@90825.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@90829.4]
  assign fifos_1_clock = clock; // @[:@90831.4]
  assign fifos_1_reset = reset; // @[:@90832.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@90858.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@90860.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@90864.4]
  assign fifos_2_clock = clock; // @[:@90866.4]
  assign fifos_2_reset = reset; // @[:@90867.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@90893.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@90895.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@90899.4]
  assign fifos_3_clock = clock; // @[:@90901.4]
  assign fifos_3_reset = reset; // @[:@90902.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@90928.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@90930.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@90934.4]
  assign fifos_4_clock = clock; // @[:@90936.4]
  assign fifos_4_reset = reset; // @[:@90937.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@90963.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@90965.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@90969.4]
  assign fifos_5_clock = clock; // @[:@90971.4]
  assign fifos_5_reset = reset; // @[:@90972.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@90998.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@91000.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@91004.4]
  assign fifos_6_clock = clock; // @[:@91006.4]
  assign fifos_6_reset = reset; // @[:@91007.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@91033.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@91035.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@91039.4]
  assign fifos_7_clock = clock; // @[:@91041.4]
  assign fifos_7_reset = reset; // @[:@91042.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@91068.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@91070.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@91074.4]
  assign fifos_8_clock = clock; // @[:@91076.4]
  assign fifos_8_reset = reset; // @[:@91077.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@91103.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@91105.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@91109.4]
  assign fifos_9_clock = clock; // @[:@91111.4]
  assign fifos_9_reset = reset; // @[:@91112.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@91138.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@91140.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@91144.4]
  assign fifos_10_clock = clock; // @[:@91146.4]
  assign fifos_10_reset = reset; // @[:@91147.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@91173.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@91175.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@91179.4]
  assign fifos_11_clock = clock; // @[:@91181.4]
  assign fifos_11_reset = reset; // @[:@91182.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@91208.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@91210.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@91214.4]
  assign fifos_12_clock = clock; // @[:@91216.4]
  assign fifos_12_reset = reset; // @[:@91217.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@91243.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@91245.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@91249.4]
  assign fifos_13_clock = clock; // @[:@91251.4]
  assign fifos_13_reset = reset; // @[:@91252.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@91278.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@91280.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@91284.4]
  assign fifos_14_clock = clock; // @[:@91286.4]
  assign fifos_14_reset = reset; // @[:@91287.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@91313.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@91315.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@91319.4]
  assign fifos_15_clock = clock; // @[:@91321.4]
  assign fifos_15_reset = reset; // @[:@91322.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@91348.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@91350.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@91354.4]
endmodule
module FIFOWidthConvert_1( // @[:@91747.2]
  input         clock, // @[:@91748.4]
  input         reset, // @[:@91749.4]
  output        io_in_ready, // @[:@91750.4]
  input         io_in_valid, // @[:@91750.4]
  input  [31:0] io_in_bits_data_0, // @[:@91750.4]
  input         io_in_bits_strobe, // @[:@91750.4]
  input         io_out_ready, // @[:@91750.4]
  output        io_out_valid, // @[:@91750.4]
  output [63:0] io_out_bits_data_0, // @[:@91750.4]
  output [63:0] io_out_bits_data_1, // @[:@91750.4]
  output [63:0] io_out_bits_data_2, // @[:@91750.4]
  output [63:0] io_out_bits_data_3, // @[:@91750.4]
  output [63:0] io_out_bits_data_4, // @[:@91750.4]
  output [63:0] io_out_bits_data_5, // @[:@91750.4]
  output [63:0] io_out_bits_data_6, // @[:@91750.4]
  output [63:0] io_out_bits_data_7, // @[:@91750.4]
  output [63:0] io_out_bits_strobe // @[:@91750.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_in_bits_1; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_in_bits_2; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_in_bits_3; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_in_bits_4; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_in_bits_5; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_in_bits_6; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_in_bits_7; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_in_bits_8; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_in_bits_9; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_in_bits_10; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_in_bits_11; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_in_bits_12; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_in_bits_13; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_in_bits_14; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_in_bits_15; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_out_bits_1; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_out_bits_2; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_out_bits_3; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_out_bits_4; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_out_bits_5; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_out_bits_6; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_out_bits_7; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_out_bits_8; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_out_bits_9; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_out_bits_10; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_out_bits_11; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_out_bits_12; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_out_bits_13; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_out_bits_14; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire [31:0] FIFOVec_io_out_bits_15; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire  FIFOVec_io_chainEnq; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire  FIFOVec_io_chainDeq; // @[FIFOWidthConvert.scala 61:22:@91752.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_in_bits_0; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_ready; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_valid; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_bits_0; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_bits_1; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_bits_2; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_bits_3; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_bits_4; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_bits_5; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_bits_6; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_bits_7; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_bits_8; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_bits_9; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_bits_10; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_bits_11; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_bits_12; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_bits_13; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_bits_14; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire  FIFOVec_1_io_out_bits_15; // @[FIFOWidthConvert.scala 62:26:@91793.4]
  wire [319:0] _T_55; // @[Cat.scala 30:58:@91852.4]
  wire [511:0] _T_61; // @[Cat.scala 30:58:@91858.4]
  wire [9:0] _T_92; // @[Cat.scala 30:58:@91892.4]
  wire [15:0] _T_98; // @[Cat.scala 30:58:@91898.4]
  wire  _T_99; // @[FIFOWidthConvert.scala 36:14:@91899.4]
  wire  _T_103; // @[FIFOWidthConvert.scala 36:14:@91903.4]
  wire  _T_107; // @[FIFOWidthConvert.scala 36:14:@91907.4]
  wire  _T_111; // @[FIFOWidthConvert.scala 36:14:@91911.4]
  wire  _T_115; // @[FIFOWidthConvert.scala 36:14:@91915.4]
  wire  _T_119; // @[FIFOWidthConvert.scala 36:14:@91919.4]
  wire  _T_123; // @[FIFOWidthConvert.scala 36:14:@91923.4]
  wire  _T_127; // @[FIFOWidthConvert.scala 36:14:@91927.4]
  wire  _T_131; // @[FIFOWidthConvert.scala 36:14:@91931.4]
  wire  _T_135; // @[FIFOWidthConvert.scala 36:14:@91935.4]
  wire  _T_139; // @[FIFOWidthConvert.scala 36:14:@91939.4]
  wire  _T_143; // @[FIFOWidthConvert.scala 36:14:@91943.4]
  wire  _T_147; // @[FIFOWidthConvert.scala 36:14:@91947.4]
  wire  _T_151; // @[FIFOWidthConvert.scala 36:14:@91951.4]
  wire  _T_155; // @[FIFOWidthConvert.scala 36:14:@91955.4]
  wire  _T_159; // @[FIFOWidthConvert.scala 36:14:@91959.4]
  wire [9:0] _T_241; // @[Cat.scala 30:58:@92036.4]
  wire [18:0] _T_250; // @[Cat.scala 30:58:@92045.4]
  wire [27:0] _T_259; // @[Cat.scala 30:58:@92054.4]
  wire [36:0] _T_268; // @[Cat.scala 30:58:@92063.4]
  wire [45:0] _T_277; // @[Cat.scala 30:58:@92072.4]
  wire [54:0] _T_286; // @[Cat.scala 30:58:@92081.4]
  wire [62:0] _T_294; // @[Cat.scala 30:58:@92089.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 61:22:@91752.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_in_bits_1(FIFOVec_io_in_bits_1),
    .io_in_bits_2(FIFOVec_io_in_bits_2),
    .io_in_bits_3(FIFOVec_io_in_bits_3),
    .io_in_bits_4(FIFOVec_io_in_bits_4),
    .io_in_bits_5(FIFOVec_io_in_bits_5),
    .io_in_bits_6(FIFOVec_io_in_bits_6),
    .io_in_bits_7(FIFOVec_io_in_bits_7),
    .io_in_bits_8(FIFOVec_io_in_bits_8),
    .io_in_bits_9(FIFOVec_io_in_bits_9),
    .io_in_bits_10(FIFOVec_io_in_bits_10),
    .io_in_bits_11(FIFOVec_io_in_bits_11),
    .io_in_bits_12(FIFOVec_io_in_bits_12),
    .io_in_bits_13(FIFOVec_io_in_bits_13),
    .io_in_bits_14(FIFOVec_io_in_bits_14),
    .io_in_bits_15(FIFOVec_io_in_bits_15),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0),
    .io_out_bits_1(FIFOVec_io_out_bits_1),
    .io_out_bits_2(FIFOVec_io_out_bits_2),
    .io_out_bits_3(FIFOVec_io_out_bits_3),
    .io_out_bits_4(FIFOVec_io_out_bits_4),
    .io_out_bits_5(FIFOVec_io_out_bits_5),
    .io_out_bits_6(FIFOVec_io_out_bits_6),
    .io_out_bits_7(FIFOVec_io_out_bits_7),
    .io_out_bits_8(FIFOVec_io_out_bits_8),
    .io_out_bits_9(FIFOVec_io_out_bits_9),
    .io_out_bits_10(FIFOVec_io_out_bits_10),
    .io_out_bits_11(FIFOVec_io_out_bits_11),
    .io_out_bits_12(FIFOVec_io_out_bits_12),
    .io_out_bits_13(FIFOVec_io_out_bits_13),
    .io_out_bits_14(FIFOVec_io_out_bits_14),
    .io_out_bits_15(FIFOVec_io_out_bits_15),
    .io_chainEnq(FIFOVec_io_chainEnq),
    .io_chainDeq(FIFOVec_io_chainDeq)
  );
  FIFOVec_3 FIFOVec_1 ( // @[FIFOWidthConvert.scala 62:26:@91793.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid),
    .io_in_bits_0(FIFOVec_1_io_in_bits_0),
    .io_out_ready(FIFOVec_1_io_out_ready),
    .io_out_valid(FIFOVec_1_io_out_valid),
    .io_out_bits_0(FIFOVec_1_io_out_bits_0),
    .io_out_bits_1(FIFOVec_1_io_out_bits_1),
    .io_out_bits_2(FIFOVec_1_io_out_bits_2),
    .io_out_bits_3(FIFOVec_1_io_out_bits_3),
    .io_out_bits_4(FIFOVec_1_io_out_bits_4),
    .io_out_bits_5(FIFOVec_1_io_out_bits_5),
    .io_out_bits_6(FIFOVec_1_io_out_bits_6),
    .io_out_bits_7(FIFOVec_1_io_out_bits_7),
    .io_out_bits_8(FIFOVec_1_io_out_bits_8),
    .io_out_bits_9(FIFOVec_1_io_out_bits_9),
    .io_out_bits_10(FIFOVec_1_io_out_bits_10),
    .io_out_bits_11(FIFOVec_1_io_out_bits_11),
    .io_out_bits_12(FIFOVec_1_io_out_bits_12),
    .io_out_bits_13(FIFOVec_1_io_out_bits_13),
    .io_out_bits_14(FIFOVec_1_io_out_bits_14),
    .io_out_bits_15(FIFOVec_1_io_out_bits_15)
  );
  assign _T_55 = {FIFOVec_io_out_bits_15,FIFOVec_io_out_bits_14,FIFOVec_io_out_bits_13,FIFOVec_io_out_bits_12,FIFOVec_io_out_bits_11,FIFOVec_io_out_bits_10,FIFOVec_io_out_bits_9,FIFOVec_io_out_bits_8,FIFOVec_io_out_bits_7,FIFOVec_io_out_bits_6}; // @[Cat.scala 30:58:@91852.4]
  assign _T_61 = {_T_55,FIFOVec_io_out_bits_5,FIFOVec_io_out_bits_4,FIFOVec_io_out_bits_3,FIFOVec_io_out_bits_2,FIFOVec_io_out_bits_1,FIFOVec_io_out_bits_0}; // @[Cat.scala 30:58:@91858.4]
  assign _T_92 = {FIFOVec_1_io_out_bits_0,FIFOVec_1_io_out_bits_1,FIFOVec_1_io_out_bits_2,FIFOVec_1_io_out_bits_3,FIFOVec_1_io_out_bits_4,FIFOVec_1_io_out_bits_5,FIFOVec_1_io_out_bits_6,FIFOVec_1_io_out_bits_7,FIFOVec_1_io_out_bits_8,FIFOVec_1_io_out_bits_9}; // @[Cat.scala 30:58:@91892.4]
  assign _T_98 = {_T_92,FIFOVec_1_io_out_bits_10,FIFOVec_1_io_out_bits_11,FIFOVec_1_io_out_bits_12,FIFOVec_1_io_out_bits_13,FIFOVec_1_io_out_bits_14,FIFOVec_1_io_out_bits_15}; // @[Cat.scala 30:58:@91898.4]
  assign _T_99 = _T_98[0]; // @[FIFOWidthConvert.scala 36:14:@91899.4]
  assign _T_103 = _T_98[1]; // @[FIFOWidthConvert.scala 36:14:@91903.4]
  assign _T_107 = _T_98[2]; // @[FIFOWidthConvert.scala 36:14:@91907.4]
  assign _T_111 = _T_98[3]; // @[FIFOWidthConvert.scala 36:14:@91911.4]
  assign _T_115 = _T_98[4]; // @[FIFOWidthConvert.scala 36:14:@91915.4]
  assign _T_119 = _T_98[5]; // @[FIFOWidthConvert.scala 36:14:@91919.4]
  assign _T_123 = _T_98[6]; // @[FIFOWidthConvert.scala 36:14:@91923.4]
  assign _T_127 = _T_98[7]; // @[FIFOWidthConvert.scala 36:14:@91927.4]
  assign _T_131 = _T_98[8]; // @[FIFOWidthConvert.scala 36:14:@91931.4]
  assign _T_135 = _T_98[9]; // @[FIFOWidthConvert.scala 36:14:@91935.4]
  assign _T_139 = _T_98[10]; // @[FIFOWidthConvert.scala 36:14:@91939.4]
  assign _T_143 = _T_98[11]; // @[FIFOWidthConvert.scala 36:14:@91943.4]
  assign _T_147 = _T_98[12]; // @[FIFOWidthConvert.scala 36:14:@91947.4]
  assign _T_151 = _T_98[13]; // @[FIFOWidthConvert.scala 36:14:@91951.4]
  assign _T_155 = _T_98[14]; // @[FIFOWidthConvert.scala 36:14:@91955.4]
  assign _T_159 = _T_98[15]; // @[FIFOWidthConvert.scala 36:14:@91959.4]
  assign _T_241 = {_T_159,_T_159,_T_159,_T_159,_T_155,_T_155,_T_155,_T_155,_T_151,_T_151}; // @[Cat.scala 30:58:@92036.4]
  assign _T_250 = {_T_241,_T_151,_T_151,_T_147,_T_147,_T_147,_T_147,_T_143,_T_143,_T_143}; // @[Cat.scala 30:58:@92045.4]
  assign _T_259 = {_T_250,_T_143,_T_139,_T_139,_T_139,_T_139,_T_135,_T_135,_T_135,_T_135}; // @[Cat.scala 30:58:@92054.4]
  assign _T_268 = {_T_259,_T_131,_T_131,_T_131,_T_131,_T_127,_T_127,_T_127,_T_127,_T_123}; // @[Cat.scala 30:58:@92063.4]
  assign _T_277 = {_T_268,_T_123,_T_123,_T_123,_T_119,_T_119,_T_119,_T_119,_T_115,_T_115}; // @[Cat.scala 30:58:@92072.4]
  assign _T_286 = {_T_277,_T_115,_T_115,_T_111,_T_111,_T_111,_T_111,_T_107,_T_107,_T_107}; // @[Cat.scala 30:58:@92081.4]
  assign _T_294 = {_T_286,_T_107,_T_103,_T_103,_T_103,_T_103,_T_99,_T_99,_T_99}; // @[Cat.scala 30:58:@92089.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 71:17:@91842.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 72:18:@91843.4]
  assign io_out_bits_data_0 = _T_61[63:0]; // @[FIFOWidthConvert.scala 73:22:@91876.4]
  assign io_out_bits_data_1 = _T_61[127:64]; // @[FIFOWidthConvert.scala 73:22:@91877.4]
  assign io_out_bits_data_2 = _T_61[191:128]; // @[FIFOWidthConvert.scala 73:22:@91878.4]
  assign io_out_bits_data_3 = _T_61[255:192]; // @[FIFOWidthConvert.scala 73:22:@91879.4]
  assign io_out_bits_data_4 = _T_61[319:256]; // @[FIFOWidthConvert.scala 73:22:@91880.4]
  assign io_out_bits_data_5 = _T_61[383:320]; // @[FIFOWidthConvert.scala 73:22:@91881.4]
  assign io_out_bits_data_6 = _T_61[447:384]; // @[FIFOWidthConvert.scala 73:22:@91882.4]
  assign io_out_bits_data_7 = _T_61[511:448]; // @[FIFOWidthConvert.scala 73:22:@91883.4]
  assign io_out_bits_strobe = {_T_294,_T_99}; // @[FIFOWidthConvert.scala 74:24:@92091.4]
  assign FIFOVec_clock = clock; // @[:@91753.4]
  assign FIFOVec_reset = reset; // @[:@91754.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 68:22:@91839.4]
  assign FIFOVec_io_in_bits_0 = io_in_bits_data_0; // @[FIFOWidthConvert.scala 67:24:@91838.4]
  assign FIFOVec_io_in_bits_1 = 32'h0;
  assign FIFOVec_io_in_bits_2 = 32'h0;
  assign FIFOVec_io_in_bits_3 = 32'h0;
  assign FIFOVec_io_in_bits_4 = 32'h0;
  assign FIFOVec_io_in_bits_5 = 32'h0;
  assign FIFOVec_io_in_bits_6 = 32'h0;
  assign FIFOVec_io_in_bits_7 = 32'h0;
  assign FIFOVec_io_in_bits_8 = 32'h0;
  assign FIFOVec_io_in_bits_9 = 32'h0;
  assign FIFOVec_io_in_bits_10 = 32'h0;
  assign FIFOVec_io_in_bits_11 = 32'h0;
  assign FIFOVec_io_in_bits_12 = 32'h0;
  assign FIFOVec_io_in_bits_13 = 32'h0;
  assign FIFOVec_io_in_bits_14 = 32'h0;
  assign FIFOVec_io_in_bits_15 = 32'h0;
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 75:23:@92092.4]
  assign FIFOVec_io_chainEnq = 1'h1; // @[FIFOWidthConvert.scala 63:22:@91834.4]
  assign FIFOVec_io_chainDeq = 1'h0; // @[FIFOWidthConvert.scala 64:22:@91835.4]
  assign FIFOVec_1_clock = clock; // @[:@91794.4]
  assign FIFOVec_1_reset = reset; // @[:@91795.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 70:26:@91841.4]
  assign FIFOVec_1_io_in_bits_0 = io_in_bits_strobe; // @[FIFOWidthConvert.scala 69:28:@91840.4]
  assign FIFOVec_1_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 76:27:@92093.4]
endmodule
module FFRAM_16( // @[:@92131.2]
  input        clock, // @[:@92132.4]
  input        reset, // @[:@92133.4]
  input  [5:0] io_raddr, // @[:@92134.4]
  input        io_wen, // @[:@92134.4]
  input  [5:0] io_waddr, // @[:@92134.4]
  output       io_rdata // @[:@92134.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@92138.4]
  reg [31:0] _RAND_0;
  wire  _T_688; // @[SRAM.scala 148:37:@92139.4]
  wire  _T_689; // @[SRAM.scala 148:25:@92140.4]
  wire  _GEN_0; // @[SRAM.scala 148:48:@92142.4]
  reg  regs_1; // @[SRAM.scala 145:20:@92149.4]
  reg [31:0] _RAND_1;
  wire  _T_697; // @[SRAM.scala 148:37:@92150.4]
  wire  _T_698; // @[SRAM.scala 148:25:@92151.4]
  wire  _GEN_1; // @[SRAM.scala 148:48:@92153.4]
  reg  regs_2; // @[SRAM.scala 145:20:@92160.4]
  reg [31:0] _RAND_2;
  wire  _T_706; // @[SRAM.scala 148:37:@92161.4]
  wire  _T_707; // @[SRAM.scala 148:25:@92162.4]
  wire  _GEN_2; // @[SRAM.scala 148:48:@92164.4]
  reg  regs_3; // @[SRAM.scala 145:20:@92171.4]
  reg [31:0] _RAND_3;
  wire  _T_715; // @[SRAM.scala 148:37:@92172.4]
  wire  _T_716; // @[SRAM.scala 148:25:@92173.4]
  wire  _GEN_3; // @[SRAM.scala 148:48:@92175.4]
  reg  regs_4; // @[SRAM.scala 145:20:@92182.4]
  reg [31:0] _RAND_4;
  wire  _T_724; // @[SRAM.scala 148:37:@92183.4]
  wire  _T_725; // @[SRAM.scala 148:25:@92184.4]
  wire  _GEN_4; // @[SRAM.scala 148:48:@92186.4]
  reg  regs_5; // @[SRAM.scala 145:20:@92193.4]
  reg [31:0] _RAND_5;
  wire  _T_733; // @[SRAM.scala 148:37:@92194.4]
  wire  _T_734; // @[SRAM.scala 148:25:@92195.4]
  wire  _GEN_5; // @[SRAM.scala 148:48:@92197.4]
  reg  regs_6; // @[SRAM.scala 145:20:@92204.4]
  reg [31:0] _RAND_6;
  wire  _T_742; // @[SRAM.scala 148:37:@92205.4]
  wire  _T_743; // @[SRAM.scala 148:25:@92206.4]
  wire  _GEN_6; // @[SRAM.scala 148:48:@92208.4]
  reg  regs_7; // @[SRAM.scala 145:20:@92215.4]
  reg [31:0] _RAND_7;
  wire  _T_751; // @[SRAM.scala 148:37:@92216.4]
  wire  _T_752; // @[SRAM.scala 148:25:@92217.4]
  wire  _GEN_7; // @[SRAM.scala 148:48:@92219.4]
  reg  regs_8; // @[SRAM.scala 145:20:@92226.4]
  reg [31:0] _RAND_8;
  wire  _T_760; // @[SRAM.scala 148:37:@92227.4]
  wire  _T_761; // @[SRAM.scala 148:25:@92228.4]
  wire  _GEN_8; // @[SRAM.scala 148:48:@92230.4]
  reg  regs_9; // @[SRAM.scala 145:20:@92237.4]
  reg [31:0] _RAND_9;
  wire  _T_769; // @[SRAM.scala 148:37:@92238.4]
  wire  _T_770; // @[SRAM.scala 148:25:@92239.4]
  wire  _GEN_9; // @[SRAM.scala 148:48:@92241.4]
  reg  regs_10; // @[SRAM.scala 145:20:@92248.4]
  reg [31:0] _RAND_10;
  wire  _T_778; // @[SRAM.scala 148:37:@92249.4]
  wire  _T_779; // @[SRAM.scala 148:25:@92250.4]
  wire  _GEN_10; // @[SRAM.scala 148:48:@92252.4]
  reg  regs_11; // @[SRAM.scala 145:20:@92259.4]
  reg [31:0] _RAND_11;
  wire  _T_787; // @[SRAM.scala 148:37:@92260.4]
  wire  _T_788; // @[SRAM.scala 148:25:@92261.4]
  wire  _GEN_11; // @[SRAM.scala 148:48:@92263.4]
  reg  regs_12; // @[SRAM.scala 145:20:@92270.4]
  reg [31:0] _RAND_12;
  wire  _T_796; // @[SRAM.scala 148:37:@92271.4]
  wire  _T_797; // @[SRAM.scala 148:25:@92272.4]
  wire  _GEN_12; // @[SRAM.scala 148:48:@92274.4]
  reg  regs_13; // @[SRAM.scala 145:20:@92281.4]
  reg [31:0] _RAND_13;
  wire  _T_805; // @[SRAM.scala 148:37:@92282.4]
  wire  _T_806; // @[SRAM.scala 148:25:@92283.4]
  wire  _GEN_13; // @[SRAM.scala 148:48:@92285.4]
  reg  regs_14; // @[SRAM.scala 145:20:@92292.4]
  reg [31:0] _RAND_14;
  wire  _T_814; // @[SRAM.scala 148:37:@92293.4]
  wire  _T_815; // @[SRAM.scala 148:25:@92294.4]
  wire  _GEN_14; // @[SRAM.scala 148:48:@92296.4]
  reg  regs_15; // @[SRAM.scala 145:20:@92303.4]
  reg [31:0] _RAND_15;
  wire  _T_823; // @[SRAM.scala 148:37:@92304.4]
  wire  _T_824; // @[SRAM.scala 148:25:@92305.4]
  wire  _GEN_15; // @[SRAM.scala 148:48:@92307.4]
  reg  regs_16; // @[SRAM.scala 145:20:@92314.4]
  reg [31:0] _RAND_16;
  wire  _T_832; // @[SRAM.scala 148:37:@92315.4]
  wire  _T_833; // @[SRAM.scala 148:25:@92316.4]
  wire  _GEN_16; // @[SRAM.scala 148:48:@92318.4]
  reg  regs_17; // @[SRAM.scala 145:20:@92325.4]
  reg [31:0] _RAND_17;
  wire  _T_841; // @[SRAM.scala 148:37:@92326.4]
  wire  _T_842; // @[SRAM.scala 148:25:@92327.4]
  wire  _GEN_17; // @[SRAM.scala 148:48:@92329.4]
  reg  regs_18; // @[SRAM.scala 145:20:@92336.4]
  reg [31:0] _RAND_18;
  wire  _T_850; // @[SRAM.scala 148:37:@92337.4]
  wire  _T_851; // @[SRAM.scala 148:25:@92338.4]
  wire  _GEN_18; // @[SRAM.scala 148:48:@92340.4]
  reg  regs_19; // @[SRAM.scala 145:20:@92347.4]
  reg [31:0] _RAND_19;
  wire  _T_859; // @[SRAM.scala 148:37:@92348.4]
  wire  _T_860; // @[SRAM.scala 148:25:@92349.4]
  wire  _GEN_19; // @[SRAM.scala 148:48:@92351.4]
  reg  regs_20; // @[SRAM.scala 145:20:@92358.4]
  reg [31:0] _RAND_20;
  wire  _T_868; // @[SRAM.scala 148:37:@92359.4]
  wire  _T_869; // @[SRAM.scala 148:25:@92360.4]
  wire  _GEN_20; // @[SRAM.scala 148:48:@92362.4]
  reg  regs_21; // @[SRAM.scala 145:20:@92369.4]
  reg [31:0] _RAND_21;
  wire  _T_877; // @[SRAM.scala 148:37:@92370.4]
  wire  _T_878; // @[SRAM.scala 148:25:@92371.4]
  wire  _GEN_21; // @[SRAM.scala 148:48:@92373.4]
  reg  regs_22; // @[SRAM.scala 145:20:@92380.4]
  reg [31:0] _RAND_22;
  wire  _T_886; // @[SRAM.scala 148:37:@92381.4]
  wire  _T_887; // @[SRAM.scala 148:25:@92382.4]
  wire  _GEN_22; // @[SRAM.scala 148:48:@92384.4]
  reg  regs_23; // @[SRAM.scala 145:20:@92391.4]
  reg [31:0] _RAND_23;
  wire  _T_895; // @[SRAM.scala 148:37:@92392.4]
  wire  _T_896; // @[SRAM.scala 148:25:@92393.4]
  wire  _GEN_23; // @[SRAM.scala 148:48:@92395.4]
  reg  regs_24; // @[SRAM.scala 145:20:@92402.4]
  reg [31:0] _RAND_24;
  wire  _T_904; // @[SRAM.scala 148:37:@92403.4]
  wire  _T_905; // @[SRAM.scala 148:25:@92404.4]
  wire  _GEN_24; // @[SRAM.scala 148:48:@92406.4]
  reg  regs_25; // @[SRAM.scala 145:20:@92413.4]
  reg [31:0] _RAND_25;
  wire  _T_913; // @[SRAM.scala 148:37:@92414.4]
  wire  _T_914; // @[SRAM.scala 148:25:@92415.4]
  wire  _GEN_25; // @[SRAM.scala 148:48:@92417.4]
  reg  regs_26; // @[SRAM.scala 145:20:@92424.4]
  reg [31:0] _RAND_26;
  wire  _T_922; // @[SRAM.scala 148:37:@92425.4]
  wire  _T_923; // @[SRAM.scala 148:25:@92426.4]
  wire  _GEN_26; // @[SRAM.scala 148:48:@92428.4]
  reg  regs_27; // @[SRAM.scala 145:20:@92435.4]
  reg [31:0] _RAND_27;
  wire  _T_931; // @[SRAM.scala 148:37:@92436.4]
  wire  _T_932; // @[SRAM.scala 148:25:@92437.4]
  wire  _GEN_27; // @[SRAM.scala 148:48:@92439.4]
  reg  regs_28; // @[SRAM.scala 145:20:@92446.4]
  reg [31:0] _RAND_28;
  wire  _T_940; // @[SRAM.scala 148:37:@92447.4]
  wire  _T_941; // @[SRAM.scala 148:25:@92448.4]
  wire  _GEN_28; // @[SRAM.scala 148:48:@92450.4]
  reg  regs_29; // @[SRAM.scala 145:20:@92457.4]
  reg [31:0] _RAND_29;
  wire  _T_949; // @[SRAM.scala 148:37:@92458.4]
  wire  _T_950; // @[SRAM.scala 148:25:@92459.4]
  wire  _GEN_29; // @[SRAM.scala 148:48:@92461.4]
  reg  regs_30; // @[SRAM.scala 145:20:@92468.4]
  reg [31:0] _RAND_30;
  wire  _T_958; // @[SRAM.scala 148:37:@92469.4]
  wire  _T_959; // @[SRAM.scala 148:25:@92470.4]
  wire  _GEN_30; // @[SRAM.scala 148:48:@92472.4]
  reg  regs_31; // @[SRAM.scala 145:20:@92479.4]
  reg [31:0] _RAND_31;
  wire  _T_967; // @[SRAM.scala 148:37:@92480.4]
  wire  _T_968; // @[SRAM.scala 148:25:@92481.4]
  wire  _GEN_31; // @[SRAM.scala 148:48:@92483.4]
  reg  regs_32; // @[SRAM.scala 145:20:@92490.4]
  reg [31:0] _RAND_32;
  wire  _T_976; // @[SRAM.scala 148:37:@92491.4]
  wire  _T_977; // @[SRAM.scala 148:25:@92492.4]
  wire  _GEN_32; // @[SRAM.scala 148:48:@92494.4]
  reg  regs_33; // @[SRAM.scala 145:20:@92501.4]
  reg [31:0] _RAND_33;
  wire  _T_985; // @[SRAM.scala 148:37:@92502.4]
  wire  _T_986; // @[SRAM.scala 148:25:@92503.4]
  wire  _GEN_33; // @[SRAM.scala 148:48:@92505.4]
  reg  regs_34; // @[SRAM.scala 145:20:@92512.4]
  reg [31:0] _RAND_34;
  wire  _T_994; // @[SRAM.scala 148:37:@92513.4]
  wire  _T_995; // @[SRAM.scala 148:25:@92514.4]
  wire  _GEN_34; // @[SRAM.scala 148:48:@92516.4]
  reg  regs_35; // @[SRAM.scala 145:20:@92523.4]
  reg [31:0] _RAND_35;
  wire  _T_1003; // @[SRAM.scala 148:37:@92524.4]
  wire  _T_1004; // @[SRAM.scala 148:25:@92525.4]
  wire  _GEN_35; // @[SRAM.scala 148:48:@92527.4]
  reg  regs_36; // @[SRAM.scala 145:20:@92534.4]
  reg [31:0] _RAND_36;
  wire  _T_1012; // @[SRAM.scala 148:37:@92535.4]
  wire  _T_1013; // @[SRAM.scala 148:25:@92536.4]
  wire  _GEN_36; // @[SRAM.scala 148:48:@92538.4]
  reg  regs_37; // @[SRAM.scala 145:20:@92545.4]
  reg [31:0] _RAND_37;
  wire  _T_1021; // @[SRAM.scala 148:37:@92546.4]
  wire  _T_1022; // @[SRAM.scala 148:25:@92547.4]
  wire  _GEN_37; // @[SRAM.scala 148:48:@92549.4]
  reg  regs_38; // @[SRAM.scala 145:20:@92556.4]
  reg [31:0] _RAND_38;
  wire  _T_1030; // @[SRAM.scala 148:37:@92557.4]
  wire  _T_1031; // @[SRAM.scala 148:25:@92558.4]
  wire  _GEN_38; // @[SRAM.scala 148:48:@92560.4]
  reg  regs_39; // @[SRAM.scala 145:20:@92567.4]
  reg [31:0] _RAND_39;
  wire  _T_1039; // @[SRAM.scala 148:37:@92568.4]
  wire  _T_1040; // @[SRAM.scala 148:25:@92569.4]
  wire  _GEN_39; // @[SRAM.scala 148:48:@92571.4]
  reg  regs_40; // @[SRAM.scala 145:20:@92578.4]
  reg [31:0] _RAND_40;
  wire  _T_1048; // @[SRAM.scala 148:37:@92579.4]
  wire  _T_1049; // @[SRAM.scala 148:25:@92580.4]
  wire  _GEN_40; // @[SRAM.scala 148:48:@92582.4]
  reg  regs_41; // @[SRAM.scala 145:20:@92589.4]
  reg [31:0] _RAND_41;
  wire  _T_1057; // @[SRAM.scala 148:37:@92590.4]
  wire  _T_1058; // @[SRAM.scala 148:25:@92591.4]
  wire  _GEN_41; // @[SRAM.scala 148:48:@92593.4]
  reg  regs_42; // @[SRAM.scala 145:20:@92600.4]
  reg [31:0] _RAND_42;
  wire  _T_1066; // @[SRAM.scala 148:37:@92601.4]
  wire  _T_1067; // @[SRAM.scala 148:25:@92602.4]
  wire  _GEN_42; // @[SRAM.scala 148:48:@92604.4]
  reg  regs_43; // @[SRAM.scala 145:20:@92611.4]
  reg [31:0] _RAND_43;
  wire  _T_1075; // @[SRAM.scala 148:37:@92612.4]
  wire  _T_1076; // @[SRAM.scala 148:25:@92613.4]
  wire  _GEN_43; // @[SRAM.scala 148:48:@92615.4]
  reg  regs_44; // @[SRAM.scala 145:20:@92622.4]
  reg [31:0] _RAND_44;
  wire  _T_1084; // @[SRAM.scala 148:37:@92623.4]
  wire  _T_1085; // @[SRAM.scala 148:25:@92624.4]
  wire  _GEN_44; // @[SRAM.scala 148:48:@92626.4]
  reg  regs_45; // @[SRAM.scala 145:20:@92633.4]
  reg [31:0] _RAND_45;
  wire  _T_1093; // @[SRAM.scala 148:37:@92634.4]
  wire  _T_1094; // @[SRAM.scala 148:25:@92635.4]
  wire  _GEN_45; // @[SRAM.scala 148:48:@92637.4]
  reg  regs_46; // @[SRAM.scala 145:20:@92644.4]
  reg [31:0] _RAND_46;
  wire  _T_1102; // @[SRAM.scala 148:37:@92645.4]
  wire  _T_1103; // @[SRAM.scala 148:25:@92646.4]
  wire  _GEN_46; // @[SRAM.scala 148:48:@92648.4]
  reg  regs_47; // @[SRAM.scala 145:20:@92655.4]
  reg [31:0] _RAND_47;
  wire  _T_1111; // @[SRAM.scala 148:37:@92656.4]
  wire  _T_1112; // @[SRAM.scala 148:25:@92657.4]
  wire  _GEN_47; // @[SRAM.scala 148:48:@92659.4]
  reg  regs_48; // @[SRAM.scala 145:20:@92666.4]
  reg [31:0] _RAND_48;
  wire  _T_1120; // @[SRAM.scala 148:37:@92667.4]
  wire  _T_1121; // @[SRAM.scala 148:25:@92668.4]
  wire  _GEN_48; // @[SRAM.scala 148:48:@92670.4]
  reg  regs_49; // @[SRAM.scala 145:20:@92677.4]
  reg [31:0] _RAND_49;
  wire  _T_1129; // @[SRAM.scala 148:37:@92678.4]
  wire  _T_1130; // @[SRAM.scala 148:25:@92679.4]
  wire  _GEN_49; // @[SRAM.scala 148:48:@92681.4]
  reg  regs_50; // @[SRAM.scala 145:20:@92688.4]
  reg [31:0] _RAND_50;
  wire  _T_1138; // @[SRAM.scala 148:37:@92689.4]
  wire  _T_1139; // @[SRAM.scala 148:25:@92690.4]
  wire  _GEN_50; // @[SRAM.scala 148:48:@92692.4]
  reg  regs_51; // @[SRAM.scala 145:20:@92699.4]
  reg [31:0] _RAND_51;
  wire  _T_1147; // @[SRAM.scala 148:37:@92700.4]
  wire  _T_1148; // @[SRAM.scala 148:25:@92701.4]
  wire  _GEN_51; // @[SRAM.scala 148:48:@92703.4]
  reg  regs_52; // @[SRAM.scala 145:20:@92710.4]
  reg [31:0] _RAND_52;
  wire  _T_1156; // @[SRAM.scala 148:37:@92711.4]
  wire  _T_1157; // @[SRAM.scala 148:25:@92712.4]
  wire  _GEN_52; // @[SRAM.scala 148:48:@92714.4]
  reg  regs_53; // @[SRAM.scala 145:20:@92721.4]
  reg [31:0] _RAND_53;
  wire  _T_1165; // @[SRAM.scala 148:37:@92722.4]
  wire  _T_1166; // @[SRAM.scala 148:25:@92723.4]
  wire  _GEN_53; // @[SRAM.scala 148:48:@92725.4]
  reg  regs_54; // @[SRAM.scala 145:20:@92732.4]
  reg [31:0] _RAND_54;
  wire  _T_1174; // @[SRAM.scala 148:37:@92733.4]
  wire  _T_1175; // @[SRAM.scala 148:25:@92734.4]
  wire  _GEN_54; // @[SRAM.scala 148:48:@92736.4]
  reg  regs_55; // @[SRAM.scala 145:20:@92743.4]
  reg [31:0] _RAND_55;
  wire  _T_1183; // @[SRAM.scala 148:37:@92744.4]
  wire  _T_1184; // @[SRAM.scala 148:25:@92745.4]
  wire  _GEN_55; // @[SRAM.scala 148:48:@92747.4]
  reg  regs_56; // @[SRAM.scala 145:20:@92754.4]
  reg [31:0] _RAND_56;
  wire  _T_1192; // @[SRAM.scala 148:37:@92755.4]
  wire  _T_1193; // @[SRAM.scala 148:25:@92756.4]
  wire  _GEN_56; // @[SRAM.scala 148:48:@92758.4]
  reg  regs_57; // @[SRAM.scala 145:20:@92765.4]
  reg [31:0] _RAND_57;
  wire  _T_1201; // @[SRAM.scala 148:37:@92766.4]
  wire  _T_1202; // @[SRAM.scala 148:25:@92767.4]
  wire  _GEN_57; // @[SRAM.scala 148:48:@92769.4]
  reg  regs_58; // @[SRAM.scala 145:20:@92776.4]
  reg [31:0] _RAND_58;
  wire  _T_1210; // @[SRAM.scala 148:37:@92777.4]
  wire  _T_1211; // @[SRAM.scala 148:25:@92778.4]
  wire  _GEN_58; // @[SRAM.scala 148:48:@92780.4]
  reg  regs_59; // @[SRAM.scala 145:20:@92787.4]
  reg [31:0] _RAND_59;
  wire  _T_1219; // @[SRAM.scala 148:37:@92788.4]
  wire  _T_1220; // @[SRAM.scala 148:25:@92789.4]
  wire  _GEN_59; // @[SRAM.scala 148:48:@92791.4]
  reg  regs_60; // @[SRAM.scala 145:20:@92798.4]
  reg [31:0] _RAND_60;
  wire  _T_1228; // @[SRAM.scala 148:37:@92799.4]
  wire  _T_1229; // @[SRAM.scala 148:25:@92800.4]
  wire  _GEN_60; // @[SRAM.scala 148:48:@92802.4]
  reg  regs_61; // @[SRAM.scala 145:20:@92809.4]
  reg [31:0] _RAND_61;
  wire  _T_1237; // @[SRAM.scala 148:37:@92810.4]
  wire  _T_1238; // @[SRAM.scala 148:25:@92811.4]
  wire  _GEN_61; // @[SRAM.scala 148:48:@92813.4]
  reg  regs_62; // @[SRAM.scala 145:20:@92820.4]
  reg [31:0] _RAND_62;
  wire  _T_1246; // @[SRAM.scala 148:37:@92821.4]
  wire  _T_1247; // @[SRAM.scala 148:25:@92822.4]
  wire  _GEN_62; // @[SRAM.scala 148:48:@92824.4]
  reg  regs_63; // @[SRAM.scala 145:20:@92831.4]
  reg [31:0] _RAND_63;
  wire  _T_1255; // @[SRAM.scala 148:37:@92832.4]
  wire  _T_1256; // @[SRAM.scala 148:25:@92833.4]
  wire  _GEN_63; // @[SRAM.scala 148:48:@92835.4]
  wire  _GEN_65; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_66; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_67; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_68; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_69; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_70; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_71; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_72; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_73; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_74; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_75; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_76; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_77; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_78; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_79; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_80; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_81; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_82; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_83; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_84; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_85; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_86; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_87; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_88; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_89; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_90; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_91; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_92; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_93; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_94; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_95; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_96; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_97; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_98; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_99; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_100; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_101; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_102; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_103; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_104; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_105; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_106; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_107; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_108; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_109; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_110; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_111; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_112; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_113; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_114; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_115; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_116; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_117; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_118; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_119; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_120; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_121; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_122; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_123; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_124; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_125; // @[SRAM.scala 155:12:@92905.4]
  wire  _GEN_126; // @[SRAM.scala 155:12:@92905.4]
  assign _T_688 = io_waddr == 6'h0; // @[SRAM.scala 148:37:@92139.4]
  assign _T_689 = io_wen & _T_688; // @[SRAM.scala 148:25:@92140.4]
  assign _GEN_0 = _T_689 ? 1'h1 : regs_0; // @[SRAM.scala 148:48:@92142.4]
  assign _T_697 = io_waddr == 6'h1; // @[SRAM.scala 148:37:@92150.4]
  assign _T_698 = io_wen & _T_697; // @[SRAM.scala 148:25:@92151.4]
  assign _GEN_1 = _T_698 ? 1'h1 : regs_1; // @[SRAM.scala 148:48:@92153.4]
  assign _T_706 = io_waddr == 6'h2; // @[SRAM.scala 148:37:@92161.4]
  assign _T_707 = io_wen & _T_706; // @[SRAM.scala 148:25:@92162.4]
  assign _GEN_2 = _T_707 ? 1'h1 : regs_2; // @[SRAM.scala 148:48:@92164.4]
  assign _T_715 = io_waddr == 6'h3; // @[SRAM.scala 148:37:@92172.4]
  assign _T_716 = io_wen & _T_715; // @[SRAM.scala 148:25:@92173.4]
  assign _GEN_3 = _T_716 ? 1'h1 : regs_3; // @[SRAM.scala 148:48:@92175.4]
  assign _T_724 = io_waddr == 6'h4; // @[SRAM.scala 148:37:@92183.4]
  assign _T_725 = io_wen & _T_724; // @[SRAM.scala 148:25:@92184.4]
  assign _GEN_4 = _T_725 ? 1'h1 : regs_4; // @[SRAM.scala 148:48:@92186.4]
  assign _T_733 = io_waddr == 6'h5; // @[SRAM.scala 148:37:@92194.4]
  assign _T_734 = io_wen & _T_733; // @[SRAM.scala 148:25:@92195.4]
  assign _GEN_5 = _T_734 ? 1'h1 : regs_5; // @[SRAM.scala 148:48:@92197.4]
  assign _T_742 = io_waddr == 6'h6; // @[SRAM.scala 148:37:@92205.4]
  assign _T_743 = io_wen & _T_742; // @[SRAM.scala 148:25:@92206.4]
  assign _GEN_6 = _T_743 ? 1'h1 : regs_6; // @[SRAM.scala 148:48:@92208.4]
  assign _T_751 = io_waddr == 6'h7; // @[SRAM.scala 148:37:@92216.4]
  assign _T_752 = io_wen & _T_751; // @[SRAM.scala 148:25:@92217.4]
  assign _GEN_7 = _T_752 ? 1'h1 : regs_7; // @[SRAM.scala 148:48:@92219.4]
  assign _T_760 = io_waddr == 6'h8; // @[SRAM.scala 148:37:@92227.4]
  assign _T_761 = io_wen & _T_760; // @[SRAM.scala 148:25:@92228.4]
  assign _GEN_8 = _T_761 ? 1'h1 : regs_8; // @[SRAM.scala 148:48:@92230.4]
  assign _T_769 = io_waddr == 6'h9; // @[SRAM.scala 148:37:@92238.4]
  assign _T_770 = io_wen & _T_769; // @[SRAM.scala 148:25:@92239.4]
  assign _GEN_9 = _T_770 ? 1'h1 : regs_9; // @[SRAM.scala 148:48:@92241.4]
  assign _T_778 = io_waddr == 6'ha; // @[SRAM.scala 148:37:@92249.4]
  assign _T_779 = io_wen & _T_778; // @[SRAM.scala 148:25:@92250.4]
  assign _GEN_10 = _T_779 ? 1'h1 : regs_10; // @[SRAM.scala 148:48:@92252.4]
  assign _T_787 = io_waddr == 6'hb; // @[SRAM.scala 148:37:@92260.4]
  assign _T_788 = io_wen & _T_787; // @[SRAM.scala 148:25:@92261.4]
  assign _GEN_11 = _T_788 ? 1'h1 : regs_11; // @[SRAM.scala 148:48:@92263.4]
  assign _T_796 = io_waddr == 6'hc; // @[SRAM.scala 148:37:@92271.4]
  assign _T_797 = io_wen & _T_796; // @[SRAM.scala 148:25:@92272.4]
  assign _GEN_12 = _T_797 ? 1'h1 : regs_12; // @[SRAM.scala 148:48:@92274.4]
  assign _T_805 = io_waddr == 6'hd; // @[SRAM.scala 148:37:@92282.4]
  assign _T_806 = io_wen & _T_805; // @[SRAM.scala 148:25:@92283.4]
  assign _GEN_13 = _T_806 ? 1'h1 : regs_13; // @[SRAM.scala 148:48:@92285.4]
  assign _T_814 = io_waddr == 6'he; // @[SRAM.scala 148:37:@92293.4]
  assign _T_815 = io_wen & _T_814; // @[SRAM.scala 148:25:@92294.4]
  assign _GEN_14 = _T_815 ? 1'h1 : regs_14; // @[SRAM.scala 148:48:@92296.4]
  assign _T_823 = io_waddr == 6'hf; // @[SRAM.scala 148:37:@92304.4]
  assign _T_824 = io_wen & _T_823; // @[SRAM.scala 148:25:@92305.4]
  assign _GEN_15 = _T_824 ? 1'h1 : regs_15; // @[SRAM.scala 148:48:@92307.4]
  assign _T_832 = io_waddr == 6'h10; // @[SRAM.scala 148:37:@92315.4]
  assign _T_833 = io_wen & _T_832; // @[SRAM.scala 148:25:@92316.4]
  assign _GEN_16 = _T_833 ? 1'h1 : regs_16; // @[SRAM.scala 148:48:@92318.4]
  assign _T_841 = io_waddr == 6'h11; // @[SRAM.scala 148:37:@92326.4]
  assign _T_842 = io_wen & _T_841; // @[SRAM.scala 148:25:@92327.4]
  assign _GEN_17 = _T_842 ? 1'h1 : regs_17; // @[SRAM.scala 148:48:@92329.4]
  assign _T_850 = io_waddr == 6'h12; // @[SRAM.scala 148:37:@92337.4]
  assign _T_851 = io_wen & _T_850; // @[SRAM.scala 148:25:@92338.4]
  assign _GEN_18 = _T_851 ? 1'h1 : regs_18; // @[SRAM.scala 148:48:@92340.4]
  assign _T_859 = io_waddr == 6'h13; // @[SRAM.scala 148:37:@92348.4]
  assign _T_860 = io_wen & _T_859; // @[SRAM.scala 148:25:@92349.4]
  assign _GEN_19 = _T_860 ? 1'h1 : regs_19; // @[SRAM.scala 148:48:@92351.4]
  assign _T_868 = io_waddr == 6'h14; // @[SRAM.scala 148:37:@92359.4]
  assign _T_869 = io_wen & _T_868; // @[SRAM.scala 148:25:@92360.4]
  assign _GEN_20 = _T_869 ? 1'h1 : regs_20; // @[SRAM.scala 148:48:@92362.4]
  assign _T_877 = io_waddr == 6'h15; // @[SRAM.scala 148:37:@92370.4]
  assign _T_878 = io_wen & _T_877; // @[SRAM.scala 148:25:@92371.4]
  assign _GEN_21 = _T_878 ? 1'h1 : regs_21; // @[SRAM.scala 148:48:@92373.4]
  assign _T_886 = io_waddr == 6'h16; // @[SRAM.scala 148:37:@92381.4]
  assign _T_887 = io_wen & _T_886; // @[SRAM.scala 148:25:@92382.4]
  assign _GEN_22 = _T_887 ? 1'h1 : regs_22; // @[SRAM.scala 148:48:@92384.4]
  assign _T_895 = io_waddr == 6'h17; // @[SRAM.scala 148:37:@92392.4]
  assign _T_896 = io_wen & _T_895; // @[SRAM.scala 148:25:@92393.4]
  assign _GEN_23 = _T_896 ? 1'h1 : regs_23; // @[SRAM.scala 148:48:@92395.4]
  assign _T_904 = io_waddr == 6'h18; // @[SRAM.scala 148:37:@92403.4]
  assign _T_905 = io_wen & _T_904; // @[SRAM.scala 148:25:@92404.4]
  assign _GEN_24 = _T_905 ? 1'h1 : regs_24; // @[SRAM.scala 148:48:@92406.4]
  assign _T_913 = io_waddr == 6'h19; // @[SRAM.scala 148:37:@92414.4]
  assign _T_914 = io_wen & _T_913; // @[SRAM.scala 148:25:@92415.4]
  assign _GEN_25 = _T_914 ? 1'h1 : regs_25; // @[SRAM.scala 148:48:@92417.4]
  assign _T_922 = io_waddr == 6'h1a; // @[SRAM.scala 148:37:@92425.4]
  assign _T_923 = io_wen & _T_922; // @[SRAM.scala 148:25:@92426.4]
  assign _GEN_26 = _T_923 ? 1'h1 : regs_26; // @[SRAM.scala 148:48:@92428.4]
  assign _T_931 = io_waddr == 6'h1b; // @[SRAM.scala 148:37:@92436.4]
  assign _T_932 = io_wen & _T_931; // @[SRAM.scala 148:25:@92437.4]
  assign _GEN_27 = _T_932 ? 1'h1 : regs_27; // @[SRAM.scala 148:48:@92439.4]
  assign _T_940 = io_waddr == 6'h1c; // @[SRAM.scala 148:37:@92447.4]
  assign _T_941 = io_wen & _T_940; // @[SRAM.scala 148:25:@92448.4]
  assign _GEN_28 = _T_941 ? 1'h1 : regs_28; // @[SRAM.scala 148:48:@92450.4]
  assign _T_949 = io_waddr == 6'h1d; // @[SRAM.scala 148:37:@92458.4]
  assign _T_950 = io_wen & _T_949; // @[SRAM.scala 148:25:@92459.4]
  assign _GEN_29 = _T_950 ? 1'h1 : regs_29; // @[SRAM.scala 148:48:@92461.4]
  assign _T_958 = io_waddr == 6'h1e; // @[SRAM.scala 148:37:@92469.4]
  assign _T_959 = io_wen & _T_958; // @[SRAM.scala 148:25:@92470.4]
  assign _GEN_30 = _T_959 ? 1'h1 : regs_30; // @[SRAM.scala 148:48:@92472.4]
  assign _T_967 = io_waddr == 6'h1f; // @[SRAM.scala 148:37:@92480.4]
  assign _T_968 = io_wen & _T_967; // @[SRAM.scala 148:25:@92481.4]
  assign _GEN_31 = _T_968 ? 1'h1 : regs_31; // @[SRAM.scala 148:48:@92483.4]
  assign _T_976 = io_waddr == 6'h20; // @[SRAM.scala 148:37:@92491.4]
  assign _T_977 = io_wen & _T_976; // @[SRAM.scala 148:25:@92492.4]
  assign _GEN_32 = _T_977 ? 1'h1 : regs_32; // @[SRAM.scala 148:48:@92494.4]
  assign _T_985 = io_waddr == 6'h21; // @[SRAM.scala 148:37:@92502.4]
  assign _T_986 = io_wen & _T_985; // @[SRAM.scala 148:25:@92503.4]
  assign _GEN_33 = _T_986 ? 1'h1 : regs_33; // @[SRAM.scala 148:48:@92505.4]
  assign _T_994 = io_waddr == 6'h22; // @[SRAM.scala 148:37:@92513.4]
  assign _T_995 = io_wen & _T_994; // @[SRAM.scala 148:25:@92514.4]
  assign _GEN_34 = _T_995 ? 1'h1 : regs_34; // @[SRAM.scala 148:48:@92516.4]
  assign _T_1003 = io_waddr == 6'h23; // @[SRAM.scala 148:37:@92524.4]
  assign _T_1004 = io_wen & _T_1003; // @[SRAM.scala 148:25:@92525.4]
  assign _GEN_35 = _T_1004 ? 1'h1 : regs_35; // @[SRAM.scala 148:48:@92527.4]
  assign _T_1012 = io_waddr == 6'h24; // @[SRAM.scala 148:37:@92535.4]
  assign _T_1013 = io_wen & _T_1012; // @[SRAM.scala 148:25:@92536.4]
  assign _GEN_36 = _T_1013 ? 1'h1 : regs_36; // @[SRAM.scala 148:48:@92538.4]
  assign _T_1021 = io_waddr == 6'h25; // @[SRAM.scala 148:37:@92546.4]
  assign _T_1022 = io_wen & _T_1021; // @[SRAM.scala 148:25:@92547.4]
  assign _GEN_37 = _T_1022 ? 1'h1 : regs_37; // @[SRAM.scala 148:48:@92549.4]
  assign _T_1030 = io_waddr == 6'h26; // @[SRAM.scala 148:37:@92557.4]
  assign _T_1031 = io_wen & _T_1030; // @[SRAM.scala 148:25:@92558.4]
  assign _GEN_38 = _T_1031 ? 1'h1 : regs_38; // @[SRAM.scala 148:48:@92560.4]
  assign _T_1039 = io_waddr == 6'h27; // @[SRAM.scala 148:37:@92568.4]
  assign _T_1040 = io_wen & _T_1039; // @[SRAM.scala 148:25:@92569.4]
  assign _GEN_39 = _T_1040 ? 1'h1 : regs_39; // @[SRAM.scala 148:48:@92571.4]
  assign _T_1048 = io_waddr == 6'h28; // @[SRAM.scala 148:37:@92579.4]
  assign _T_1049 = io_wen & _T_1048; // @[SRAM.scala 148:25:@92580.4]
  assign _GEN_40 = _T_1049 ? 1'h1 : regs_40; // @[SRAM.scala 148:48:@92582.4]
  assign _T_1057 = io_waddr == 6'h29; // @[SRAM.scala 148:37:@92590.4]
  assign _T_1058 = io_wen & _T_1057; // @[SRAM.scala 148:25:@92591.4]
  assign _GEN_41 = _T_1058 ? 1'h1 : regs_41; // @[SRAM.scala 148:48:@92593.4]
  assign _T_1066 = io_waddr == 6'h2a; // @[SRAM.scala 148:37:@92601.4]
  assign _T_1067 = io_wen & _T_1066; // @[SRAM.scala 148:25:@92602.4]
  assign _GEN_42 = _T_1067 ? 1'h1 : regs_42; // @[SRAM.scala 148:48:@92604.4]
  assign _T_1075 = io_waddr == 6'h2b; // @[SRAM.scala 148:37:@92612.4]
  assign _T_1076 = io_wen & _T_1075; // @[SRAM.scala 148:25:@92613.4]
  assign _GEN_43 = _T_1076 ? 1'h1 : regs_43; // @[SRAM.scala 148:48:@92615.4]
  assign _T_1084 = io_waddr == 6'h2c; // @[SRAM.scala 148:37:@92623.4]
  assign _T_1085 = io_wen & _T_1084; // @[SRAM.scala 148:25:@92624.4]
  assign _GEN_44 = _T_1085 ? 1'h1 : regs_44; // @[SRAM.scala 148:48:@92626.4]
  assign _T_1093 = io_waddr == 6'h2d; // @[SRAM.scala 148:37:@92634.4]
  assign _T_1094 = io_wen & _T_1093; // @[SRAM.scala 148:25:@92635.4]
  assign _GEN_45 = _T_1094 ? 1'h1 : regs_45; // @[SRAM.scala 148:48:@92637.4]
  assign _T_1102 = io_waddr == 6'h2e; // @[SRAM.scala 148:37:@92645.4]
  assign _T_1103 = io_wen & _T_1102; // @[SRAM.scala 148:25:@92646.4]
  assign _GEN_46 = _T_1103 ? 1'h1 : regs_46; // @[SRAM.scala 148:48:@92648.4]
  assign _T_1111 = io_waddr == 6'h2f; // @[SRAM.scala 148:37:@92656.4]
  assign _T_1112 = io_wen & _T_1111; // @[SRAM.scala 148:25:@92657.4]
  assign _GEN_47 = _T_1112 ? 1'h1 : regs_47; // @[SRAM.scala 148:48:@92659.4]
  assign _T_1120 = io_waddr == 6'h30; // @[SRAM.scala 148:37:@92667.4]
  assign _T_1121 = io_wen & _T_1120; // @[SRAM.scala 148:25:@92668.4]
  assign _GEN_48 = _T_1121 ? 1'h1 : regs_48; // @[SRAM.scala 148:48:@92670.4]
  assign _T_1129 = io_waddr == 6'h31; // @[SRAM.scala 148:37:@92678.4]
  assign _T_1130 = io_wen & _T_1129; // @[SRAM.scala 148:25:@92679.4]
  assign _GEN_49 = _T_1130 ? 1'h1 : regs_49; // @[SRAM.scala 148:48:@92681.4]
  assign _T_1138 = io_waddr == 6'h32; // @[SRAM.scala 148:37:@92689.4]
  assign _T_1139 = io_wen & _T_1138; // @[SRAM.scala 148:25:@92690.4]
  assign _GEN_50 = _T_1139 ? 1'h1 : regs_50; // @[SRAM.scala 148:48:@92692.4]
  assign _T_1147 = io_waddr == 6'h33; // @[SRAM.scala 148:37:@92700.4]
  assign _T_1148 = io_wen & _T_1147; // @[SRAM.scala 148:25:@92701.4]
  assign _GEN_51 = _T_1148 ? 1'h1 : regs_51; // @[SRAM.scala 148:48:@92703.4]
  assign _T_1156 = io_waddr == 6'h34; // @[SRAM.scala 148:37:@92711.4]
  assign _T_1157 = io_wen & _T_1156; // @[SRAM.scala 148:25:@92712.4]
  assign _GEN_52 = _T_1157 ? 1'h1 : regs_52; // @[SRAM.scala 148:48:@92714.4]
  assign _T_1165 = io_waddr == 6'h35; // @[SRAM.scala 148:37:@92722.4]
  assign _T_1166 = io_wen & _T_1165; // @[SRAM.scala 148:25:@92723.4]
  assign _GEN_53 = _T_1166 ? 1'h1 : regs_53; // @[SRAM.scala 148:48:@92725.4]
  assign _T_1174 = io_waddr == 6'h36; // @[SRAM.scala 148:37:@92733.4]
  assign _T_1175 = io_wen & _T_1174; // @[SRAM.scala 148:25:@92734.4]
  assign _GEN_54 = _T_1175 ? 1'h1 : regs_54; // @[SRAM.scala 148:48:@92736.4]
  assign _T_1183 = io_waddr == 6'h37; // @[SRAM.scala 148:37:@92744.4]
  assign _T_1184 = io_wen & _T_1183; // @[SRAM.scala 148:25:@92745.4]
  assign _GEN_55 = _T_1184 ? 1'h1 : regs_55; // @[SRAM.scala 148:48:@92747.4]
  assign _T_1192 = io_waddr == 6'h38; // @[SRAM.scala 148:37:@92755.4]
  assign _T_1193 = io_wen & _T_1192; // @[SRAM.scala 148:25:@92756.4]
  assign _GEN_56 = _T_1193 ? 1'h1 : regs_56; // @[SRAM.scala 148:48:@92758.4]
  assign _T_1201 = io_waddr == 6'h39; // @[SRAM.scala 148:37:@92766.4]
  assign _T_1202 = io_wen & _T_1201; // @[SRAM.scala 148:25:@92767.4]
  assign _GEN_57 = _T_1202 ? 1'h1 : regs_57; // @[SRAM.scala 148:48:@92769.4]
  assign _T_1210 = io_waddr == 6'h3a; // @[SRAM.scala 148:37:@92777.4]
  assign _T_1211 = io_wen & _T_1210; // @[SRAM.scala 148:25:@92778.4]
  assign _GEN_58 = _T_1211 ? 1'h1 : regs_58; // @[SRAM.scala 148:48:@92780.4]
  assign _T_1219 = io_waddr == 6'h3b; // @[SRAM.scala 148:37:@92788.4]
  assign _T_1220 = io_wen & _T_1219; // @[SRAM.scala 148:25:@92789.4]
  assign _GEN_59 = _T_1220 ? 1'h1 : regs_59; // @[SRAM.scala 148:48:@92791.4]
  assign _T_1228 = io_waddr == 6'h3c; // @[SRAM.scala 148:37:@92799.4]
  assign _T_1229 = io_wen & _T_1228; // @[SRAM.scala 148:25:@92800.4]
  assign _GEN_60 = _T_1229 ? 1'h1 : regs_60; // @[SRAM.scala 148:48:@92802.4]
  assign _T_1237 = io_waddr == 6'h3d; // @[SRAM.scala 148:37:@92810.4]
  assign _T_1238 = io_wen & _T_1237; // @[SRAM.scala 148:25:@92811.4]
  assign _GEN_61 = _T_1238 ? 1'h1 : regs_61; // @[SRAM.scala 148:48:@92813.4]
  assign _T_1246 = io_waddr == 6'h3e; // @[SRAM.scala 148:37:@92821.4]
  assign _T_1247 = io_wen & _T_1246; // @[SRAM.scala 148:25:@92822.4]
  assign _GEN_62 = _T_1247 ? 1'h1 : regs_62; // @[SRAM.scala 148:48:@92824.4]
  assign _T_1255 = io_waddr == 6'h3f; // @[SRAM.scala 148:37:@92832.4]
  assign _T_1256 = io_wen & _T_1255; // @[SRAM.scala 148:25:@92833.4]
  assign _GEN_63 = _T_1256 ? 1'h1 : regs_63; // @[SRAM.scala 148:48:@92835.4]
  assign _GEN_65 = 6'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_66 = 6'h2 == io_raddr ? regs_2 : _GEN_65; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_67 = 6'h3 == io_raddr ? regs_3 : _GEN_66; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_68 = 6'h4 == io_raddr ? regs_4 : _GEN_67; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_69 = 6'h5 == io_raddr ? regs_5 : _GEN_68; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_70 = 6'h6 == io_raddr ? regs_6 : _GEN_69; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_71 = 6'h7 == io_raddr ? regs_7 : _GEN_70; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_72 = 6'h8 == io_raddr ? regs_8 : _GEN_71; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_73 = 6'h9 == io_raddr ? regs_9 : _GEN_72; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_74 = 6'ha == io_raddr ? regs_10 : _GEN_73; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_75 = 6'hb == io_raddr ? regs_11 : _GEN_74; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_76 = 6'hc == io_raddr ? regs_12 : _GEN_75; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_77 = 6'hd == io_raddr ? regs_13 : _GEN_76; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_78 = 6'he == io_raddr ? regs_14 : _GEN_77; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_79 = 6'hf == io_raddr ? regs_15 : _GEN_78; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_80 = 6'h10 == io_raddr ? regs_16 : _GEN_79; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_81 = 6'h11 == io_raddr ? regs_17 : _GEN_80; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_82 = 6'h12 == io_raddr ? regs_18 : _GEN_81; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_83 = 6'h13 == io_raddr ? regs_19 : _GEN_82; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_84 = 6'h14 == io_raddr ? regs_20 : _GEN_83; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_85 = 6'h15 == io_raddr ? regs_21 : _GEN_84; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_86 = 6'h16 == io_raddr ? regs_22 : _GEN_85; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_87 = 6'h17 == io_raddr ? regs_23 : _GEN_86; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_88 = 6'h18 == io_raddr ? regs_24 : _GEN_87; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_89 = 6'h19 == io_raddr ? regs_25 : _GEN_88; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_90 = 6'h1a == io_raddr ? regs_26 : _GEN_89; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_91 = 6'h1b == io_raddr ? regs_27 : _GEN_90; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_92 = 6'h1c == io_raddr ? regs_28 : _GEN_91; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_93 = 6'h1d == io_raddr ? regs_29 : _GEN_92; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_94 = 6'h1e == io_raddr ? regs_30 : _GEN_93; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_95 = 6'h1f == io_raddr ? regs_31 : _GEN_94; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_96 = 6'h20 == io_raddr ? regs_32 : _GEN_95; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_97 = 6'h21 == io_raddr ? regs_33 : _GEN_96; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_98 = 6'h22 == io_raddr ? regs_34 : _GEN_97; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_99 = 6'h23 == io_raddr ? regs_35 : _GEN_98; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_100 = 6'h24 == io_raddr ? regs_36 : _GEN_99; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_101 = 6'h25 == io_raddr ? regs_37 : _GEN_100; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_102 = 6'h26 == io_raddr ? regs_38 : _GEN_101; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_103 = 6'h27 == io_raddr ? regs_39 : _GEN_102; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_104 = 6'h28 == io_raddr ? regs_40 : _GEN_103; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_105 = 6'h29 == io_raddr ? regs_41 : _GEN_104; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_106 = 6'h2a == io_raddr ? regs_42 : _GEN_105; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_107 = 6'h2b == io_raddr ? regs_43 : _GEN_106; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_108 = 6'h2c == io_raddr ? regs_44 : _GEN_107; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_109 = 6'h2d == io_raddr ? regs_45 : _GEN_108; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_110 = 6'h2e == io_raddr ? regs_46 : _GEN_109; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_111 = 6'h2f == io_raddr ? regs_47 : _GEN_110; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_112 = 6'h30 == io_raddr ? regs_48 : _GEN_111; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_113 = 6'h31 == io_raddr ? regs_49 : _GEN_112; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_114 = 6'h32 == io_raddr ? regs_50 : _GEN_113; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_115 = 6'h33 == io_raddr ? regs_51 : _GEN_114; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_116 = 6'h34 == io_raddr ? regs_52 : _GEN_115; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_117 = 6'h35 == io_raddr ? regs_53 : _GEN_116; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_118 = 6'h36 == io_raddr ? regs_54 : _GEN_117; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_119 = 6'h37 == io_raddr ? regs_55 : _GEN_118; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_120 = 6'h38 == io_raddr ? regs_56 : _GEN_119; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_121 = 6'h39 == io_raddr ? regs_57 : _GEN_120; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_122 = 6'h3a == io_raddr ? regs_58 : _GEN_121; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_123 = 6'h3b == io_raddr ? regs_59 : _GEN_122; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_124 = 6'h3c == io_raddr ? regs_60 : _GEN_123; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_125 = 6'h3d == io_raddr ? regs_61 : _GEN_124; // @[SRAM.scala 155:12:@92905.4]
  assign _GEN_126 = 6'h3e == io_raddr ? regs_62 : _GEN_125; // @[SRAM.scala 155:12:@92905.4]
  assign io_rdata = 6'h3f == io_raddr ? regs_63 : _GEN_126; // @[SRAM.scala 155:12:@92905.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_689) begin
        regs_0 <= 1'h1;
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_698) begin
        regs_1 <= 1'h1;
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_707) begin
        regs_2 <= 1'h1;
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_716) begin
        regs_3 <= 1'h1;
      end
    end
    if (reset) begin
      regs_4 <= 1'h0;
    end else begin
      if (_T_725) begin
        regs_4 <= 1'h1;
      end
    end
    if (reset) begin
      regs_5 <= 1'h0;
    end else begin
      if (_T_734) begin
        regs_5 <= 1'h1;
      end
    end
    if (reset) begin
      regs_6 <= 1'h0;
    end else begin
      if (_T_743) begin
        regs_6 <= 1'h1;
      end
    end
    if (reset) begin
      regs_7 <= 1'h0;
    end else begin
      if (_T_752) begin
        regs_7 <= 1'h1;
      end
    end
    if (reset) begin
      regs_8 <= 1'h0;
    end else begin
      if (_T_761) begin
        regs_8 <= 1'h1;
      end
    end
    if (reset) begin
      regs_9 <= 1'h0;
    end else begin
      if (_T_770) begin
        regs_9 <= 1'h1;
      end
    end
    if (reset) begin
      regs_10 <= 1'h0;
    end else begin
      if (_T_779) begin
        regs_10 <= 1'h1;
      end
    end
    if (reset) begin
      regs_11 <= 1'h0;
    end else begin
      if (_T_788) begin
        regs_11 <= 1'h1;
      end
    end
    if (reset) begin
      regs_12 <= 1'h0;
    end else begin
      if (_T_797) begin
        regs_12 <= 1'h1;
      end
    end
    if (reset) begin
      regs_13 <= 1'h0;
    end else begin
      if (_T_806) begin
        regs_13 <= 1'h1;
      end
    end
    if (reset) begin
      regs_14 <= 1'h0;
    end else begin
      if (_T_815) begin
        regs_14 <= 1'h1;
      end
    end
    if (reset) begin
      regs_15 <= 1'h0;
    end else begin
      if (_T_824) begin
        regs_15 <= 1'h1;
      end
    end
    if (reset) begin
      regs_16 <= 1'h0;
    end else begin
      if (_T_833) begin
        regs_16 <= 1'h1;
      end
    end
    if (reset) begin
      regs_17 <= 1'h0;
    end else begin
      if (_T_842) begin
        regs_17 <= 1'h1;
      end
    end
    if (reset) begin
      regs_18 <= 1'h0;
    end else begin
      if (_T_851) begin
        regs_18 <= 1'h1;
      end
    end
    if (reset) begin
      regs_19 <= 1'h0;
    end else begin
      if (_T_860) begin
        regs_19 <= 1'h1;
      end
    end
    if (reset) begin
      regs_20 <= 1'h0;
    end else begin
      if (_T_869) begin
        regs_20 <= 1'h1;
      end
    end
    if (reset) begin
      regs_21 <= 1'h0;
    end else begin
      if (_T_878) begin
        regs_21 <= 1'h1;
      end
    end
    if (reset) begin
      regs_22 <= 1'h0;
    end else begin
      if (_T_887) begin
        regs_22 <= 1'h1;
      end
    end
    if (reset) begin
      regs_23 <= 1'h0;
    end else begin
      if (_T_896) begin
        regs_23 <= 1'h1;
      end
    end
    if (reset) begin
      regs_24 <= 1'h0;
    end else begin
      if (_T_905) begin
        regs_24 <= 1'h1;
      end
    end
    if (reset) begin
      regs_25 <= 1'h0;
    end else begin
      if (_T_914) begin
        regs_25 <= 1'h1;
      end
    end
    if (reset) begin
      regs_26 <= 1'h0;
    end else begin
      if (_T_923) begin
        regs_26 <= 1'h1;
      end
    end
    if (reset) begin
      regs_27 <= 1'h0;
    end else begin
      if (_T_932) begin
        regs_27 <= 1'h1;
      end
    end
    if (reset) begin
      regs_28 <= 1'h0;
    end else begin
      if (_T_941) begin
        regs_28 <= 1'h1;
      end
    end
    if (reset) begin
      regs_29 <= 1'h0;
    end else begin
      if (_T_950) begin
        regs_29 <= 1'h1;
      end
    end
    if (reset) begin
      regs_30 <= 1'h0;
    end else begin
      if (_T_959) begin
        regs_30 <= 1'h1;
      end
    end
    if (reset) begin
      regs_31 <= 1'h0;
    end else begin
      if (_T_968) begin
        regs_31 <= 1'h1;
      end
    end
    if (reset) begin
      regs_32 <= 1'h0;
    end else begin
      if (_T_977) begin
        regs_32 <= 1'h1;
      end
    end
    if (reset) begin
      regs_33 <= 1'h0;
    end else begin
      if (_T_986) begin
        regs_33 <= 1'h1;
      end
    end
    if (reset) begin
      regs_34 <= 1'h0;
    end else begin
      if (_T_995) begin
        regs_34 <= 1'h1;
      end
    end
    if (reset) begin
      regs_35 <= 1'h0;
    end else begin
      if (_T_1004) begin
        regs_35 <= 1'h1;
      end
    end
    if (reset) begin
      regs_36 <= 1'h0;
    end else begin
      if (_T_1013) begin
        regs_36 <= 1'h1;
      end
    end
    if (reset) begin
      regs_37 <= 1'h0;
    end else begin
      if (_T_1022) begin
        regs_37 <= 1'h1;
      end
    end
    if (reset) begin
      regs_38 <= 1'h0;
    end else begin
      if (_T_1031) begin
        regs_38 <= 1'h1;
      end
    end
    if (reset) begin
      regs_39 <= 1'h0;
    end else begin
      if (_T_1040) begin
        regs_39 <= 1'h1;
      end
    end
    if (reset) begin
      regs_40 <= 1'h0;
    end else begin
      if (_T_1049) begin
        regs_40 <= 1'h1;
      end
    end
    if (reset) begin
      regs_41 <= 1'h0;
    end else begin
      if (_T_1058) begin
        regs_41 <= 1'h1;
      end
    end
    if (reset) begin
      regs_42 <= 1'h0;
    end else begin
      if (_T_1067) begin
        regs_42 <= 1'h1;
      end
    end
    if (reset) begin
      regs_43 <= 1'h0;
    end else begin
      if (_T_1076) begin
        regs_43 <= 1'h1;
      end
    end
    if (reset) begin
      regs_44 <= 1'h0;
    end else begin
      if (_T_1085) begin
        regs_44 <= 1'h1;
      end
    end
    if (reset) begin
      regs_45 <= 1'h0;
    end else begin
      if (_T_1094) begin
        regs_45 <= 1'h1;
      end
    end
    if (reset) begin
      regs_46 <= 1'h0;
    end else begin
      if (_T_1103) begin
        regs_46 <= 1'h1;
      end
    end
    if (reset) begin
      regs_47 <= 1'h0;
    end else begin
      if (_T_1112) begin
        regs_47 <= 1'h1;
      end
    end
    if (reset) begin
      regs_48 <= 1'h0;
    end else begin
      if (_T_1121) begin
        regs_48 <= 1'h1;
      end
    end
    if (reset) begin
      regs_49 <= 1'h0;
    end else begin
      if (_T_1130) begin
        regs_49 <= 1'h1;
      end
    end
    if (reset) begin
      regs_50 <= 1'h0;
    end else begin
      if (_T_1139) begin
        regs_50 <= 1'h1;
      end
    end
    if (reset) begin
      regs_51 <= 1'h0;
    end else begin
      if (_T_1148) begin
        regs_51 <= 1'h1;
      end
    end
    if (reset) begin
      regs_52 <= 1'h0;
    end else begin
      if (_T_1157) begin
        regs_52 <= 1'h1;
      end
    end
    if (reset) begin
      regs_53 <= 1'h0;
    end else begin
      if (_T_1166) begin
        regs_53 <= 1'h1;
      end
    end
    if (reset) begin
      regs_54 <= 1'h0;
    end else begin
      if (_T_1175) begin
        regs_54 <= 1'h1;
      end
    end
    if (reset) begin
      regs_55 <= 1'h0;
    end else begin
      if (_T_1184) begin
        regs_55 <= 1'h1;
      end
    end
    if (reset) begin
      regs_56 <= 1'h0;
    end else begin
      if (_T_1193) begin
        regs_56 <= 1'h1;
      end
    end
    if (reset) begin
      regs_57 <= 1'h0;
    end else begin
      if (_T_1202) begin
        regs_57 <= 1'h1;
      end
    end
    if (reset) begin
      regs_58 <= 1'h0;
    end else begin
      if (_T_1211) begin
        regs_58 <= 1'h1;
      end
    end
    if (reset) begin
      regs_59 <= 1'h0;
    end else begin
      if (_T_1220) begin
        regs_59 <= 1'h1;
      end
    end
    if (reset) begin
      regs_60 <= 1'h0;
    end else begin
      if (_T_1229) begin
        regs_60 <= 1'h1;
      end
    end
    if (reset) begin
      regs_61 <= 1'h0;
    end else begin
      if (_T_1238) begin
        regs_61 <= 1'h1;
      end
    end
    if (reset) begin
      regs_62 <= 1'h0;
    end else begin
      if (_T_1247) begin
        regs_62 <= 1'h1;
      end
    end
    if (reset) begin
      regs_63 <= 1'h0;
    end else begin
      if (_T_1256) begin
        regs_63 <= 1'h1;
      end
    end
  end
endmodule
module FIFO_51( // @[:@92907.2]
  input   clock, // @[:@92908.4]
  input   reset, // @[:@92909.4]
  output  io_in_ready, // @[:@92910.4]
  input   io_in_valid, // @[:@92910.4]
  input   io_out_ready, // @[:@92910.4]
  output  io_out_valid, // @[:@92910.4]
  output  io_out_bits // @[:@92910.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@93176.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@93176.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@93176.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@93176.4]
  wire [5:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@93176.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@93176.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@93176.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@93186.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@93186.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@93186.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@93186.4]
  wire [5:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@93186.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@93186.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@93186.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@93201.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@93201.4]
  wire [5:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@93201.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@93201.4]
  wire [5:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@93201.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@93201.4]
  wire  writeEn; // @[FIFO.scala 30:29:@93174.4]
  wire  readEn; // @[FIFO.scala 31:29:@93175.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@93196.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@93197.4]
  wire  _T_824; // @[FIFO.scala 45:27:@93198.4]
  wire  empty; // @[FIFO.scala 45:24:@93199.4]
  wire  full; // @[FIFO.scala 46:23:@93200.4]
  wire  _T_1657; // @[FIFO.scala 83:17:@94367.4]
  wire  _GEN_64; // @[FIFO.scala 83:29:@94368.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@93176.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@93186.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM_16 FFRAM ( // @[FIFO.scala 49:19:@93201.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_rdata(FFRAM_io_rdata)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@93174.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@93175.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@93197.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@93198.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@93199.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@93200.4]
  assign _T_1657 = writeEn != readEn; // @[FIFO.scala 83:17:@94367.4]
  assign _GEN_64 = _T_1657 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@94368.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@94374.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@94372.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@93406.4]
  assign enqCounter_clock = clock; // @[:@93177.4]
  assign enqCounter_reset = reset; // @[:@93178.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@93184.4]
  assign enqCounter_io_stride = 6'h1; // @[FIFO.scala 37:24:@93185.4]
  assign deqCounter_clock = clock; // @[:@93187.4]
  assign deqCounter_reset = reset; // @[:@93188.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@93194.4]
  assign deqCounter_io_stride = 6'h1; // @[FIFO.scala 41:24:@93195.4]
  assign FFRAM_clock = clock; // @[:@93202.4]
  assign FFRAM_reset = reset; // @[:@93203.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@93402.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@93403.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@93404.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_1657) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module StreamControllerStore( // @[:@94376.2]
  input         clock, // @[:@94377.4]
  input         reset, // @[:@94378.4]
  input         io_dram_cmd_ready, // @[:@94379.4]
  output        io_dram_cmd_valid, // @[:@94379.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@94379.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@94379.4]
  input         io_dram_wdata_ready, // @[:@94379.4]
  output        io_dram_wdata_valid, // @[:@94379.4]
  output [63:0] io_dram_wdata_bits_wdata_0, // @[:@94379.4]
  output [63:0] io_dram_wdata_bits_wdata_1, // @[:@94379.4]
  output [63:0] io_dram_wdata_bits_wdata_2, // @[:@94379.4]
  output [63:0] io_dram_wdata_bits_wdata_3, // @[:@94379.4]
  output [63:0] io_dram_wdata_bits_wdata_4, // @[:@94379.4]
  output [63:0] io_dram_wdata_bits_wdata_5, // @[:@94379.4]
  output [63:0] io_dram_wdata_bits_wdata_6, // @[:@94379.4]
  output [63:0] io_dram_wdata_bits_wdata_7, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@94379.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@94379.4]
  output        io_dram_wresp_ready, // @[:@94379.4]
  input         io_dram_wresp_valid, // @[:@94379.4]
  output        io_store_cmd_ready, // @[:@94379.4]
  input         io_store_cmd_valid, // @[:@94379.4]
  input  [63:0] io_store_cmd_bits_addr, // @[:@94379.4]
  input  [31:0] io_store_cmd_bits_size, // @[:@94379.4]
  output        io_store_data_ready, // @[:@94379.4]
  input         io_store_data_valid, // @[:@94379.4]
  input  [31:0] io_store_data_bits_wdata_0, // @[:@94379.4]
  input         io_store_data_bits_wstrb, // @[:@94379.4]
  input         io_store_wresp_ready, // @[:@94379.4]
  output        io_store_wresp_valid, // @[:@94379.4]
  output        io_store_wresp_bits // @[:@94379.4]
);
  wire  cmd_clock; // @[StreamController.scala 75:19:@94488.4]
  wire  cmd_reset; // @[StreamController.scala 75:19:@94488.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 75:19:@94488.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 75:19:@94488.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 75:19:@94488.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 75:19:@94488.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 75:19:@94488.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 75:19:@94488.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 75:19:@94488.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 75:19:@94488.4]
  wire  wdata_clock; // @[StreamController.scala 88:21:@94894.4]
  wire  wdata_reset; // @[StreamController.scala 88:21:@94894.4]
  wire  wdata_io_in_ready; // @[StreamController.scala 88:21:@94894.4]
  wire  wdata_io_in_valid; // @[StreamController.scala 88:21:@94894.4]
  wire [31:0] wdata_io_in_bits_data_0; // @[StreamController.scala 88:21:@94894.4]
  wire  wdata_io_in_bits_strobe; // @[StreamController.scala 88:21:@94894.4]
  wire  wdata_io_out_ready; // @[StreamController.scala 88:21:@94894.4]
  wire  wdata_io_out_valid; // @[StreamController.scala 88:21:@94894.4]
  wire [63:0] wdata_io_out_bits_data_0; // @[StreamController.scala 88:21:@94894.4]
  wire [63:0] wdata_io_out_bits_data_1; // @[StreamController.scala 88:21:@94894.4]
  wire [63:0] wdata_io_out_bits_data_2; // @[StreamController.scala 88:21:@94894.4]
  wire [63:0] wdata_io_out_bits_data_3; // @[StreamController.scala 88:21:@94894.4]
  wire [63:0] wdata_io_out_bits_data_4; // @[StreamController.scala 88:21:@94894.4]
  wire [63:0] wdata_io_out_bits_data_5; // @[StreamController.scala 88:21:@94894.4]
  wire [63:0] wdata_io_out_bits_data_6; // @[StreamController.scala 88:21:@94894.4]
  wire [63:0] wdata_io_out_bits_data_7; // @[StreamController.scala 88:21:@94894.4]
  wire [63:0] wdata_io_out_bits_strobe; // @[StreamController.scala 88:21:@94894.4]
  wire  wresp_clock; // @[StreamController.scala 100:21:@95119.4]
  wire  wresp_reset; // @[StreamController.scala 100:21:@95119.4]
  wire  wresp_io_in_ready; // @[StreamController.scala 100:21:@95119.4]
  wire  wresp_io_in_valid; // @[StreamController.scala 100:21:@95119.4]
  wire  wresp_io_out_ready; // @[StreamController.scala 100:21:@95119.4]
  wire  wresp_io_out_valid; // @[StreamController.scala 100:21:@95119.4]
  wire  wresp_io_out_bits; // @[StreamController.scala 100:21:@95119.4]
  wire [25:0] _T_111; // @[StreamController.scala 21:10:@94891.4]
  FIFO cmd ( // @[StreamController.scala 75:19:@94488.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert_1 wdata ( // @[StreamController.scala 88:21:@94894.4]
    .clock(wdata_clock),
    .reset(wdata_reset),
    .io_in_ready(wdata_io_in_ready),
    .io_in_valid(wdata_io_in_valid),
    .io_in_bits_data_0(wdata_io_in_bits_data_0),
    .io_in_bits_strobe(wdata_io_in_bits_strobe),
    .io_out_ready(wdata_io_out_ready),
    .io_out_valid(wdata_io_out_valid),
    .io_out_bits_data_0(wdata_io_out_bits_data_0),
    .io_out_bits_data_1(wdata_io_out_bits_data_1),
    .io_out_bits_data_2(wdata_io_out_bits_data_2),
    .io_out_bits_data_3(wdata_io_out_bits_data_3),
    .io_out_bits_data_4(wdata_io_out_bits_data_4),
    .io_out_bits_data_5(wdata_io_out_bits_data_5),
    .io_out_bits_data_6(wdata_io_out_bits_data_6),
    .io_out_bits_data_7(wdata_io_out_bits_data_7),
    .io_out_bits_strobe(wdata_io_out_bits_strobe)
  );
  FIFO_51 wresp ( // @[StreamController.scala 100:21:@95119.4]
    .clock(wresp_clock),
    .reset(wresp_reset),
    .io_in_ready(wresp_io_in_ready),
    .io_in_valid(wresp_io_in_valid),
    .io_out_ready(wresp_io_out_ready),
    .io_out_valid(wresp_io_out_valid),
    .io_out_bits(wresp_io_out_bits)
  );
  assign _T_111 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@94891.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 81:21:@94888.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 83:25:@94889.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_111}; // @[StreamController.scala 85:25:@94892.4]
  assign io_dram_wdata_valid = wdata_io_out_valid; // @[StreamController.scala 95:23:@94916.4]
  assign io_dram_wdata_bits_wdata_0 = wdata_io_out_bits_data_0; // @[StreamController.scala 96:28:@94917.4]
  assign io_dram_wdata_bits_wdata_1 = wdata_io_out_bits_data_1; // @[StreamController.scala 96:28:@94918.4]
  assign io_dram_wdata_bits_wdata_2 = wdata_io_out_bits_data_2; // @[StreamController.scala 96:28:@94919.4]
  assign io_dram_wdata_bits_wdata_3 = wdata_io_out_bits_data_3; // @[StreamController.scala 96:28:@94920.4]
  assign io_dram_wdata_bits_wdata_4 = wdata_io_out_bits_data_4; // @[StreamController.scala 96:28:@94921.4]
  assign io_dram_wdata_bits_wdata_5 = wdata_io_out_bits_data_5; // @[StreamController.scala 96:28:@94922.4]
  assign io_dram_wdata_bits_wdata_6 = wdata_io_out_bits_data_6; // @[StreamController.scala 96:28:@94923.4]
  assign io_dram_wdata_bits_wdata_7 = wdata_io_out_bits_data_7; // @[StreamController.scala 96:28:@94924.4]
  assign io_dram_wdata_bits_wstrb_0 = wdata_io_out_bits_strobe[63]; // @[StreamController.scala 97:28:@95054.4]
  assign io_dram_wdata_bits_wstrb_1 = wdata_io_out_bits_strobe[62]; // @[StreamController.scala 97:28:@95055.4]
  assign io_dram_wdata_bits_wstrb_2 = wdata_io_out_bits_strobe[61]; // @[StreamController.scala 97:28:@95056.4]
  assign io_dram_wdata_bits_wstrb_3 = wdata_io_out_bits_strobe[60]; // @[StreamController.scala 97:28:@95057.4]
  assign io_dram_wdata_bits_wstrb_4 = wdata_io_out_bits_strobe[59]; // @[StreamController.scala 97:28:@95058.4]
  assign io_dram_wdata_bits_wstrb_5 = wdata_io_out_bits_strobe[58]; // @[StreamController.scala 97:28:@95059.4]
  assign io_dram_wdata_bits_wstrb_6 = wdata_io_out_bits_strobe[57]; // @[StreamController.scala 97:28:@95060.4]
  assign io_dram_wdata_bits_wstrb_7 = wdata_io_out_bits_strobe[56]; // @[StreamController.scala 97:28:@95061.4]
  assign io_dram_wdata_bits_wstrb_8 = wdata_io_out_bits_strobe[55]; // @[StreamController.scala 97:28:@95062.4]
  assign io_dram_wdata_bits_wstrb_9 = wdata_io_out_bits_strobe[54]; // @[StreamController.scala 97:28:@95063.4]
  assign io_dram_wdata_bits_wstrb_10 = wdata_io_out_bits_strobe[53]; // @[StreamController.scala 97:28:@95064.4]
  assign io_dram_wdata_bits_wstrb_11 = wdata_io_out_bits_strobe[52]; // @[StreamController.scala 97:28:@95065.4]
  assign io_dram_wdata_bits_wstrb_12 = wdata_io_out_bits_strobe[51]; // @[StreamController.scala 97:28:@95066.4]
  assign io_dram_wdata_bits_wstrb_13 = wdata_io_out_bits_strobe[50]; // @[StreamController.scala 97:28:@95067.4]
  assign io_dram_wdata_bits_wstrb_14 = wdata_io_out_bits_strobe[49]; // @[StreamController.scala 97:28:@95068.4]
  assign io_dram_wdata_bits_wstrb_15 = wdata_io_out_bits_strobe[48]; // @[StreamController.scala 97:28:@95069.4]
  assign io_dram_wdata_bits_wstrb_16 = wdata_io_out_bits_strobe[47]; // @[StreamController.scala 97:28:@95070.4]
  assign io_dram_wdata_bits_wstrb_17 = wdata_io_out_bits_strobe[46]; // @[StreamController.scala 97:28:@95071.4]
  assign io_dram_wdata_bits_wstrb_18 = wdata_io_out_bits_strobe[45]; // @[StreamController.scala 97:28:@95072.4]
  assign io_dram_wdata_bits_wstrb_19 = wdata_io_out_bits_strobe[44]; // @[StreamController.scala 97:28:@95073.4]
  assign io_dram_wdata_bits_wstrb_20 = wdata_io_out_bits_strobe[43]; // @[StreamController.scala 97:28:@95074.4]
  assign io_dram_wdata_bits_wstrb_21 = wdata_io_out_bits_strobe[42]; // @[StreamController.scala 97:28:@95075.4]
  assign io_dram_wdata_bits_wstrb_22 = wdata_io_out_bits_strobe[41]; // @[StreamController.scala 97:28:@95076.4]
  assign io_dram_wdata_bits_wstrb_23 = wdata_io_out_bits_strobe[40]; // @[StreamController.scala 97:28:@95077.4]
  assign io_dram_wdata_bits_wstrb_24 = wdata_io_out_bits_strobe[39]; // @[StreamController.scala 97:28:@95078.4]
  assign io_dram_wdata_bits_wstrb_25 = wdata_io_out_bits_strobe[38]; // @[StreamController.scala 97:28:@95079.4]
  assign io_dram_wdata_bits_wstrb_26 = wdata_io_out_bits_strobe[37]; // @[StreamController.scala 97:28:@95080.4]
  assign io_dram_wdata_bits_wstrb_27 = wdata_io_out_bits_strobe[36]; // @[StreamController.scala 97:28:@95081.4]
  assign io_dram_wdata_bits_wstrb_28 = wdata_io_out_bits_strobe[35]; // @[StreamController.scala 97:28:@95082.4]
  assign io_dram_wdata_bits_wstrb_29 = wdata_io_out_bits_strobe[34]; // @[StreamController.scala 97:28:@95083.4]
  assign io_dram_wdata_bits_wstrb_30 = wdata_io_out_bits_strobe[33]; // @[StreamController.scala 97:28:@95084.4]
  assign io_dram_wdata_bits_wstrb_31 = wdata_io_out_bits_strobe[32]; // @[StreamController.scala 97:28:@95085.4]
  assign io_dram_wdata_bits_wstrb_32 = wdata_io_out_bits_strobe[31]; // @[StreamController.scala 97:28:@95086.4]
  assign io_dram_wdata_bits_wstrb_33 = wdata_io_out_bits_strobe[30]; // @[StreamController.scala 97:28:@95087.4]
  assign io_dram_wdata_bits_wstrb_34 = wdata_io_out_bits_strobe[29]; // @[StreamController.scala 97:28:@95088.4]
  assign io_dram_wdata_bits_wstrb_35 = wdata_io_out_bits_strobe[28]; // @[StreamController.scala 97:28:@95089.4]
  assign io_dram_wdata_bits_wstrb_36 = wdata_io_out_bits_strobe[27]; // @[StreamController.scala 97:28:@95090.4]
  assign io_dram_wdata_bits_wstrb_37 = wdata_io_out_bits_strobe[26]; // @[StreamController.scala 97:28:@95091.4]
  assign io_dram_wdata_bits_wstrb_38 = wdata_io_out_bits_strobe[25]; // @[StreamController.scala 97:28:@95092.4]
  assign io_dram_wdata_bits_wstrb_39 = wdata_io_out_bits_strobe[24]; // @[StreamController.scala 97:28:@95093.4]
  assign io_dram_wdata_bits_wstrb_40 = wdata_io_out_bits_strobe[23]; // @[StreamController.scala 97:28:@95094.4]
  assign io_dram_wdata_bits_wstrb_41 = wdata_io_out_bits_strobe[22]; // @[StreamController.scala 97:28:@95095.4]
  assign io_dram_wdata_bits_wstrb_42 = wdata_io_out_bits_strobe[21]; // @[StreamController.scala 97:28:@95096.4]
  assign io_dram_wdata_bits_wstrb_43 = wdata_io_out_bits_strobe[20]; // @[StreamController.scala 97:28:@95097.4]
  assign io_dram_wdata_bits_wstrb_44 = wdata_io_out_bits_strobe[19]; // @[StreamController.scala 97:28:@95098.4]
  assign io_dram_wdata_bits_wstrb_45 = wdata_io_out_bits_strobe[18]; // @[StreamController.scala 97:28:@95099.4]
  assign io_dram_wdata_bits_wstrb_46 = wdata_io_out_bits_strobe[17]; // @[StreamController.scala 97:28:@95100.4]
  assign io_dram_wdata_bits_wstrb_47 = wdata_io_out_bits_strobe[16]; // @[StreamController.scala 97:28:@95101.4]
  assign io_dram_wdata_bits_wstrb_48 = wdata_io_out_bits_strobe[15]; // @[StreamController.scala 97:28:@95102.4]
  assign io_dram_wdata_bits_wstrb_49 = wdata_io_out_bits_strobe[14]; // @[StreamController.scala 97:28:@95103.4]
  assign io_dram_wdata_bits_wstrb_50 = wdata_io_out_bits_strobe[13]; // @[StreamController.scala 97:28:@95104.4]
  assign io_dram_wdata_bits_wstrb_51 = wdata_io_out_bits_strobe[12]; // @[StreamController.scala 97:28:@95105.4]
  assign io_dram_wdata_bits_wstrb_52 = wdata_io_out_bits_strobe[11]; // @[StreamController.scala 97:28:@95106.4]
  assign io_dram_wdata_bits_wstrb_53 = wdata_io_out_bits_strobe[10]; // @[StreamController.scala 97:28:@95107.4]
  assign io_dram_wdata_bits_wstrb_54 = wdata_io_out_bits_strobe[9]; // @[StreamController.scala 97:28:@95108.4]
  assign io_dram_wdata_bits_wstrb_55 = wdata_io_out_bits_strobe[8]; // @[StreamController.scala 97:28:@95109.4]
  assign io_dram_wdata_bits_wstrb_56 = wdata_io_out_bits_strobe[7]; // @[StreamController.scala 97:28:@95110.4]
  assign io_dram_wdata_bits_wstrb_57 = wdata_io_out_bits_strobe[6]; // @[StreamController.scala 97:28:@95111.4]
  assign io_dram_wdata_bits_wstrb_58 = wdata_io_out_bits_strobe[5]; // @[StreamController.scala 97:28:@95112.4]
  assign io_dram_wdata_bits_wstrb_59 = wdata_io_out_bits_strobe[4]; // @[StreamController.scala 97:28:@95113.4]
  assign io_dram_wdata_bits_wstrb_60 = wdata_io_out_bits_strobe[3]; // @[StreamController.scala 97:28:@95114.4]
  assign io_dram_wdata_bits_wstrb_61 = wdata_io_out_bits_strobe[2]; // @[StreamController.scala 97:28:@95115.4]
  assign io_dram_wdata_bits_wstrb_62 = wdata_io_out_bits_strobe[1]; // @[StreamController.scala 97:28:@95116.4]
  assign io_dram_wdata_bits_wstrb_63 = wdata_io_out_bits_strobe[0]; // @[StreamController.scala 97:28:@95117.4]
  assign io_dram_wresp_ready = wresp_io_in_ready; // @[StreamController.scala 104:23:@95386.4]
  assign io_store_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 79:22:@94886.4]
  assign io_store_data_ready = wdata_io_in_ready; // @[StreamController.scala 93:23:@94915.4]
  assign io_store_wresp_valid = wresp_io_out_valid; // @[StreamController.scala 106:24:@95387.4]
  assign io_store_wresp_bits = wresp_io_out_bits; // @[StreamController.scala 107:23:@95388.4]
  assign cmd_clock = clock; // @[:@94489.4]
  assign cmd_reset = reset; // @[:@94490.4]
  assign cmd_io_in_valid = io_store_cmd_valid; // @[StreamController.scala 77:19:@94883.4]
  assign cmd_io_in_bits_addr = io_store_cmd_bits_addr; // @[StreamController.scala 78:18:@94885.4]
  assign cmd_io_in_bits_size = io_store_cmd_bits_size; // @[StreamController.scala 78:18:@94884.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 80:20:@94887.4]
  assign wdata_clock = clock; // @[:@94895.4]
  assign wdata_reset = reset; // @[:@94896.4]
  assign wdata_io_in_valid = io_store_data_valid; // @[StreamController.scala 90:21:@94912.4]
  assign wdata_io_in_bits_data_0 = io_store_data_bits_wdata_0; // @[StreamController.scala 91:25:@94913.4]
  assign wdata_io_in_bits_strobe = io_store_data_bits_wstrb; // @[StreamController.scala 92:27:@94914.4]
  assign wdata_io_out_ready = io_dram_wdata_ready; // @[StreamController.scala 98:22:@95118.4]
  assign wresp_clock = clock; // @[:@95120.4]
  assign wresp_reset = reset; // @[:@95121.4]
  assign wresp_io_in_valid = io_dram_wresp_valid; // @[StreamController.scala 102:21:@95384.4]
  assign wresp_io_out_ready = io_store_wresp_ready; // @[StreamController.scala 108:22:@95389.4]
endmodule
module MuxN( // @[:@95455.2]
  input  [63:0] io_ins_0_addr, // @[:@95458.4]
  input  [31:0] io_ins_0_size, // @[:@95458.4]
  input         io_ins_0_isWr, // @[:@95458.4]
  input  [31:0] io_ins_0_tag, // @[:@95458.4]
  input  [63:0] io_ins_1_addr, // @[:@95458.4]
  input  [31:0] io_ins_1_size, // @[:@95458.4]
  input         io_ins_1_isWr, // @[:@95458.4]
  input  [31:0] io_ins_1_tag, // @[:@95458.4]
  input         io_sel, // @[:@95458.4]
  output [63:0] io_out_addr, // @[:@95458.4]
  output [31:0] io_out_size, // @[:@95458.4]
  output        io_out_isWr, // @[:@95458.4]
  output [31:0] io_out_tag // @[:@95458.4]
);
  assign io_out_addr = io_sel ? io_ins_1_addr : io_ins_0_addr; // @[MuxN.scala 16:10:@95464.4]
  assign io_out_size = io_sel ? io_ins_1_size : io_ins_0_size; // @[MuxN.scala 16:10:@95463.4]
  assign io_out_isWr = io_sel ? io_ins_1_isWr : io_ins_0_isWr; // @[MuxN.scala 16:10:@95461.4]
  assign io_out_tag = io_sel ? io_ins_1_tag : io_ins_0_tag; // @[MuxN.scala 16:10:@95460.4]
endmodule
module MuxPipe( // @[:@95466.2]
  output        io_in_ready, // @[:@95469.4]
  input         io_in_valid, // @[:@95469.4]
  input  [63:0] io_in_bits_0_addr, // @[:@95469.4]
  input  [31:0] io_in_bits_0_size, // @[:@95469.4]
  input         io_in_bits_0_isWr, // @[:@95469.4]
  input  [31:0] io_in_bits_0_tag, // @[:@95469.4]
  input  [63:0] io_in_bits_1_addr, // @[:@95469.4]
  input  [31:0] io_in_bits_1_size, // @[:@95469.4]
  input         io_in_bits_1_isWr, // @[:@95469.4]
  input  [31:0] io_in_bits_1_tag, // @[:@95469.4]
  input         io_sel, // @[:@95469.4]
  input         io_out_ready, // @[:@95469.4]
  output        io_out_valid, // @[:@95469.4]
  output [63:0] io_out_bits_addr, // @[:@95469.4]
  output [31:0] io_out_bits_size, // @[:@95469.4]
  output        io_out_bits_isWr, // @[:@95469.4]
  output [31:0] io_out_bits_tag // @[:@95469.4]
);
  wire [63:0] MuxN_io_ins_0_addr; // @[MuxN.scala 40:23:@95484.4]
  wire [31:0] MuxN_io_ins_0_size; // @[MuxN.scala 40:23:@95484.4]
  wire  MuxN_io_ins_0_isWr; // @[MuxN.scala 40:23:@95484.4]
  wire [31:0] MuxN_io_ins_0_tag; // @[MuxN.scala 40:23:@95484.4]
  wire [63:0] MuxN_io_ins_1_addr; // @[MuxN.scala 40:23:@95484.4]
  wire [31:0] MuxN_io_ins_1_size; // @[MuxN.scala 40:23:@95484.4]
  wire  MuxN_io_ins_1_isWr; // @[MuxN.scala 40:23:@95484.4]
  wire [31:0] MuxN_io_ins_1_tag; // @[MuxN.scala 40:23:@95484.4]
  wire  MuxN_io_sel; // @[MuxN.scala 40:23:@95484.4]
  wire [63:0] MuxN_io_out_addr; // @[MuxN.scala 40:23:@95484.4]
  wire [31:0] MuxN_io_out_size; // @[MuxN.scala 40:23:@95484.4]
  wire  MuxN_io_out_isWr; // @[MuxN.scala 40:23:@95484.4]
  wire [31:0] MuxN_io_out_tag; // @[MuxN.scala 40:23:@95484.4]
  wire  _T_46; // @[MuxN.scala 28:31:@95471.4]
  MuxN MuxN ( // @[MuxN.scala 40:23:@95484.4]
    .io_ins_0_addr(MuxN_io_ins_0_addr),
    .io_ins_0_size(MuxN_io_ins_0_size),
    .io_ins_0_isWr(MuxN_io_ins_0_isWr),
    .io_ins_0_tag(MuxN_io_ins_0_tag),
    .io_ins_1_addr(MuxN_io_ins_1_addr),
    .io_ins_1_size(MuxN_io_ins_1_size),
    .io_ins_1_isWr(MuxN_io_ins_1_isWr),
    .io_ins_1_tag(MuxN_io_ins_1_tag),
    .io_sel(MuxN_io_sel),
    .io_out_addr(MuxN_io_out_addr),
    .io_out_size(MuxN_io_out_size),
    .io_out_isWr(MuxN_io_out_isWr),
    .io_out_tag(MuxN_io_out_tag)
  );
  assign _T_46 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@95471.4]
  assign io_in_ready = io_out_ready | _T_46; // @[MuxN.scala 71:15:@95500.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@95499.4]
  assign io_out_bits_addr = MuxN_io_out_addr; // @[MuxN.scala 72:15:@95505.4]
  assign io_out_bits_size = MuxN_io_out_size; // @[MuxN.scala 72:15:@95504.4]
  assign io_out_bits_isWr = MuxN_io_out_isWr; // @[MuxN.scala 72:15:@95502.4]
  assign io_out_bits_tag = MuxN_io_out_tag; // @[MuxN.scala 72:15:@95501.4]
  assign MuxN_io_ins_0_addr = io_in_bits_0_addr; // @[MuxN.scala 41:18:@95491.4]
  assign MuxN_io_ins_0_size = io_in_bits_0_size; // @[MuxN.scala 41:18:@95490.4]
  assign MuxN_io_ins_0_isWr = io_in_bits_0_isWr; // @[MuxN.scala 41:18:@95488.4]
  assign MuxN_io_ins_0_tag = io_in_bits_0_tag; // @[MuxN.scala 41:18:@95487.4]
  assign MuxN_io_ins_1_addr = io_in_bits_1_addr; // @[MuxN.scala 41:18:@95496.4]
  assign MuxN_io_ins_1_size = io_in_bits_1_size; // @[MuxN.scala 41:18:@95495.4]
  assign MuxN_io_ins_1_isWr = io_in_bits_1_isWr; // @[MuxN.scala 41:18:@95493.4]
  assign MuxN_io_ins_1_tag = io_in_bits_1_tag; // @[MuxN.scala 41:18:@95492.4]
  assign MuxN_io_sel = io_sel; // @[MuxN.scala 44:18:@95498.4]
endmodule
module MuxN_1( // @[:@95507.2]
  input  [63:0] io_ins_0_wdata_0, // @[:@95510.4]
  input  [63:0] io_ins_0_wdata_1, // @[:@95510.4]
  input  [63:0] io_ins_0_wdata_2, // @[:@95510.4]
  input  [63:0] io_ins_0_wdata_3, // @[:@95510.4]
  input  [63:0] io_ins_0_wdata_4, // @[:@95510.4]
  input  [63:0] io_ins_0_wdata_5, // @[:@95510.4]
  input  [63:0] io_ins_0_wdata_6, // @[:@95510.4]
  input  [63:0] io_ins_0_wdata_7, // @[:@95510.4]
  input         io_ins_0_wstrb_0, // @[:@95510.4]
  input         io_ins_0_wstrb_1, // @[:@95510.4]
  input         io_ins_0_wstrb_2, // @[:@95510.4]
  input         io_ins_0_wstrb_3, // @[:@95510.4]
  input         io_ins_0_wstrb_4, // @[:@95510.4]
  input         io_ins_0_wstrb_5, // @[:@95510.4]
  input         io_ins_0_wstrb_6, // @[:@95510.4]
  input         io_ins_0_wstrb_7, // @[:@95510.4]
  input         io_ins_0_wstrb_8, // @[:@95510.4]
  input         io_ins_0_wstrb_9, // @[:@95510.4]
  input         io_ins_0_wstrb_10, // @[:@95510.4]
  input         io_ins_0_wstrb_11, // @[:@95510.4]
  input         io_ins_0_wstrb_12, // @[:@95510.4]
  input         io_ins_0_wstrb_13, // @[:@95510.4]
  input         io_ins_0_wstrb_14, // @[:@95510.4]
  input         io_ins_0_wstrb_15, // @[:@95510.4]
  input         io_ins_0_wstrb_16, // @[:@95510.4]
  input         io_ins_0_wstrb_17, // @[:@95510.4]
  input         io_ins_0_wstrb_18, // @[:@95510.4]
  input         io_ins_0_wstrb_19, // @[:@95510.4]
  input         io_ins_0_wstrb_20, // @[:@95510.4]
  input         io_ins_0_wstrb_21, // @[:@95510.4]
  input         io_ins_0_wstrb_22, // @[:@95510.4]
  input         io_ins_0_wstrb_23, // @[:@95510.4]
  input         io_ins_0_wstrb_24, // @[:@95510.4]
  input         io_ins_0_wstrb_25, // @[:@95510.4]
  input         io_ins_0_wstrb_26, // @[:@95510.4]
  input         io_ins_0_wstrb_27, // @[:@95510.4]
  input         io_ins_0_wstrb_28, // @[:@95510.4]
  input         io_ins_0_wstrb_29, // @[:@95510.4]
  input         io_ins_0_wstrb_30, // @[:@95510.4]
  input         io_ins_0_wstrb_31, // @[:@95510.4]
  input         io_ins_0_wstrb_32, // @[:@95510.4]
  input         io_ins_0_wstrb_33, // @[:@95510.4]
  input         io_ins_0_wstrb_34, // @[:@95510.4]
  input         io_ins_0_wstrb_35, // @[:@95510.4]
  input         io_ins_0_wstrb_36, // @[:@95510.4]
  input         io_ins_0_wstrb_37, // @[:@95510.4]
  input         io_ins_0_wstrb_38, // @[:@95510.4]
  input         io_ins_0_wstrb_39, // @[:@95510.4]
  input         io_ins_0_wstrb_40, // @[:@95510.4]
  input         io_ins_0_wstrb_41, // @[:@95510.4]
  input         io_ins_0_wstrb_42, // @[:@95510.4]
  input         io_ins_0_wstrb_43, // @[:@95510.4]
  input         io_ins_0_wstrb_44, // @[:@95510.4]
  input         io_ins_0_wstrb_45, // @[:@95510.4]
  input         io_ins_0_wstrb_46, // @[:@95510.4]
  input         io_ins_0_wstrb_47, // @[:@95510.4]
  input         io_ins_0_wstrb_48, // @[:@95510.4]
  input         io_ins_0_wstrb_49, // @[:@95510.4]
  input         io_ins_0_wstrb_50, // @[:@95510.4]
  input         io_ins_0_wstrb_51, // @[:@95510.4]
  input         io_ins_0_wstrb_52, // @[:@95510.4]
  input         io_ins_0_wstrb_53, // @[:@95510.4]
  input         io_ins_0_wstrb_54, // @[:@95510.4]
  input         io_ins_0_wstrb_55, // @[:@95510.4]
  input         io_ins_0_wstrb_56, // @[:@95510.4]
  input         io_ins_0_wstrb_57, // @[:@95510.4]
  input         io_ins_0_wstrb_58, // @[:@95510.4]
  input         io_ins_0_wstrb_59, // @[:@95510.4]
  input         io_ins_0_wstrb_60, // @[:@95510.4]
  input         io_ins_0_wstrb_61, // @[:@95510.4]
  input         io_ins_0_wstrb_62, // @[:@95510.4]
  input         io_ins_0_wstrb_63, // @[:@95510.4]
  input  [63:0] io_ins_1_wdata_0, // @[:@95510.4]
  input  [63:0] io_ins_1_wdata_1, // @[:@95510.4]
  input  [63:0] io_ins_1_wdata_2, // @[:@95510.4]
  input  [63:0] io_ins_1_wdata_3, // @[:@95510.4]
  input  [63:0] io_ins_1_wdata_4, // @[:@95510.4]
  input  [63:0] io_ins_1_wdata_5, // @[:@95510.4]
  input  [63:0] io_ins_1_wdata_6, // @[:@95510.4]
  input  [63:0] io_ins_1_wdata_7, // @[:@95510.4]
  input         io_ins_1_wstrb_0, // @[:@95510.4]
  input         io_ins_1_wstrb_1, // @[:@95510.4]
  input         io_ins_1_wstrb_2, // @[:@95510.4]
  input         io_ins_1_wstrb_3, // @[:@95510.4]
  input         io_ins_1_wstrb_4, // @[:@95510.4]
  input         io_ins_1_wstrb_5, // @[:@95510.4]
  input         io_ins_1_wstrb_6, // @[:@95510.4]
  input         io_ins_1_wstrb_7, // @[:@95510.4]
  input         io_ins_1_wstrb_8, // @[:@95510.4]
  input         io_ins_1_wstrb_9, // @[:@95510.4]
  input         io_ins_1_wstrb_10, // @[:@95510.4]
  input         io_ins_1_wstrb_11, // @[:@95510.4]
  input         io_ins_1_wstrb_12, // @[:@95510.4]
  input         io_ins_1_wstrb_13, // @[:@95510.4]
  input         io_ins_1_wstrb_14, // @[:@95510.4]
  input         io_ins_1_wstrb_15, // @[:@95510.4]
  input         io_ins_1_wstrb_16, // @[:@95510.4]
  input         io_ins_1_wstrb_17, // @[:@95510.4]
  input         io_ins_1_wstrb_18, // @[:@95510.4]
  input         io_ins_1_wstrb_19, // @[:@95510.4]
  input         io_ins_1_wstrb_20, // @[:@95510.4]
  input         io_ins_1_wstrb_21, // @[:@95510.4]
  input         io_ins_1_wstrb_22, // @[:@95510.4]
  input         io_ins_1_wstrb_23, // @[:@95510.4]
  input         io_ins_1_wstrb_24, // @[:@95510.4]
  input         io_ins_1_wstrb_25, // @[:@95510.4]
  input         io_ins_1_wstrb_26, // @[:@95510.4]
  input         io_ins_1_wstrb_27, // @[:@95510.4]
  input         io_ins_1_wstrb_28, // @[:@95510.4]
  input         io_ins_1_wstrb_29, // @[:@95510.4]
  input         io_ins_1_wstrb_30, // @[:@95510.4]
  input         io_ins_1_wstrb_31, // @[:@95510.4]
  input         io_ins_1_wstrb_32, // @[:@95510.4]
  input         io_ins_1_wstrb_33, // @[:@95510.4]
  input         io_ins_1_wstrb_34, // @[:@95510.4]
  input         io_ins_1_wstrb_35, // @[:@95510.4]
  input         io_ins_1_wstrb_36, // @[:@95510.4]
  input         io_ins_1_wstrb_37, // @[:@95510.4]
  input         io_ins_1_wstrb_38, // @[:@95510.4]
  input         io_ins_1_wstrb_39, // @[:@95510.4]
  input         io_ins_1_wstrb_40, // @[:@95510.4]
  input         io_ins_1_wstrb_41, // @[:@95510.4]
  input         io_ins_1_wstrb_42, // @[:@95510.4]
  input         io_ins_1_wstrb_43, // @[:@95510.4]
  input         io_ins_1_wstrb_44, // @[:@95510.4]
  input         io_ins_1_wstrb_45, // @[:@95510.4]
  input         io_ins_1_wstrb_46, // @[:@95510.4]
  input         io_ins_1_wstrb_47, // @[:@95510.4]
  input         io_ins_1_wstrb_48, // @[:@95510.4]
  input         io_ins_1_wstrb_49, // @[:@95510.4]
  input         io_ins_1_wstrb_50, // @[:@95510.4]
  input         io_ins_1_wstrb_51, // @[:@95510.4]
  input         io_ins_1_wstrb_52, // @[:@95510.4]
  input         io_ins_1_wstrb_53, // @[:@95510.4]
  input         io_ins_1_wstrb_54, // @[:@95510.4]
  input         io_ins_1_wstrb_55, // @[:@95510.4]
  input         io_ins_1_wstrb_56, // @[:@95510.4]
  input         io_ins_1_wstrb_57, // @[:@95510.4]
  input         io_ins_1_wstrb_58, // @[:@95510.4]
  input         io_ins_1_wstrb_59, // @[:@95510.4]
  input         io_ins_1_wstrb_60, // @[:@95510.4]
  input         io_ins_1_wstrb_61, // @[:@95510.4]
  input         io_ins_1_wstrb_62, // @[:@95510.4]
  input         io_ins_1_wstrb_63, // @[:@95510.4]
  input         io_sel, // @[:@95510.4]
  output [63:0] io_out_wdata_0, // @[:@95510.4]
  output [63:0] io_out_wdata_1, // @[:@95510.4]
  output [63:0] io_out_wdata_2, // @[:@95510.4]
  output [63:0] io_out_wdata_3, // @[:@95510.4]
  output [63:0] io_out_wdata_4, // @[:@95510.4]
  output [63:0] io_out_wdata_5, // @[:@95510.4]
  output [63:0] io_out_wdata_6, // @[:@95510.4]
  output [63:0] io_out_wdata_7, // @[:@95510.4]
  output        io_out_wstrb_0, // @[:@95510.4]
  output        io_out_wstrb_1, // @[:@95510.4]
  output        io_out_wstrb_2, // @[:@95510.4]
  output        io_out_wstrb_3, // @[:@95510.4]
  output        io_out_wstrb_4, // @[:@95510.4]
  output        io_out_wstrb_5, // @[:@95510.4]
  output        io_out_wstrb_6, // @[:@95510.4]
  output        io_out_wstrb_7, // @[:@95510.4]
  output        io_out_wstrb_8, // @[:@95510.4]
  output        io_out_wstrb_9, // @[:@95510.4]
  output        io_out_wstrb_10, // @[:@95510.4]
  output        io_out_wstrb_11, // @[:@95510.4]
  output        io_out_wstrb_12, // @[:@95510.4]
  output        io_out_wstrb_13, // @[:@95510.4]
  output        io_out_wstrb_14, // @[:@95510.4]
  output        io_out_wstrb_15, // @[:@95510.4]
  output        io_out_wstrb_16, // @[:@95510.4]
  output        io_out_wstrb_17, // @[:@95510.4]
  output        io_out_wstrb_18, // @[:@95510.4]
  output        io_out_wstrb_19, // @[:@95510.4]
  output        io_out_wstrb_20, // @[:@95510.4]
  output        io_out_wstrb_21, // @[:@95510.4]
  output        io_out_wstrb_22, // @[:@95510.4]
  output        io_out_wstrb_23, // @[:@95510.4]
  output        io_out_wstrb_24, // @[:@95510.4]
  output        io_out_wstrb_25, // @[:@95510.4]
  output        io_out_wstrb_26, // @[:@95510.4]
  output        io_out_wstrb_27, // @[:@95510.4]
  output        io_out_wstrb_28, // @[:@95510.4]
  output        io_out_wstrb_29, // @[:@95510.4]
  output        io_out_wstrb_30, // @[:@95510.4]
  output        io_out_wstrb_31, // @[:@95510.4]
  output        io_out_wstrb_32, // @[:@95510.4]
  output        io_out_wstrb_33, // @[:@95510.4]
  output        io_out_wstrb_34, // @[:@95510.4]
  output        io_out_wstrb_35, // @[:@95510.4]
  output        io_out_wstrb_36, // @[:@95510.4]
  output        io_out_wstrb_37, // @[:@95510.4]
  output        io_out_wstrb_38, // @[:@95510.4]
  output        io_out_wstrb_39, // @[:@95510.4]
  output        io_out_wstrb_40, // @[:@95510.4]
  output        io_out_wstrb_41, // @[:@95510.4]
  output        io_out_wstrb_42, // @[:@95510.4]
  output        io_out_wstrb_43, // @[:@95510.4]
  output        io_out_wstrb_44, // @[:@95510.4]
  output        io_out_wstrb_45, // @[:@95510.4]
  output        io_out_wstrb_46, // @[:@95510.4]
  output        io_out_wstrb_47, // @[:@95510.4]
  output        io_out_wstrb_48, // @[:@95510.4]
  output        io_out_wstrb_49, // @[:@95510.4]
  output        io_out_wstrb_50, // @[:@95510.4]
  output        io_out_wstrb_51, // @[:@95510.4]
  output        io_out_wstrb_52, // @[:@95510.4]
  output        io_out_wstrb_53, // @[:@95510.4]
  output        io_out_wstrb_54, // @[:@95510.4]
  output        io_out_wstrb_55, // @[:@95510.4]
  output        io_out_wstrb_56, // @[:@95510.4]
  output        io_out_wstrb_57, // @[:@95510.4]
  output        io_out_wstrb_58, // @[:@95510.4]
  output        io_out_wstrb_59, // @[:@95510.4]
  output        io_out_wstrb_60, // @[:@95510.4]
  output        io_out_wstrb_61, // @[:@95510.4]
  output        io_out_wstrb_62, // @[:@95510.4]
  output        io_out_wstrb_63 // @[:@95510.4]
);
  assign io_out_wdata_0 = io_sel ? io_ins_1_wdata_0 : io_ins_0_wdata_0; // @[MuxN.scala 16:10:@95577.4]
  assign io_out_wdata_1 = io_sel ? io_ins_1_wdata_1 : io_ins_0_wdata_1; // @[MuxN.scala 16:10:@95578.4]
  assign io_out_wdata_2 = io_sel ? io_ins_1_wdata_2 : io_ins_0_wdata_2; // @[MuxN.scala 16:10:@95579.4]
  assign io_out_wdata_3 = io_sel ? io_ins_1_wdata_3 : io_ins_0_wdata_3; // @[MuxN.scala 16:10:@95580.4]
  assign io_out_wdata_4 = io_sel ? io_ins_1_wdata_4 : io_ins_0_wdata_4; // @[MuxN.scala 16:10:@95581.4]
  assign io_out_wdata_5 = io_sel ? io_ins_1_wdata_5 : io_ins_0_wdata_5; // @[MuxN.scala 16:10:@95582.4]
  assign io_out_wdata_6 = io_sel ? io_ins_1_wdata_6 : io_ins_0_wdata_6; // @[MuxN.scala 16:10:@95583.4]
  assign io_out_wdata_7 = io_sel ? io_ins_1_wdata_7 : io_ins_0_wdata_7; // @[MuxN.scala 16:10:@95584.4]
  assign io_out_wstrb_0 = io_sel ? io_ins_1_wstrb_0 : io_ins_0_wstrb_0; // @[MuxN.scala 16:10:@95513.4]
  assign io_out_wstrb_1 = io_sel ? io_ins_1_wstrb_1 : io_ins_0_wstrb_1; // @[MuxN.scala 16:10:@95514.4]
  assign io_out_wstrb_2 = io_sel ? io_ins_1_wstrb_2 : io_ins_0_wstrb_2; // @[MuxN.scala 16:10:@95515.4]
  assign io_out_wstrb_3 = io_sel ? io_ins_1_wstrb_3 : io_ins_0_wstrb_3; // @[MuxN.scala 16:10:@95516.4]
  assign io_out_wstrb_4 = io_sel ? io_ins_1_wstrb_4 : io_ins_0_wstrb_4; // @[MuxN.scala 16:10:@95517.4]
  assign io_out_wstrb_5 = io_sel ? io_ins_1_wstrb_5 : io_ins_0_wstrb_5; // @[MuxN.scala 16:10:@95518.4]
  assign io_out_wstrb_6 = io_sel ? io_ins_1_wstrb_6 : io_ins_0_wstrb_6; // @[MuxN.scala 16:10:@95519.4]
  assign io_out_wstrb_7 = io_sel ? io_ins_1_wstrb_7 : io_ins_0_wstrb_7; // @[MuxN.scala 16:10:@95520.4]
  assign io_out_wstrb_8 = io_sel ? io_ins_1_wstrb_8 : io_ins_0_wstrb_8; // @[MuxN.scala 16:10:@95521.4]
  assign io_out_wstrb_9 = io_sel ? io_ins_1_wstrb_9 : io_ins_0_wstrb_9; // @[MuxN.scala 16:10:@95522.4]
  assign io_out_wstrb_10 = io_sel ? io_ins_1_wstrb_10 : io_ins_0_wstrb_10; // @[MuxN.scala 16:10:@95523.4]
  assign io_out_wstrb_11 = io_sel ? io_ins_1_wstrb_11 : io_ins_0_wstrb_11; // @[MuxN.scala 16:10:@95524.4]
  assign io_out_wstrb_12 = io_sel ? io_ins_1_wstrb_12 : io_ins_0_wstrb_12; // @[MuxN.scala 16:10:@95525.4]
  assign io_out_wstrb_13 = io_sel ? io_ins_1_wstrb_13 : io_ins_0_wstrb_13; // @[MuxN.scala 16:10:@95526.4]
  assign io_out_wstrb_14 = io_sel ? io_ins_1_wstrb_14 : io_ins_0_wstrb_14; // @[MuxN.scala 16:10:@95527.4]
  assign io_out_wstrb_15 = io_sel ? io_ins_1_wstrb_15 : io_ins_0_wstrb_15; // @[MuxN.scala 16:10:@95528.4]
  assign io_out_wstrb_16 = io_sel ? io_ins_1_wstrb_16 : io_ins_0_wstrb_16; // @[MuxN.scala 16:10:@95529.4]
  assign io_out_wstrb_17 = io_sel ? io_ins_1_wstrb_17 : io_ins_0_wstrb_17; // @[MuxN.scala 16:10:@95530.4]
  assign io_out_wstrb_18 = io_sel ? io_ins_1_wstrb_18 : io_ins_0_wstrb_18; // @[MuxN.scala 16:10:@95531.4]
  assign io_out_wstrb_19 = io_sel ? io_ins_1_wstrb_19 : io_ins_0_wstrb_19; // @[MuxN.scala 16:10:@95532.4]
  assign io_out_wstrb_20 = io_sel ? io_ins_1_wstrb_20 : io_ins_0_wstrb_20; // @[MuxN.scala 16:10:@95533.4]
  assign io_out_wstrb_21 = io_sel ? io_ins_1_wstrb_21 : io_ins_0_wstrb_21; // @[MuxN.scala 16:10:@95534.4]
  assign io_out_wstrb_22 = io_sel ? io_ins_1_wstrb_22 : io_ins_0_wstrb_22; // @[MuxN.scala 16:10:@95535.4]
  assign io_out_wstrb_23 = io_sel ? io_ins_1_wstrb_23 : io_ins_0_wstrb_23; // @[MuxN.scala 16:10:@95536.4]
  assign io_out_wstrb_24 = io_sel ? io_ins_1_wstrb_24 : io_ins_0_wstrb_24; // @[MuxN.scala 16:10:@95537.4]
  assign io_out_wstrb_25 = io_sel ? io_ins_1_wstrb_25 : io_ins_0_wstrb_25; // @[MuxN.scala 16:10:@95538.4]
  assign io_out_wstrb_26 = io_sel ? io_ins_1_wstrb_26 : io_ins_0_wstrb_26; // @[MuxN.scala 16:10:@95539.4]
  assign io_out_wstrb_27 = io_sel ? io_ins_1_wstrb_27 : io_ins_0_wstrb_27; // @[MuxN.scala 16:10:@95540.4]
  assign io_out_wstrb_28 = io_sel ? io_ins_1_wstrb_28 : io_ins_0_wstrb_28; // @[MuxN.scala 16:10:@95541.4]
  assign io_out_wstrb_29 = io_sel ? io_ins_1_wstrb_29 : io_ins_0_wstrb_29; // @[MuxN.scala 16:10:@95542.4]
  assign io_out_wstrb_30 = io_sel ? io_ins_1_wstrb_30 : io_ins_0_wstrb_30; // @[MuxN.scala 16:10:@95543.4]
  assign io_out_wstrb_31 = io_sel ? io_ins_1_wstrb_31 : io_ins_0_wstrb_31; // @[MuxN.scala 16:10:@95544.4]
  assign io_out_wstrb_32 = io_sel ? io_ins_1_wstrb_32 : io_ins_0_wstrb_32; // @[MuxN.scala 16:10:@95545.4]
  assign io_out_wstrb_33 = io_sel ? io_ins_1_wstrb_33 : io_ins_0_wstrb_33; // @[MuxN.scala 16:10:@95546.4]
  assign io_out_wstrb_34 = io_sel ? io_ins_1_wstrb_34 : io_ins_0_wstrb_34; // @[MuxN.scala 16:10:@95547.4]
  assign io_out_wstrb_35 = io_sel ? io_ins_1_wstrb_35 : io_ins_0_wstrb_35; // @[MuxN.scala 16:10:@95548.4]
  assign io_out_wstrb_36 = io_sel ? io_ins_1_wstrb_36 : io_ins_0_wstrb_36; // @[MuxN.scala 16:10:@95549.4]
  assign io_out_wstrb_37 = io_sel ? io_ins_1_wstrb_37 : io_ins_0_wstrb_37; // @[MuxN.scala 16:10:@95550.4]
  assign io_out_wstrb_38 = io_sel ? io_ins_1_wstrb_38 : io_ins_0_wstrb_38; // @[MuxN.scala 16:10:@95551.4]
  assign io_out_wstrb_39 = io_sel ? io_ins_1_wstrb_39 : io_ins_0_wstrb_39; // @[MuxN.scala 16:10:@95552.4]
  assign io_out_wstrb_40 = io_sel ? io_ins_1_wstrb_40 : io_ins_0_wstrb_40; // @[MuxN.scala 16:10:@95553.4]
  assign io_out_wstrb_41 = io_sel ? io_ins_1_wstrb_41 : io_ins_0_wstrb_41; // @[MuxN.scala 16:10:@95554.4]
  assign io_out_wstrb_42 = io_sel ? io_ins_1_wstrb_42 : io_ins_0_wstrb_42; // @[MuxN.scala 16:10:@95555.4]
  assign io_out_wstrb_43 = io_sel ? io_ins_1_wstrb_43 : io_ins_0_wstrb_43; // @[MuxN.scala 16:10:@95556.4]
  assign io_out_wstrb_44 = io_sel ? io_ins_1_wstrb_44 : io_ins_0_wstrb_44; // @[MuxN.scala 16:10:@95557.4]
  assign io_out_wstrb_45 = io_sel ? io_ins_1_wstrb_45 : io_ins_0_wstrb_45; // @[MuxN.scala 16:10:@95558.4]
  assign io_out_wstrb_46 = io_sel ? io_ins_1_wstrb_46 : io_ins_0_wstrb_46; // @[MuxN.scala 16:10:@95559.4]
  assign io_out_wstrb_47 = io_sel ? io_ins_1_wstrb_47 : io_ins_0_wstrb_47; // @[MuxN.scala 16:10:@95560.4]
  assign io_out_wstrb_48 = io_sel ? io_ins_1_wstrb_48 : io_ins_0_wstrb_48; // @[MuxN.scala 16:10:@95561.4]
  assign io_out_wstrb_49 = io_sel ? io_ins_1_wstrb_49 : io_ins_0_wstrb_49; // @[MuxN.scala 16:10:@95562.4]
  assign io_out_wstrb_50 = io_sel ? io_ins_1_wstrb_50 : io_ins_0_wstrb_50; // @[MuxN.scala 16:10:@95563.4]
  assign io_out_wstrb_51 = io_sel ? io_ins_1_wstrb_51 : io_ins_0_wstrb_51; // @[MuxN.scala 16:10:@95564.4]
  assign io_out_wstrb_52 = io_sel ? io_ins_1_wstrb_52 : io_ins_0_wstrb_52; // @[MuxN.scala 16:10:@95565.4]
  assign io_out_wstrb_53 = io_sel ? io_ins_1_wstrb_53 : io_ins_0_wstrb_53; // @[MuxN.scala 16:10:@95566.4]
  assign io_out_wstrb_54 = io_sel ? io_ins_1_wstrb_54 : io_ins_0_wstrb_54; // @[MuxN.scala 16:10:@95567.4]
  assign io_out_wstrb_55 = io_sel ? io_ins_1_wstrb_55 : io_ins_0_wstrb_55; // @[MuxN.scala 16:10:@95568.4]
  assign io_out_wstrb_56 = io_sel ? io_ins_1_wstrb_56 : io_ins_0_wstrb_56; // @[MuxN.scala 16:10:@95569.4]
  assign io_out_wstrb_57 = io_sel ? io_ins_1_wstrb_57 : io_ins_0_wstrb_57; // @[MuxN.scala 16:10:@95570.4]
  assign io_out_wstrb_58 = io_sel ? io_ins_1_wstrb_58 : io_ins_0_wstrb_58; // @[MuxN.scala 16:10:@95571.4]
  assign io_out_wstrb_59 = io_sel ? io_ins_1_wstrb_59 : io_ins_0_wstrb_59; // @[MuxN.scala 16:10:@95572.4]
  assign io_out_wstrb_60 = io_sel ? io_ins_1_wstrb_60 : io_ins_0_wstrb_60; // @[MuxN.scala 16:10:@95573.4]
  assign io_out_wstrb_61 = io_sel ? io_ins_1_wstrb_61 : io_ins_0_wstrb_61; // @[MuxN.scala 16:10:@95574.4]
  assign io_out_wstrb_62 = io_sel ? io_ins_1_wstrb_62 : io_ins_0_wstrb_62; // @[MuxN.scala 16:10:@95575.4]
  assign io_out_wstrb_63 = io_sel ? io_ins_1_wstrb_63 : io_ins_0_wstrb_63; // @[MuxN.scala 16:10:@95576.4]
endmodule
module MuxPipe_1( // @[:@95586.2]
  output        io_in_ready, // @[:@95589.4]
  input         io_in_valid, // @[:@95589.4]
  input  [63:0] io_in_bits_0_wdata_0, // @[:@95589.4]
  input  [63:0] io_in_bits_0_wdata_1, // @[:@95589.4]
  input  [63:0] io_in_bits_0_wdata_2, // @[:@95589.4]
  input  [63:0] io_in_bits_0_wdata_3, // @[:@95589.4]
  input  [63:0] io_in_bits_0_wdata_4, // @[:@95589.4]
  input  [63:0] io_in_bits_0_wdata_5, // @[:@95589.4]
  input  [63:0] io_in_bits_0_wdata_6, // @[:@95589.4]
  input  [63:0] io_in_bits_0_wdata_7, // @[:@95589.4]
  input         io_in_bits_0_wstrb_0, // @[:@95589.4]
  input         io_in_bits_0_wstrb_1, // @[:@95589.4]
  input         io_in_bits_0_wstrb_2, // @[:@95589.4]
  input         io_in_bits_0_wstrb_3, // @[:@95589.4]
  input         io_in_bits_0_wstrb_4, // @[:@95589.4]
  input         io_in_bits_0_wstrb_5, // @[:@95589.4]
  input         io_in_bits_0_wstrb_6, // @[:@95589.4]
  input         io_in_bits_0_wstrb_7, // @[:@95589.4]
  input         io_in_bits_0_wstrb_8, // @[:@95589.4]
  input         io_in_bits_0_wstrb_9, // @[:@95589.4]
  input         io_in_bits_0_wstrb_10, // @[:@95589.4]
  input         io_in_bits_0_wstrb_11, // @[:@95589.4]
  input         io_in_bits_0_wstrb_12, // @[:@95589.4]
  input         io_in_bits_0_wstrb_13, // @[:@95589.4]
  input         io_in_bits_0_wstrb_14, // @[:@95589.4]
  input         io_in_bits_0_wstrb_15, // @[:@95589.4]
  input         io_in_bits_0_wstrb_16, // @[:@95589.4]
  input         io_in_bits_0_wstrb_17, // @[:@95589.4]
  input         io_in_bits_0_wstrb_18, // @[:@95589.4]
  input         io_in_bits_0_wstrb_19, // @[:@95589.4]
  input         io_in_bits_0_wstrb_20, // @[:@95589.4]
  input         io_in_bits_0_wstrb_21, // @[:@95589.4]
  input         io_in_bits_0_wstrb_22, // @[:@95589.4]
  input         io_in_bits_0_wstrb_23, // @[:@95589.4]
  input         io_in_bits_0_wstrb_24, // @[:@95589.4]
  input         io_in_bits_0_wstrb_25, // @[:@95589.4]
  input         io_in_bits_0_wstrb_26, // @[:@95589.4]
  input         io_in_bits_0_wstrb_27, // @[:@95589.4]
  input         io_in_bits_0_wstrb_28, // @[:@95589.4]
  input         io_in_bits_0_wstrb_29, // @[:@95589.4]
  input         io_in_bits_0_wstrb_30, // @[:@95589.4]
  input         io_in_bits_0_wstrb_31, // @[:@95589.4]
  input         io_in_bits_0_wstrb_32, // @[:@95589.4]
  input         io_in_bits_0_wstrb_33, // @[:@95589.4]
  input         io_in_bits_0_wstrb_34, // @[:@95589.4]
  input         io_in_bits_0_wstrb_35, // @[:@95589.4]
  input         io_in_bits_0_wstrb_36, // @[:@95589.4]
  input         io_in_bits_0_wstrb_37, // @[:@95589.4]
  input         io_in_bits_0_wstrb_38, // @[:@95589.4]
  input         io_in_bits_0_wstrb_39, // @[:@95589.4]
  input         io_in_bits_0_wstrb_40, // @[:@95589.4]
  input         io_in_bits_0_wstrb_41, // @[:@95589.4]
  input         io_in_bits_0_wstrb_42, // @[:@95589.4]
  input         io_in_bits_0_wstrb_43, // @[:@95589.4]
  input         io_in_bits_0_wstrb_44, // @[:@95589.4]
  input         io_in_bits_0_wstrb_45, // @[:@95589.4]
  input         io_in_bits_0_wstrb_46, // @[:@95589.4]
  input         io_in_bits_0_wstrb_47, // @[:@95589.4]
  input         io_in_bits_0_wstrb_48, // @[:@95589.4]
  input         io_in_bits_0_wstrb_49, // @[:@95589.4]
  input         io_in_bits_0_wstrb_50, // @[:@95589.4]
  input         io_in_bits_0_wstrb_51, // @[:@95589.4]
  input         io_in_bits_0_wstrb_52, // @[:@95589.4]
  input         io_in_bits_0_wstrb_53, // @[:@95589.4]
  input         io_in_bits_0_wstrb_54, // @[:@95589.4]
  input         io_in_bits_0_wstrb_55, // @[:@95589.4]
  input         io_in_bits_0_wstrb_56, // @[:@95589.4]
  input         io_in_bits_0_wstrb_57, // @[:@95589.4]
  input         io_in_bits_0_wstrb_58, // @[:@95589.4]
  input         io_in_bits_0_wstrb_59, // @[:@95589.4]
  input         io_in_bits_0_wstrb_60, // @[:@95589.4]
  input         io_in_bits_0_wstrb_61, // @[:@95589.4]
  input         io_in_bits_0_wstrb_62, // @[:@95589.4]
  input         io_in_bits_0_wstrb_63, // @[:@95589.4]
  input  [63:0] io_in_bits_1_wdata_0, // @[:@95589.4]
  input  [63:0] io_in_bits_1_wdata_1, // @[:@95589.4]
  input  [63:0] io_in_bits_1_wdata_2, // @[:@95589.4]
  input  [63:0] io_in_bits_1_wdata_3, // @[:@95589.4]
  input  [63:0] io_in_bits_1_wdata_4, // @[:@95589.4]
  input  [63:0] io_in_bits_1_wdata_5, // @[:@95589.4]
  input  [63:0] io_in_bits_1_wdata_6, // @[:@95589.4]
  input  [63:0] io_in_bits_1_wdata_7, // @[:@95589.4]
  input         io_in_bits_1_wstrb_0, // @[:@95589.4]
  input         io_in_bits_1_wstrb_1, // @[:@95589.4]
  input         io_in_bits_1_wstrb_2, // @[:@95589.4]
  input         io_in_bits_1_wstrb_3, // @[:@95589.4]
  input         io_in_bits_1_wstrb_4, // @[:@95589.4]
  input         io_in_bits_1_wstrb_5, // @[:@95589.4]
  input         io_in_bits_1_wstrb_6, // @[:@95589.4]
  input         io_in_bits_1_wstrb_7, // @[:@95589.4]
  input         io_in_bits_1_wstrb_8, // @[:@95589.4]
  input         io_in_bits_1_wstrb_9, // @[:@95589.4]
  input         io_in_bits_1_wstrb_10, // @[:@95589.4]
  input         io_in_bits_1_wstrb_11, // @[:@95589.4]
  input         io_in_bits_1_wstrb_12, // @[:@95589.4]
  input         io_in_bits_1_wstrb_13, // @[:@95589.4]
  input         io_in_bits_1_wstrb_14, // @[:@95589.4]
  input         io_in_bits_1_wstrb_15, // @[:@95589.4]
  input         io_in_bits_1_wstrb_16, // @[:@95589.4]
  input         io_in_bits_1_wstrb_17, // @[:@95589.4]
  input         io_in_bits_1_wstrb_18, // @[:@95589.4]
  input         io_in_bits_1_wstrb_19, // @[:@95589.4]
  input         io_in_bits_1_wstrb_20, // @[:@95589.4]
  input         io_in_bits_1_wstrb_21, // @[:@95589.4]
  input         io_in_bits_1_wstrb_22, // @[:@95589.4]
  input         io_in_bits_1_wstrb_23, // @[:@95589.4]
  input         io_in_bits_1_wstrb_24, // @[:@95589.4]
  input         io_in_bits_1_wstrb_25, // @[:@95589.4]
  input         io_in_bits_1_wstrb_26, // @[:@95589.4]
  input         io_in_bits_1_wstrb_27, // @[:@95589.4]
  input         io_in_bits_1_wstrb_28, // @[:@95589.4]
  input         io_in_bits_1_wstrb_29, // @[:@95589.4]
  input         io_in_bits_1_wstrb_30, // @[:@95589.4]
  input         io_in_bits_1_wstrb_31, // @[:@95589.4]
  input         io_in_bits_1_wstrb_32, // @[:@95589.4]
  input         io_in_bits_1_wstrb_33, // @[:@95589.4]
  input         io_in_bits_1_wstrb_34, // @[:@95589.4]
  input         io_in_bits_1_wstrb_35, // @[:@95589.4]
  input         io_in_bits_1_wstrb_36, // @[:@95589.4]
  input         io_in_bits_1_wstrb_37, // @[:@95589.4]
  input         io_in_bits_1_wstrb_38, // @[:@95589.4]
  input         io_in_bits_1_wstrb_39, // @[:@95589.4]
  input         io_in_bits_1_wstrb_40, // @[:@95589.4]
  input         io_in_bits_1_wstrb_41, // @[:@95589.4]
  input         io_in_bits_1_wstrb_42, // @[:@95589.4]
  input         io_in_bits_1_wstrb_43, // @[:@95589.4]
  input         io_in_bits_1_wstrb_44, // @[:@95589.4]
  input         io_in_bits_1_wstrb_45, // @[:@95589.4]
  input         io_in_bits_1_wstrb_46, // @[:@95589.4]
  input         io_in_bits_1_wstrb_47, // @[:@95589.4]
  input         io_in_bits_1_wstrb_48, // @[:@95589.4]
  input         io_in_bits_1_wstrb_49, // @[:@95589.4]
  input         io_in_bits_1_wstrb_50, // @[:@95589.4]
  input         io_in_bits_1_wstrb_51, // @[:@95589.4]
  input         io_in_bits_1_wstrb_52, // @[:@95589.4]
  input         io_in_bits_1_wstrb_53, // @[:@95589.4]
  input         io_in_bits_1_wstrb_54, // @[:@95589.4]
  input         io_in_bits_1_wstrb_55, // @[:@95589.4]
  input         io_in_bits_1_wstrb_56, // @[:@95589.4]
  input         io_in_bits_1_wstrb_57, // @[:@95589.4]
  input         io_in_bits_1_wstrb_58, // @[:@95589.4]
  input         io_in_bits_1_wstrb_59, // @[:@95589.4]
  input         io_in_bits_1_wstrb_60, // @[:@95589.4]
  input         io_in_bits_1_wstrb_61, // @[:@95589.4]
  input         io_in_bits_1_wstrb_62, // @[:@95589.4]
  input         io_in_bits_1_wstrb_63, // @[:@95589.4]
  input         io_sel, // @[:@95589.4]
  input         io_out_ready, // @[:@95589.4]
  output        io_out_valid, // @[:@95589.4]
  output [63:0] io_out_bits_wdata_0, // @[:@95589.4]
  output [63:0] io_out_bits_wdata_1, // @[:@95589.4]
  output [63:0] io_out_bits_wdata_2, // @[:@95589.4]
  output [63:0] io_out_bits_wdata_3, // @[:@95589.4]
  output [63:0] io_out_bits_wdata_4, // @[:@95589.4]
  output [63:0] io_out_bits_wdata_5, // @[:@95589.4]
  output [63:0] io_out_bits_wdata_6, // @[:@95589.4]
  output [63:0] io_out_bits_wdata_7, // @[:@95589.4]
  output        io_out_bits_wstrb_0, // @[:@95589.4]
  output        io_out_bits_wstrb_1, // @[:@95589.4]
  output        io_out_bits_wstrb_2, // @[:@95589.4]
  output        io_out_bits_wstrb_3, // @[:@95589.4]
  output        io_out_bits_wstrb_4, // @[:@95589.4]
  output        io_out_bits_wstrb_5, // @[:@95589.4]
  output        io_out_bits_wstrb_6, // @[:@95589.4]
  output        io_out_bits_wstrb_7, // @[:@95589.4]
  output        io_out_bits_wstrb_8, // @[:@95589.4]
  output        io_out_bits_wstrb_9, // @[:@95589.4]
  output        io_out_bits_wstrb_10, // @[:@95589.4]
  output        io_out_bits_wstrb_11, // @[:@95589.4]
  output        io_out_bits_wstrb_12, // @[:@95589.4]
  output        io_out_bits_wstrb_13, // @[:@95589.4]
  output        io_out_bits_wstrb_14, // @[:@95589.4]
  output        io_out_bits_wstrb_15, // @[:@95589.4]
  output        io_out_bits_wstrb_16, // @[:@95589.4]
  output        io_out_bits_wstrb_17, // @[:@95589.4]
  output        io_out_bits_wstrb_18, // @[:@95589.4]
  output        io_out_bits_wstrb_19, // @[:@95589.4]
  output        io_out_bits_wstrb_20, // @[:@95589.4]
  output        io_out_bits_wstrb_21, // @[:@95589.4]
  output        io_out_bits_wstrb_22, // @[:@95589.4]
  output        io_out_bits_wstrb_23, // @[:@95589.4]
  output        io_out_bits_wstrb_24, // @[:@95589.4]
  output        io_out_bits_wstrb_25, // @[:@95589.4]
  output        io_out_bits_wstrb_26, // @[:@95589.4]
  output        io_out_bits_wstrb_27, // @[:@95589.4]
  output        io_out_bits_wstrb_28, // @[:@95589.4]
  output        io_out_bits_wstrb_29, // @[:@95589.4]
  output        io_out_bits_wstrb_30, // @[:@95589.4]
  output        io_out_bits_wstrb_31, // @[:@95589.4]
  output        io_out_bits_wstrb_32, // @[:@95589.4]
  output        io_out_bits_wstrb_33, // @[:@95589.4]
  output        io_out_bits_wstrb_34, // @[:@95589.4]
  output        io_out_bits_wstrb_35, // @[:@95589.4]
  output        io_out_bits_wstrb_36, // @[:@95589.4]
  output        io_out_bits_wstrb_37, // @[:@95589.4]
  output        io_out_bits_wstrb_38, // @[:@95589.4]
  output        io_out_bits_wstrb_39, // @[:@95589.4]
  output        io_out_bits_wstrb_40, // @[:@95589.4]
  output        io_out_bits_wstrb_41, // @[:@95589.4]
  output        io_out_bits_wstrb_42, // @[:@95589.4]
  output        io_out_bits_wstrb_43, // @[:@95589.4]
  output        io_out_bits_wstrb_44, // @[:@95589.4]
  output        io_out_bits_wstrb_45, // @[:@95589.4]
  output        io_out_bits_wstrb_46, // @[:@95589.4]
  output        io_out_bits_wstrb_47, // @[:@95589.4]
  output        io_out_bits_wstrb_48, // @[:@95589.4]
  output        io_out_bits_wstrb_49, // @[:@95589.4]
  output        io_out_bits_wstrb_50, // @[:@95589.4]
  output        io_out_bits_wstrb_51, // @[:@95589.4]
  output        io_out_bits_wstrb_52, // @[:@95589.4]
  output        io_out_bits_wstrb_53, // @[:@95589.4]
  output        io_out_bits_wstrb_54, // @[:@95589.4]
  output        io_out_bits_wstrb_55, // @[:@95589.4]
  output        io_out_bits_wstrb_56, // @[:@95589.4]
  output        io_out_bits_wstrb_57, // @[:@95589.4]
  output        io_out_bits_wstrb_58, // @[:@95589.4]
  output        io_out_bits_wstrb_59, // @[:@95589.4]
  output        io_out_bits_wstrb_60, // @[:@95589.4]
  output        io_out_bits_wstrb_61, // @[:@95589.4]
  output        io_out_bits_wstrb_62, // @[:@95589.4]
  output        io_out_bits_wstrb_63 // @[:@95589.4]
);
  wire [63:0] MuxN_io_ins_0_wdata_0; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_ins_0_wdata_1; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_ins_0_wdata_2; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_ins_0_wdata_3; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_ins_0_wdata_4; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_ins_0_wdata_5; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_ins_0_wdata_6; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_ins_0_wdata_7; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_0; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_1; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_2; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_3; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_4; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_5; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_6; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_7; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_8; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_9; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_10; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_11; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_12; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_13; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_14; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_15; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_16; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_17; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_18; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_19; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_20; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_21; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_22; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_23; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_24; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_25; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_26; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_27; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_28; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_29; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_30; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_31; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_32; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_33; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_34; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_35; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_36; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_37; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_38; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_39; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_40; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_41; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_42; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_43; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_44; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_45; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_46; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_47; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_48; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_49; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_50; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_51; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_52; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_53; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_54; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_55; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_56; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_57; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_58; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_59; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_60; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_61; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_62; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_0_wstrb_63; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_ins_1_wdata_0; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_ins_1_wdata_1; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_ins_1_wdata_2; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_ins_1_wdata_3; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_ins_1_wdata_4; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_ins_1_wdata_5; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_ins_1_wdata_6; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_ins_1_wdata_7; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_0; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_1; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_2; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_3; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_4; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_5; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_6; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_7; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_8; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_9; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_10; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_11; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_12; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_13; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_14; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_15; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_16; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_17; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_18; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_19; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_20; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_21; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_22; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_23; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_24; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_25; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_26; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_27; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_28; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_29; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_30; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_31; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_32; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_33; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_34; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_35; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_36; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_37; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_38; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_39; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_40; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_41; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_42; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_43; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_44; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_45; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_46; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_47; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_48; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_49; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_50; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_51; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_52; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_53; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_54; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_55; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_56; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_57; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_58; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_59; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_60; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_61; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_62; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_ins_1_wstrb_63; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_sel; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_out_wdata_0; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_out_wdata_1; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_out_wdata_2; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_out_wdata_3; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_out_wdata_4; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_out_wdata_5; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_out_wdata_6; // @[MuxN.scala 40:23:@95740.4]
  wire [63:0] MuxN_io_out_wdata_7; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_0; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_1; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_2; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_3; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_4; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_5; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_6; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_7; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_8; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_9; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_10; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_11; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_12; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_13; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_14; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_15; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_16; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_17; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_18; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_19; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_20; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_21; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_22; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_23; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_24; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_25; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_26; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_27; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_28; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_29; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_30; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_31; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_32; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_33; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_34; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_35; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_36; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_37; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_38; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_39; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_40; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_41; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_42; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_43; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_44; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_45; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_46; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_47; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_48; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_49; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_50; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_51; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_52; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_53; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_54; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_55; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_56; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_57; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_58; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_59; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_60; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_61; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_62; // @[MuxN.scala 40:23:@95740.4]
  wire  MuxN_io_out_wstrb_63; // @[MuxN.scala 40:23:@95740.4]
  wire  _T_190; // @[MuxN.scala 28:31:@95591.4]
  MuxN_1 MuxN ( // @[MuxN.scala 40:23:@95740.4]
    .io_ins_0_wdata_0(MuxN_io_ins_0_wdata_0),
    .io_ins_0_wdata_1(MuxN_io_ins_0_wdata_1),
    .io_ins_0_wdata_2(MuxN_io_ins_0_wdata_2),
    .io_ins_0_wdata_3(MuxN_io_ins_0_wdata_3),
    .io_ins_0_wdata_4(MuxN_io_ins_0_wdata_4),
    .io_ins_0_wdata_5(MuxN_io_ins_0_wdata_5),
    .io_ins_0_wdata_6(MuxN_io_ins_0_wdata_6),
    .io_ins_0_wdata_7(MuxN_io_ins_0_wdata_7),
    .io_ins_0_wstrb_0(MuxN_io_ins_0_wstrb_0),
    .io_ins_0_wstrb_1(MuxN_io_ins_0_wstrb_1),
    .io_ins_0_wstrb_2(MuxN_io_ins_0_wstrb_2),
    .io_ins_0_wstrb_3(MuxN_io_ins_0_wstrb_3),
    .io_ins_0_wstrb_4(MuxN_io_ins_0_wstrb_4),
    .io_ins_0_wstrb_5(MuxN_io_ins_0_wstrb_5),
    .io_ins_0_wstrb_6(MuxN_io_ins_0_wstrb_6),
    .io_ins_0_wstrb_7(MuxN_io_ins_0_wstrb_7),
    .io_ins_0_wstrb_8(MuxN_io_ins_0_wstrb_8),
    .io_ins_0_wstrb_9(MuxN_io_ins_0_wstrb_9),
    .io_ins_0_wstrb_10(MuxN_io_ins_0_wstrb_10),
    .io_ins_0_wstrb_11(MuxN_io_ins_0_wstrb_11),
    .io_ins_0_wstrb_12(MuxN_io_ins_0_wstrb_12),
    .io_ins_0_wstrb_13(MuxN_io_ins_0_wstrb_13),
    .io_ins_0_wstrb_14(MuxN_io_ins_0_wstrb_14),
    .io_ins_0_wstrb_15(MuxN_io_ins_0_wstrb_15),
    .io_ins_0_wstrb_16(MuxN_io_ins_0_wstrb_16),
    .io_ins_0_wstrb_17(MuxN_io_ins_0_wstrb_17),
    .io_ins_0_wstrb_18(MuxN_io_ins_0_wstrb_18),
    .io_ins_0_wstrb_19(MuxN_io_ins_0_wstrb_19),
    .io_ins_0_wstrb_20(MuxN_io_ins_0_wstrb_20),
    .io_ins_0_wstrb_21(MuxN_io_ins_0_wstrb_21),
    .io_ins_0_wstrb_22(MuxN_io_ins_0_wstrb_22),
    .io_ins_0_wstrb_23(MuxN_io_ins_0_wstrb_23),
    .io_ins_0_wstrb_24(MuxN_io_ins_0_wstrb_24),
    .io_ins_0_wstrb_25(MuxN_io_ins_0_wstrb_25),
    .io_ins_0_wstrb_26(MuxN_io_ins_0_wstrb_26),
    .io_ins_0_wstrb_27(MuxN_io_ins_0_wstrb_27),
    .io_ins_0_wstrb_28(MuxN_io_ins_0_wstrb_28),
    .io_ins_0_wstrb_29(MuxN_io_ins_0_wstrb_29),
    .io_ins_0_wstrb_30(MuxN_io_ins_0_wstrb_30),
    .io_ins_0_wstrb_31(MuxN_io_ins_0_wstrb_31),
    .io_ins_0_wstrb_32(MuxN_io_ins_0_wstrb_32),
    .io_ins_0_wstrb_33(MuxN_io_ins_0_wstrb_33),
    .io_ins_0_wstrb_34(MuxN_io_ins_0_wstrb_34),
    .io_ins_0_wstrb_35(MuxN_io_ins_0_wstrb_35),
    .io_ins_0_wstrb_36(MuxN_io_ins_0_wstrb_36),
    .io_ins_0_wstrb_37(MuxN_io_ins_0_wstrb_37),
    .io_ins_0_wstrb_38(MuxN_io_ins_0_wstrb_38),
    .io_ins_0_wstrb_39(MuxN_io_ins_0_wstrb_39),
    .io_ins_0_wstrb_40(MuxN_io_ins_0_wstrb_40),
    .io_ins_0_wstrb_41(MuxN_io_ins_0_wstrb_41),
    .io_ins_0_wstrb_42(MuxN_io_ins_0_wstrb_42),
    .io_ins_0_wstrb_43(MuxN_io_ins_0_wstrb_43),
    .io_ins_0_wstrb_44(MuxN_io_ins_0_wstrb_44),
    .io_ins_0_wstrb_45(MuxN_io_ins_0_wstrb_45),
    .io_ins_0_wstrb_46(MuxN_io_ins_0_wstrb_46),
    .io_ins_0_wstrb_47(MuxN_io_ins_0_wstrb_47),
    .io_ins_0_wstrb_48(MuxN_io_ins_0_wstrb_48),
    .io_ins_0_wstrb_49(MuxN_io_ins_0_wstrb_49),
    .io_ins_0_wstrb_50(MuxN_io_ins_0_wstrb_50),
    .io_ins_0_wstrb_51(MuxN_io_ins_0_wstrb_51),
    .io_ins_0_wstrb_52(MuxN_io_ins_0_wstrb_52),
    .io_ins_0_wstrb_53(MuxN_io_ins_0_wstrb_53),
    .io_ins_0_wstrb_54(MuxN_io_ins_0_wstrb_54),
    .io_ins_0_wstrb_55(MuxN_io_ins_0_wstrb_55),
    .io_ins_0_wstrb_56(MuxN_io_ins_0_wstrb_56),
    .io_ins_0_wstrb_57(MuxN_io_ins_0_wstrb_57),
    .io_ins_0_wstrb_58(MuxN_io_ins_0_wstrb_58),
    .io_ins_0_wstrb_59(MuxN_io_ins_0_wstrb_59),
    .io_ins_0_wstrb_60(MuxN_io_ins_0_wstrb_60),
    .io_ins_0_wstrb_61(MuxN_io_ins_0_wstrb_61),
    .io_ins_0_wstrb_62(MuxN_io_ins_0_wstrb_62),
    .io_ins_0_wstrb_63(MuxN_io_ins_0_wstrb_63),
    .io_ins_1_wdata_0(MuxN_io_ins_1_wdata_0),
    .io_ins_1_wdata_1(MuxN_io_ins_1_wdata_1),
    .io_ins_1_wdata_2(MuxN_io_ins_1_wdata_2),
    .io_ins_1_wdata_3(MuxN_io_ins_1_wdata_3),
    .io_ins_1_wdata_4(MuxN_io_ins_1_wdata_4),
    .io_ins_1_wdata_5(MuxN_io_ins_1_wdata_5),
    .io_ins_1_wdata_6(MuxN_io_ins_1_wdata_6),
    .io_ins_1_wdata_7(MuxN_io_ins_1_wdata_7),
    .io_ins_1_wstrb_0(MuxN_io_ins_1_wstrb_0),
    .io_ins_1_wstrb_1(MuxN_io_ins_1_wstrb_1),
    .io_ins_1_wstrb_2(MuxN_io_ins_1_wstrb_2),
    .io_ins_1_wstrb_3(MuxN_io_ins_1_wstrb_3),
    .io_ins_1_wstrb_4(MuxN_io_ins_1_wstrb_4),
    .io_ins_1_wstrb_5(MuxN_io_ins_1_wstrb_5),
    .io_ins_1_wstrb_6(MuxN_io_ins_1_wstrb_6),
    .io_ins_1_wstrb_7(MuxN_io_ins_1_wstrb_7),
    .io_ins_1_wstrb_8(MuxN_io_ins_1_wstrb_8),
    .io_ins_1_wstrb_9(MuxN_io_ins_1_wstrb_9),
    .io_ins_1_wstrb_10(MuxN_io_ins_1_wstrb_10),
    .io_ins_1_wstrb_11(MuxN_io_ins_1_wstrb_11),
    .io_ins_1_wstrb_12(MuxN_io_ins_1_wstrb_12),
    .io_ins_1_wstrb_13(MuxN_io_ins_1_wstrb_13),
    .io_ins_1_wstrb_14(MuxN_io_ins_1_wstrb_14),
    .io_ins_1_wstrb_15(MuxN_io_ins_1_wstrb_15),
    .io_ins_1_wstrb_16(MuxN_io_ins_1_wstrb_16),
    .io_ins_1_wstrb_17(MuxN_io_ins_1_wstrb_17),
    .io_ins_1_wstrb_18(MuxN_io_ins_1_wstrb_18),
    .io_ins_1_wstrb_19(MuxN_io_ins_1_wstrb_19),
    .io_ins_1_wstrb_20(MuxN_io_ins_1_wstrb_20),
    .io_ins_1_wstrb_21(MuxN_io_ins_1_wstrb_21),
    .io_ins_1_wstrb_22(MuxN_io_ins_1_wstrb_22),
    .io_ins_1_wstrb_23(MuxN_io_ins_1_wstrb_23),
    .io_ins_1_wstrb_24(MuxN_io_ins_1_wstrb_24),
    .io_ins_1_wstrb_25(MuxN_io_ins_1_wstrb_25),
    .io_ins_1_wstrb_26(MuxN_io_ins_1_wstrb_26),
    .io_ins_1_wstrb_27(MuxN_io_ins_1_wstrb_27),
    .io_ins_1_wstrb_28(MuxN_io_ins_1_wstrb_28),
    .io_ins_1_wstrb_29(MuxN_io_ins_1_wstrb_29),
    .io_ins_1_wstrb_30(MuxN_io_ins_1_wstrb_30),
    .io_ins_1_wstrb_31(MuxN_io_ins_1_wstrb_31),
    .io_ins_1_wstrb_32(MuxN_io_ins_1_wstrb_32),
    .io_ins_1_wstrb_33(MuxN_io_ins_1_wstrb_33),
    .io_ins_1_wstrb_34(MuxN_io_ins_1_wstrb_34),
    .io_ins_1_wstrb_35(MuxN_io_ins_1_wstrb_35),
    .io_ins_1_wstrb_36(MuxN_io_ins_1_wstrb_36),
    .io_ins_1_wstrb_37(MuxN_io_ins_1_wstrb_37),
    .io_ins_1_wstrb_38(MuxN_io_ins_1_wstrb_38),
    .io_ins_1_wstrb_39(MuxN_io_ins_1_wstrb_39),
    .io_ins_1_wstrb_40(MuxN_io_ins_1_wstrb_40),
    .io_ins_1_wstrb_41(MuxN_io_ins_1_wstrb_41),
    .io_ins_1_wstrb_42(MuxN_io_ins_1_wstrb_42),
    .io_ins_1_wstrb_43(MuxN_io_ins_1_wstrb_43),
    .io_ins_1_wstrb_44(MuxN_io_ins_1_wstrb_44),
    .io_ins_1_wstrb_45(MuxN_io_ins_1_wstrb_45),
    .io_ins_1_wstrb_46(MuxN_io_ins_1_wstrb_46),
    .io_ins_1_wstrb_47(MuxN_io_ins_1_wstrb_47),
    .io_ins_1_wstrb_48(MuxN_io_ins_1_wstrb_48),
    .io_ins_1_wstrb_49(MuxN_io_ins_1_wstrb_49),
    .io_ins_1_wstrb_50(MuxN_io_ins_1_wstrb_50),
    .io_ins_1_wstrb_51(MuxN_io_ins_1_wstrb_51),
    .io_ins_1_wstrb_52(MuxN_io_ins_1_wstrb_52),
    .io_ins_1_wstrb_53(MuxN_io_ins_1_wstrb_53),
    .io_ins_1_wstrb_54(MuxN_io_ins_1_wstrb_54),
    .io_ins_1_wstrb_55(MuxN_io_ins_1_wstrb_55),
    .io_ins_1_wstrb_56(MuxN_io_ins_1_wstrb_56),
    .io_ins_1_wstrb_57(MuxN_io_ins_1_wstrb_57),
    .io_ins_1_wstrb_58(MuxN_io_ins_1_wstrb_58),
    .io_ins_1_wstrb_59(MuxN_io_ins_1_wstrb_59),
    .io_ins_1_wstrb_60(MuxN_io_ins_1_wstrb_60),
    .io_ins_1_wstrb_61(MuxN_io_ins_1_wstrb_61),
    .io_ins_1_wstrb_62(MuxN_io_ins_1_wstrb_62),
    .io_ins_1_wstrb_63(MuxN_io_ins_1_wstrb_63),
    .io_sel(MuxN_io_sel),
    .io_out_wdata_0(MuxN_io_out_wdata_0),
    .io_out_wdata_1(MuxN_io_out_wdata_1),
    .io_out_wdata_2(MuxN_io_out_wdata_2),
    .io_out_wdata_3(MuxN_io_out_wdata_3),
    .io_out_wdata_4(MuxN_io_out_wdata_4),
    .io_out_wdata_5(MuxN_io_out_wdata_5),
    .io_out_wdata_6(MuxN_io_out_wdata_6),
    .io_out_wdata_7(MuxN_io_out_wdata_7),
    .io_out_wstrb_0(MuxN_io_out_wstrb_0),
    .io_out_wstrb_1(MuxN_io_out_wstrb_1),
    .io_out_wstrb_2(MuxN_io_out_wstrb_2),
    .io_out_wstrb_3(MuxN_io_out_wstrb_3),
    .io_out_wstrb_4(MuxN_io_out_wstrb_4),
    .io_out_wstrb_5(MuxN_io_out_wstrb_5),
    .io_out_wstrb_6(MuxN_io_out_wstrb_6),
    .io_out_wstrb_7(MuxN_io_out_wstrb_7),
    .io_out_wstrb_8(MuxN_io_out_wstrb_8),
    .io_out_wstrb_9(MuxN_io_out_wstrb_9),
    .io_out_wstrb_10(MuxN_io_out_wstrb_10),
    .io_out_wstrb_11(MuxN_io_out_wstrb_11),
    .io_out_wstrb_12(MuxN_io_out_wstrb_12),
    .io_out_wstrb_13(MuxN_io_out_wstrb_13),
    .io_out_wstrb_14(MuxN_io_out_wstrb_14),
    .io_out_wstrb_15(MuxN_io_out_wstrb_15),
    .io_out_wstrb_16(MuxN_io_out_wstrb_16),
    .io_out_wstrb_17(MuxN_io_out_wstrb_17),
    .io_out_wstrb_18(MuxN_io_out_wstrb_18),
    .io_out_wstrb_19(MuxN_io_out_wstrb_19),
    .io_out_wstrb_20(MuxN_io_out_wstrb_20),
    .io_out_wstrb_21(MuxN_io_out_wstrb_21),
    .io_out_wstrb_22(MuxN_io_out_wstrb_22),
    .io_out_wstrb_23(MuxN_io_out_wstrb_23),
    .io_out_wstrb_24(MuxN_io_out_wstrb_24),
    .io_out_wstrb_25(MuxN_io_out_wstrb_25),
    .io_out_wstrb_26(MuxN_io_out_wstrb_26),
    .io_out_wstrb_27(MuxN_io_out_wstrb_27),
    .io_out_wstrb_28(MuxN_io_out_wstrb_28),
    .io_out_wstrb_29(MuxN_io_out_wstrb_29),
    .io_out_wstrb_30(MuxN_io_out_wstrb_30),
    .io_out_wstrb_31(MuxN_io_out_wstrb_31),
    .io_out_wstrb_32(MuxN_io_out_wstrb_32),
    .io_out_wstrb_33(MuxN_io_out_wstrb_33),
    .io_out_wstrb_34(MuxN_io_out_wstrb_34),
    .io_out_wstrb_35(MuxN_io_out_wstrb_35),
    .io_out_wstrb_36(MuxN_io_out_wstrb_36),
    .io_out_wstrb_37(MuxN_io_out_wstrb_37),
    .io_out_wstrb_38(MuxN_io_out_wstrb_38),
    .io_out_wstrb_39(MuxN_io_out_wstrb_39),
    .io_out_wstrb_40(MuxN_io_out_wstrb_40),
    .io_out_wstrb_41(MuxN_io_out_wstrb_41),
    .io_out_wstrb_42(MuxN_io_out_wstrb_42),
    .io_out_wstrb_43(MuxN_io_out_wstrb_43),
    .io_out_wstrb_44(MuxN_io_out_wstrb_44),
    .io_out_wstrb_45(MuxN_io_out_wstrb_45),
    .io_out_wstrb_46(MuxN_io_out_wstrb_46),
    .io_out_wstrb_47(MuxN_io_out_wstrb_47),
    .io_out_wstrb_48(MuxN_io_out_wstrb_48),
    .io_out_wstrb_49(MuxN_io_out_wstrb_49),
    .io_out_wstrb_50(MuxN_io_out_wstrb_50),
    .io_out_wstrb_51(MuxN_io_out_wstrb_51),
    .io_out_wstrb_52(MuxN_io_out_wstrb_52),
    .io_out_wstrb_53(MuxN_io_out_wstrb_53),
    .io_out_wstrb_54(MuxN_io_out_wstrb_54),
    .io_out_wstrb_55(MuxN_io_out_wstrb_55),
    .io_out_wstrb_56(MuxN_io_out_wstrb_56),
    .io_out_wstrb_57(MuxN_io_out_wstrb_57),
    .io_out_wstrb_58(MuxN_io_out_wstrb_58),
    .io_out_wstrb_59(MuxN_io_out_wstrb_59),
    .io_out_wstrb_60(MuxN_io_out_wstrb_60),
    .io_out_wstrb_61(MuxN_io_out_wstrb_61),
    .io_out_wstrb_62(MuxN_io_out_wstrb_62),
    .io_out_wstrb_63(MuxN_io_out_wstrb_63)
  );
  assign _T_190 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@95591.4]
  assign io_in_ready = io_out_ready | _T_190; // @[MuxN.scala 71:15:@95892.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@95891.4]
  assign io_out_bits_wdata_0 = MuxN_io_out_wdata_0; // @[MuxN.scala 72:15:@95958.4]
  assign io_out_bits_wdata_1 = MuxN_io_out_wdata_1; // @[MuxN.scala 72:15:@95959.4]
  assign io_out_bits_wdata_2 = MuxN_io_out_wdata_2; // @[MuxN.scala 72:15:@95960.4]
  assign io_out_bits_wdata_3 = MuxN_io_out_wdata_3; // @[MuxN.scala 72:15:@95961.4]
  assign io_out_bits_wdata_4 = MuxN_io_out_wdata_4; // @[MuxN.scala 72:15:@95962.4]
  assign io_out_bits_wdata_5 = MuxN_io_out_wdata_5; // @[MuxN.scala 72:15:@95963.4]
  assign io_out_bits_wdata_6 = MuxN_io_out_wdata_6; // @[MuxN.scala 72:15:@95964.4]
  assign io_out_bits_wdata_7 = MuxN_io_out_wdata_7; // @[MuxN.scala 72:15:@95965.4]
  assign io_out_bits_wstrb_0 = MuxN_io_out_wstrb_0; // @[MuxN.scala 72:15:@95894.4]
  assign io_out_bits_wstrb_1 = MuxN_io_out_wstrb_1; // @[MuxN.scala 72:15:@95895.4]
  assign io_out_bits_wstrb_2 = MuxN_io_out_wstrb_2; // @[MuxN.scala 72:15:@95896.4]
  assign io_out_bits_wstrb_3 = MuxN_io_out_wstrb_3; // @[MuxN.scala 72:15:@95897.4]
  assign io_out_bits_wstrb_4 = MuxN_io_out_wstrb_4; // @[MuxN.scala 72:15:@95898.4]
  assign io_out_bits_wstrb_5 = MuxN_io_out_wstrb_5; // @[MuxN.scala 72:15:@95899.4]
  assign io_out_bits_wstrb_6 = MuxN_io_out_wstrb_6; // @[MuxN.scala 72:15:@95900.4]
  assign io_out_bits_wstrb_7 = MuxN_io_out_wstrb_7; // @[MuxN.scala 72:15:@95901.4]
  assign io_out_bits_wstrb_8 = MuxN_io_out_wstrb_8; // @[MuxN.scala 72:15:@95902.4]
  assign io_out_bits_wstrb_9 = MuxN_io_out_wstrb_9; // @[MuxN.scala 72:15:@95903.4]
  assign io_out_bits_wstrb_10 = MuxN_io_out_wstrb_10; // @[MuxN.scala 72:15:@95904.4]
  assign io_out_bits_wstrb_11 = MuxN_io_out_wstrb_11; // @[MuxN.scala 72:15:@95905.4]
  assign io_out_bits_wstrb_12 = MuxN_io_out_wstrb_12; // @[MuxN.scala 72:15:@95906.4]
  assign io_out_bits_wstrb_13 = MuxN_io_out_wstrb_13; // @[MuxN.scala 72:15:@95907.4]
  assign io_out_bits_wstrb_14 = MuxN_io_out_wstrb_14; // @[MuxN.scala 72:15:@95908.4]
  assign io_out_bits_wstrb_15 = MuxN_io_out_wstrb_15; // @[MuxN.scala 72:15:@95909.4]
  assign io_out_bits_wstrb_16 = MuxN_io_out_wstrb_16; // @[MuxN.scala 72:15:@95910.4]
  assign io_out_bits_wstrb_17 = MuxN_io_out_wstrb_17; // @[MuxN.scala 72:15:@95911.4]
  assign io_out_bits_wstrb_18 = MuxN_io_out_wstrb_18; // @[MuxN.scala 72:15:@95912.4]
  assign io_out_bits_wstrb_19 = MuxN_io_out_wstrb_19; // @[MuxN.scala 72:15:@95913.4]
  assign io_out_bits_wstrb_20 = MuxN_io_out_wstrb_20; // @[MuxN.scala 72:15:@95914.4]
  assign io_out_bits_wstrb_21 = MuxN_io_out_wstrb_21; // @[MuxN.scala 72:15:@95915.4]
  assign io_out_bits_wstrb_22 = MuxN_io_out_wstrb_22; // @[MuxN.scala 72:15:@95916.4]
  assign io_out_bits_wstrb_23 = MuxN_io_out_wstrb_23; // @[MuxN.scala 72:15:@95917.4]
  assign io_out_bits_wstrb_24 = MuxN_io_out_wstrb_24; // @[MuxN.scala 72:15:@95918.4]
  assign io_out_bits_wstrb_25 = MuxN_io_out_wstrb_25; // @[MuxN.scala 72:15:@95919.4]
  assign io_out_bits_wstrb_26 = MuxN_io_out_wstrb_26; // @[MuxN.scala 72:15:@95920.4]
  assign io_out_bits_wstrb_27 = MuxN_io_out_wstrb_27; // @[MuxN.scala 72:15:@95921.4]
  assign io_out_bits_wstrb_28 = MuxN_io_out_wstrb_28; // @[MuxN.scala 72:15:@95922.4]
  assign io_out_bits_wstrb_29 = MuxN_io_out_wstrb_29; // @[MuxN.scala 72:15:@95923.4]
  assign io_out_bits_wstrb_30 = MuxN_io_out_wstrb_30; // @[MuxN.scala 72:15:@95924.4]
  assign io_out_bits_wstrb_31 = MuxN_io_out_wstrb_31; // @[MuxN.scala 72:15:@95925.4]
  assign io_out_bits_wstrb_32 = MuxN_io_out_wstrb_32; // @[MuxN.scala 72:15:@95926.4]
  assign io_out_bits_wstrb_33 = MuxN_io_out_wstrb_33; // @[MuxN.scala 72:15:@95927.4]
  assign io_out_bits_wstrb_34 = MuxN_io_out_wstrb_34; // @[MuxN.scala 72:15:@95928.4]
  assign io_out_bits_wstrb_35 = MuxN_io_out_wstrb_35; // @[MuxN.scala 72:15:@95929.4]
  assign io_out_bits_wstrb_36 = MuxN_io_out_wstrb_36; // @[MuxN.scala 72:15:@95930.4]
  assign io_out_bits_wstrb_37 = MuxN_io_out_wstrb_37; // @[MuxN.scala 72:15:@95931.4]
  assign io_out_bits_wstrb_38 = MuxN_io_out_wstrb_38; // @[MuxN.scala 72:15:@95932.4]
  assign io_out_bits_wstrb_39 = MuxN_io_out_wstrb_39; // @[MuxN.scala 72:15:@95933.4]
  assign io_out_bits_wstrb_40 = MuxN_io_out_wstrb_40; // @[MuxN.scala 72:15:@95934.4]
  assign io_out_bits_wstrb_41 = MuxN_io_out_wstrb_41; // @[MuxN.scala 72:15:@95935.4]
  assign io_out_bits_wstrb_42 = MuxN_io_out_wstrb_42; // @[MuxN.scala 72:15:@95936.4]
  assign io_out_bits_wstrb_43 = MuxN_io_out_wstrb_43; // @[MuxN.scala 72:15:@95937.4]
  assign io_out_bits_wstrb_44 = MuxN_io_out_wstrb_44; // @[MuxN.scala 72:15:@95938.4]
  assign io_out_bits_wstrb_45 = MuxN_io_out_wstrb_45; // @[MuxN.scala 72:15:@95939.4]
  assign io_out_bits_wstrb_46 = MuxN_io_out_wstrb_46; // @[MuxN.scala 72:15:@95940.4]
  assign io_out_bits_wstrb_47 = MuxN_io_out_wstrb_47; // @[MuxN.scala 72:15:@95941.4]
  assign io_out_bits_wstrb_48 = MuxN_io_out_wstrb_48; // @[MuxN.scala 72:15:@95942.4]
  assign io_out_bits_wstrb_49 = MuxN_io_out_wstrb_49; // @[MuxN.scala 72:15:@95943.4]
  assign io_out_bits_wstrb_50 = MuxN_io_out_wstrb_50; // @[MuxN.scala 72:15:@95944.4]
  assign io_out_bits_wstrb_51 = MuxN_io_out_wstrb_51; // @[MuxN.scala 72:15:@95945.4]
  assign io_out_bits_wstrb_52 = MuxN_io_out_wstrb_52; // @[MuxN.scala 72:15:@95946.4]
  assign io_out_bits_wstrb_53 = MuxN_io_out_wstrb_53; // @[MuxN.scala 72:15:@95947.4]
  assign io_out_bits_wstrb_54 = MuxN_io_out_wstrb_54; // @[MuxN.scala 72:15:@95948.4]
  assign io_out_bits_wstrb_55 = MuxN_io_out_wstrb_55; // @[MuxN.scala 72:15:@95949.4]
  assign io_out_bits_wstrb_56 = MuxN_io_out_wstrb_56; // @[MuxN.scala 72:15:@95950.4]
  assign io_out_bits_wstrb_57 = MuxN_io_out_wstrb_57; // @[MuxN.scala 72:15:@95951.4]
  assign io_out_bits_wstrb_58 = MuxN_io_out_wstrb_58; // @[MuxN.scala 72:15:@95952.4]
  assign io_out_bits_wstrb_59 = MuxN_io_out_wstrb_59; // @[MuxN.scala 72:15:@95953.4]
  assign io_out_bits_wstrb_60 = MuxN_io_out_wstrb_60; // @[MuxN.scala 72:15:@95954.4]
  assign io_out_bits_wstrb_61 = MuxN_io_out_wstrb_61; // @[MuxN.scala 72:15:@95955.4]
  assign io_out_bits_wstrb_62 = MuxN_io_out_wstrb_62; // @[MuxN.scala 72:15:@95956.4]
  assign io_out_bits_wstrb_63 = MuxN_io_out_wstrb_63; // @[MuxN.scala 72:15:@95957.4]
  assign MuxN_io_ins_0_wdata_0 = io_in_bits_0_wdata_0; // @[MuxN.scala 41:18:@95808.4]
  assign MuxN_io_ins_0_wdata_1 = io_in_bits_0_wdata_1; // @[MuxN.scala 41:18:@95809.4]
  assign MuxN_io_ins_0_wdata_2 = io_in_bits_0_wdata_2; // @[MuxN.scala 41:18:@95810.4]
  assign MuxN_io_ins_0_wdata_3 = io_in_bits_0_wdata_3; // @[MuxN.scala 41:18:@95811.4]
  assign MuxN_io_ins_0_wdata_4 = io_in_bits_0_wdata_4; // @[MuxN.scala 41:18:@95812.4]
  assign MuxN_io_ins_0_wdata_5 = io_in_bits_0_wdata_5; // @[MuxN.scala 41:18:@95813.4]
  assign MuxN_io_ins_0_wdata_6 = io_in_bits_0_wdata_6; // @[MuxN.scala 41:18:@95814.4]
  assign MuxN_io_ins_0_wdata_7 = io_in_bits_0_wdata_7; // @[MuxN.scala 41:18:@95815.4]
  assign MuxN_io_ins_0_wstrb_0 = io_in_bits_0_wstrb_0; // @[MuxN.scala 41:18:@95744.4]
  assign MuxN_io_ins_0_wstrb_1 = io_in_bits_0_wstrb_1; // @[MuxN.scala 41:18:@95745.4]
  assign MuxN_io_ins_0_wstrb_2 = io_in_bits_0_wstrb_2; // @[MuxN.scala 41:18:@95746.4]
  assign MuxN_io_ins_0_wstrb_3 = io_in_bits_0_wstrb_3; // @[MuxN.scala 41:18:@95747.4]
  assign MuxN_io_ins_0_wstrb_4 = io_in_bits_0_wstrb_4; // @[MuxN.scala 41:18:@95748.4]
  assign MuxN_io_ins_0_wstrb_5 = io_in_bits_0_wstrb_5; // @[MuxN.scala 41:18:@95749.4]
  assign MuxN_io_ins_0_wstrb_6 = io_in_bits_0_wstrb_6; // @[MuxN.scala 41:18:@95750.4]
  assign MuxN_io_ins_0_wstrb_7 = io_in_bits_0_wstrb_7; // @[MuxN.scala 41:18:@95751.4]
  assign MuxN_io_ins_0_wstrb_8 = io_in_bits_0_wstrb_8; // @[MuxN.scala 41:18:@95752.4]
  assign MuxN_io_ins_0_wstrb_9 = io_in_bits_0_wstrb_9; // @[MuxN.scala 41:18:@95753.4]
  assign MuxN_io_ins_0_wstrb_10 = io_in_bits_0_wstrb_10; // @[MuxN.scala 41:18:@95754.4]
  assign MuxN_io_ins_0_wstrb_11 = io_in_bits_0_wstrb_11; // @[MuxN.scala 41:18:@95755.4]
  assign MuxN_io_ins_0_wstrb_12 = io_in_bits_0_wstrb_12; // @[MuxN.scala 41:18:@95756.4]
  assign MuxN_io_ins_0_wstrb_13 = io_in_bits_0_wstrb_13; // @[MuxN.scala 41:18:@95757.4]
  assign MuxN_io_ins_0_wstrb_14 = io_in_bits_0_wstrb_14; // @[MuxN.scala 41:18:@95758.4]
  assign MuxN_io_ins_0_wstrb_15 = io_in_bits_0_wstrb_15; // @[MuxN.scala 41:18:@95759.4]
  assign MuxN_io_ins_0_wstrb_16 = io_in_bits_0_wstrb_16; // @[MuxN.scala 41:18:@95760.4]
  assign MuxN_io_ins_0_wstrb_17 = io_in_bits_0_wstrb_17; // @[MuxN.scala 41:18:@95761.4]
  assign MuxN_io_ins_0_wstrb_18 = io_in_bits_0_wstrb_18; // @[MuxN.scala 41:18:@95762.4]
  assign MuxN_io_ins_0_wstrb_19 = io_in_bits_0_wstrb_19; // @[MuxN.scala 41:18:@95763.4]
  assign MuxN_io_ins_0_wstrb_20 = io_in_bits_0_wstrb_20; // @[MuxN.scala 41:18:@95764.4]
  assign MuxN_io_ins_0_wstrb_21 = io_in_bits_0_wstrb_21; // @[MuxN.scala 41:18:@95765.4]
  assign MuxN_io_ins_0_wstrb_22 = io_in_bits_0_wstrb_22; // @[MuxN.scala 41:18:@95766.4]
  assign MuxN_io_ins_0_wstrb_23 = io_in_bits_0_wstrb_23; // @[MuxN.scala 41:18:@95767.4]
  assign MuxN_io_ins_0_wstrb_24 = io_in_bits_0_wstrb_24; // @[MuxN.scala 41:18:@95768.4]
  assign MuxN_io_ins_0_wstrb_25 = io_in_bits_0_wstrb_25; // @[MuxN.scala 41:18:@95769.4]
  assign MuxN_io_ins_0_wstrb_26 = io_in_bits_0_wstrb_26; // @[MuxN.scala 41:18:@95770.4]
  assign MuxN_io_ins_0_wstrb_27 = io_in_bits_0_wstrb_27; // @[MuxN.scala 41:18:@95771.4]
  assign MuxN_io_ins_0_wstrb_28 = io_in_bits_0_wstrb_28; // @[MuxN.scala 41:18:@95772.4]
  assign MuxN_io_ins_0_wstrb_29 = io_in_bits_0_wstrb_29; // @[MuxN.scala 41:18:@95773.4]
  assign MuxN_io_ins_0_wstrb_30 = io_in_bits_0_wstrb_30; // @[MuxN.scala 41:18:@95774.4]
  assign MuxN_io_ins_0_wstrb_31 = io_in_bits_0_wstrb_31; // @[MuxN.scala 41:18:@95775.4]
  assign MuxN_io_ins_0_wstrb_32 = io_in_bits_0_wstrb_32; // @[MuxN.scala 41:18:@95776.4]
  assign MuxN_io_ins_0_wstrb_33 = io_in_bits_0_wstrb_33; // @[MuxN.scala 41:18:@95777.4]
  assign MuxN_io_ins_0_wstrb_34 = io_in_bits_0_wstrb_34; // @[MuxN.scala 41:18:@95778.4]
  assign MuxN_io_ins_0_wstrb_35 = io_in_bits_0_wstrb_35; // @[MuxN.scala 41:18:@95779.4]
  assign MuxN_io_ins_0_wstrb_36 = io_in_bits_0_wstrb_36; // @[MuxN.scala 41:18:@95780.4]
  assign MuxN_io_ins_0_wstrb_37 = io_in_bits_0_wstrb_37; // @[MuxN.scala 41:18:@95781.4]
  assign MuxN_io_ins_0_wstrb_38 = io_in_bits_0_wstrb_38; // @[MuxN.scala 41:18:@95782.4]
  assign MuxN_io_ins_0_wstrb_39 = io_in_bits_0_wstrb_39; // @[MuxN.scala 41:18:@95783.4]
  assign MuxN_io_ins_0_wstrb_40 = io_in_bits_0_wstrb_40; // @[MuxN.scala 41:18:@95784.4]
  assign MuxN_io_ins_0_wstrb_41 = io_in_bits_0_wstrb_41; // @[MuxN.scala 41:18:@95785.4]
  assign MuxN_io_ins_0_wstrb_42 = io_in_bits_0_wstrb_42; // @[MuxN.scala 41:18:@95786.4]
  assign MuxN_io_ins_0_wstrb_43 = io_in_bits_0_wstrb_43; // @[MuxN.scala 41:18:@95787.4]
  assign MuxN_io_ins_0_wstrb_44 = io_in_bits_0_wstrb_44; // @[MuxN.scala 41:18:@95788.4]
  assign MuxN_io_ins_0_wstrb_45 = io_in_bits_0_wstrb_45; // @[MuxN.scala 41:18:@95789.4]
  assign MuxN_io_ins_0_wstrb_46 = io_in_bits_0_wstrb_46; // @[MuxN.scala 41:18:@95790.4]
  assign MuxN_io_ins_0_wstrb_47 = io_in_bits_0_wstrb_47; // @[MuxN.scala 41:18:@95791.4]
  assign MuxN_io_ins_0_wstrb_48 = io_in_bits_0_wstrb_48; // @[MuxN.scala 41:18:@95792.4]
  assign MuxN_io_ins_0_wstrb_49 = io_in_bits_0_wstrb_49; // @[MuxN.scala 41:18:@95793.4]
  assign MuxN_io_ins_0_wstrb_50 = io_in_bits_0_wstrb_50; // @[MuxN.scala 41:18:@95794.4]
  assign MuxN_io_ins_0_wstrb_51 = io_in_bits_0_wstrb_51; // @[MuxN.scala 41:18:@95795.4]
  assign MuxN_io_ins_0_wstrb_52 = io_in_bits_0_wstrb_52; // @[MuxN.scala 41:18:@95796.4]
  assign MuxN_io_ins_0_wstrb_53 = io_in_bits_0_wstrb_53; // @[MuxN.scala 41:18:@95797.4]
  assign MuxN_io_ins_0_wstrb_54 = io_in_bits_0_wstrb_54; // @[MuxN.scala 41:18:@95798.4]
  assign MuxN_io_ins_0_wstrb_55 = io_in_bits_0_wstrb_55; // @[MuxN.scala 41:18:@95799.4]
  assign MuxN_io_ins_0_wstrb_56 = io_in_bits_0_wstrb_56; // @[MuxN.scala 41:18:@95800.4]
  assign MuxN_io_ins_0_wstrb_57 = io_in_bits_0_wstrb_57; // @[MuxN.scala 41:18:@95801.4]
  assign MuxN_io_ins_0_wstrb_58 = io_in_bits_0_wstrb_58; // @[MuxN.scala 41:18:@95802.4]
  assign MuxN_io_ins_0_wstrb_59 = io_in_bits_0_wstrb_59; // @[MuxN.scala 41:18:@95803.4]
  assign MuxN_io_ins_0_wstrb_60 = io_in_bits_0_wstrb_60; // @[MuxN.scala 41:18:@95804.4]
  assign MuxN_io_ins_0_wstrb_61 = io_in_bits_0_wstrb_61; // @[MuxN.scala 41:18:@95805.4]
  assign MuxN_io_ins_0_wstrb_62 = io_in_bits_0_wstrb_62; // @[MuxN.scala 41:18:@95806.4]
  assign MuxN_io_ins_0_wstrb_63 = io_in_bits_0_wstrb_63; // @[MuxN.scala 41:18:@95807.4]
  assign MuxN_io_ins_1_wdata_0 = io_in_bits_1_wdata_0; // @[MuxN.scala 41:18:@95881.4]
  assign MuxN_io_ins_1_wdata_1 = io_in_bits_1_wdata_1; // @[MuxN.scala 41:18:@95882.4]
  assign MuxN_io_ins_1_wdata_2 = io_in_bits_1_wdata_2; // @[MuxN.scala 41:18:@95883.4]
  assign MuxN_io_ins_1_wdata_3 = io_in_bits_1_wdata_3; // @[MuxN.scala 41:18:@95884.4]
  assign MuxN_io_ins_1_wdata_4 = io_in_bits_1_wdata_4; // @[MuxN.scala 41:18:@95885.4]
  assign MuxN_io_ins_1_wdata_5 = io_in_bits_1_wdata_5; // @[MuxN.scala 41:18:@95886.4]
  assign MuxN_io_ins_1_wdata_6 = io_in_bits_1_wdata_6; // @[MuxN.scala 41:18:@95887.4]
  assign MuxN_io_ins_1_wdata_7 = io_in_bits_1_wdata_7; // @[MuxN.scala 41:18:@95888.4]
  assign MuxN_io_ins_1_wstrb_0 = io_in_bits_1_wstrb_0; // @[MuxN.scala 41:18:@95817.4]
  assign MuxN_io_ins_1_wstrb_1 = io_in_bits_1_wstrb_1; // @[MuxN.scala 41:18:@95818.4]
  assign MuxN_io_ins_1_wstrb_2 = io_in_bits_1_wstrb_2; // @[MuxN.scala 41:18:@95819.4]
  assign MuxN_io_ins_1_wstrb_3 = io_in_bits_1_wstrb_3; // @[MuxN.scala 41:18:@95820.4]
  assign MuxN_io_ins_1_wstrb_4 = io_in_bits_1_wstrb_4; // @[MuxN.scala 41:18:@95821.4]
  assign MuxN_io_ins_1_wstrb_5 = io_in_bits_1_wstrb_5; // @[MuxN.scala 41:18:@95822.4]
  assign MuxN_io_ins_1_wstrb_6 = io_in_bits_1_wstrb_6; // @[MuxN.scala 41:18:@95823.4]
  assign MuxN_io_ins_1_wstrb_7 = io_in_bits_1_wstrb_7; // @[MuxN.scala 41:18:@95824.4]
  assign MuxN_io_ins_1_wstrb_8 = io_in_bits_1_wstrb_8; // @[MuxN.scala 41:18:@95825.4]
  assign MuxN_io_ins_1_wstrb_9 = io_in_bits_1_wstrb_9; // @[MuxN.scala 41:18:@95826.4]
  assign MuxN_io_ins_1_wstrb_10 = io_in_bits_1_wstrb_10; // @[MuxN.scala 41:18:@95827.4]
  assign MuxN_io_ins_1_wstrb_11 = io_in_bits_1_wstrb_11; // @[MuxN.scala 41:18:@95828.4]
  assign MuxN_io_ins_1_wstrb_12 = io_in_bits_1_wstrb_12; // @[MuxN.scala 41:18:@95829.4]
  assign MuxN_io_ins_1_wstrb_13 = io_in_bits_1_wstrb_13; // @[MuxN.scala 41:18:@95830.4]
  assign MuxN_io_ins_1_wstrb_14 = io_in_bits_1_wstrb_14; // @[MuxN.scala 41:18:@95831.4]
  assign MuxN_io_ins_1_wstrb_15 = io_in_bits_1_wstrb_15; // @[MuxN.scala 41:18:@95832.4]
  assign MuxN_io_ins_1_wstrb_16 = io_in_bits_1_wstrb_16; // @[MuxN.scala 41:18:@95833.4]
  assign MuxN_io_ins_1_wstrb_17 = io_in_bits_1_wstrb_17; // @[MuxN.scala 41:18:@95834.4]
  assign MuxN_io_ins_1_wstrb_18 = io_in_bits_1_wstrb_18; // @[MuxN.scala 41:18:@95835.4]
  assign MuxN_io_ins_1_wstrb_19 = io_in_bits_1_wstrb_19; // @[MuxN.scala 41:18:@95836.4]
  assign MuxN_io_ins_1_wstrb_20 = io_in_bits_1_wstrb_20; // @[MuxN.scala 41:18:@95837.4]
  assign MuxN_io_ins_1_wstrb_21 = io_in_bits_1_wstrb_21; // @[MuxN.scala 41:18:@95838.4]
  assign MuxN_io_ins_1_wstrb_22 = io_in_bits_1_wstrb_22; // @[MuxN.scala 41:18:@95839.4]
  assign MuxN_io_ins_1_wstrb_23 = io_in_bits_1_wstrb_23; // @[MuxN.scala 41:18:@95840.4]
  assign MuxN_io_ins_1_wstrb_24 = io_in_bits_1_wstrb_24; // @[MuxN.scala 41:18:@95841.4]
  assign MuxN_io_ins_1_wstrb_25 = io_in_bits_1_wstrb_25; // @[MuxN.scala 41:18:@95842.4]
  assign MuxN_io_ins_1_wstrb_26 = io_in_bits_1_wstrb_26; // @[MuxN.scala 41:18:@95843.4]
  assign MuxN_io_ins_1_wstrb_27 = io_in_bits_1_wstrb_27; // @[MuxN.scala 41:18:@95844.4]
  assign MuxN_io_ins_1_wstrb_28 = io_in_bits_1_wstrb_28; // @[MuxN.scala 41:18:@95845.4]
  assign MuxN_io_ins_1_wstrb_29 = io_in_bits_1_wstrb_29; // @[MuxN.scala 41:18:@95846.4]
  assign MuxN_io_ins_1_wstrb_30 = io_in_bits_1_wstrb_30; // @[MuxN.scala 41:18:@95847.4]
  assign MuxN_io_ins_1_wstrb_31 = io_in_bits_1_wstrb_31; // @[MuxN.scala 41:18:@95848.4]
  assign MuxN_io_ins_1_wstrb_32 = io_in_bits_1_wstrb_32; // @[MuxN.scala 41:18:@95849.4]
  assign MuxN_io_ins_1_wstrb_33 = io_in_bits_1_wstrb_33; // @[MuxN.scala 41:18:@95850.4]
  assign MuxN_io_ins_1_wstrb_34 = io_in_bits_1_wstrb_34; // @[MuxN.scala 41:18:@95851.4]
  assign MuxN_io_ins_1_wstrb_35 = io_in_bits_1_wstrb_35; // @[MuxN.scala 41:18:@95852.4]
  assign MuxN_io_ins_1_wstrb_36 = io_in_bits_1_wstrb_36; // @[MuxN.scala 41:18:@95853.4]
  assign MuxN_io_ins_1_wstrb_37 = io_in_bits_1_wstrb_37; // @[MuxN.scala 41:18:@95854.4]
  assign MuxN_io_ins_1_wstrb_38 = io_in_bits_1_wstrb_38; // @[MuxN.scala 41:18:@95855.4]
  assign MuxN_io_ins_1_wstrb_39 = io_in_bits_1_wstrb_39; // @[MuxN.scala 41:18:@95856.4]
  assign MuxN_io_ins_1_wstrb_40 = io_in_bits_1_wstrb_40; // @[MuxN.scala 41:18:@95857.4]
  assign MuxN_io_ins_1_wstrb_41 = io_in_bits_1_wstrb_41; // @[MuxN.scala 41:18:@95858.4]
  assign MuxN_io_ins_1_wstrb_42 = io_in_bits_1_wstrb_42; // @[MuxN.scala 41:18:@95859.4]
  assign MuxN_io_ins_1_wstrb_43 = io_in_bits_1_wstrb_43; // @[MuxN.scala 41:18:@95860.4]
  assign MuxN_io_ins_1_wstrb_44 = io_in_bits_1_wstrb_44; // @[MuxN.scala 41:18:@95861.4]
  assign MuxN_io_ins_1_wstrb_45 = io_in_bits_1_wstrb_45; // @[MuxN.scala 41:18:@95862.4]
  assign MuxN_io_ins_1_wstrb_46 = io_in_bits_1_wstrb_46; // @[MuxN.scala 41:18:@95863.4]
  assign MuxN_io_ins_1_wstrb_47 = io_in_bits_1_wstrb_47; // @[MuxN.scala 41:18:@95864.4]
  assign MuxN_io_ins_1_wstrb_48 = io_in_bits_1_wstrb_48; // @[MuxN.scala 41:18:@95865.4]
  assign MuxN_io_ins_1_wstrb_49 = io_in_bits_1_wstrb_49; // @[MuxN.scala 41:18:@95866.4]
  assign MuxN_io_ins_1_wstrb_50 = io_in_bits_1_wstrb_50; // @[MuxN.scala 41:18:@95867.4]
  assign MuxN_io_ins_1_wstrb_51 = io_in_bits_1_wstrb_51; // @[MuxN.scala 41:18:@95868.4]
  assign MuxN_io_ins_1_wstrb_52 = io_in_bits_1_wstrb_52; // @[MuxN.scala 41:18:@95869.4]
  assign MuxN_io_ins_1_wstrb_53 = io_in_bits_1_wstrb_53; // @[MuxN.scala 41:18:@95870.4]
  assign MuxN_io_ins_1_wstrb_54 = io_in_bits_1_wstrb_54; // @[MuxN.scala 41:18:@95871.4]
  assign MuxN_io_ins_1_wstrb_55 = io_in_bits_1_wstrb_55; // @[MuxN.scala 41:18:@95872.4]
  assign MuxN_io_ins_1_wstrb_56 = io_in_bits_1_wstrb_56; // @[MuxN.scala 41:18:@95873.4]
  assign MuxN_io_ins_1_wstrb_57 = io_in_bits_1_wstrb_57; // @[MuxN.scala 41:18:@95874.4]
  assign MuxN_io_ins_1_wstrb_58 = io_in_bits_1_wstrb_58; // @[MuxN.scala 41:18:@95875.4]
  assign MuxN_io_ins_1_wstrb_59 = io_in_bits_1_wstrb_59; // @[MuxN.scala 41:18:@95876.4]
  assign MuxN_io_ins_1_wstrb_60 = io_in_bits_1_wstrb_60; // @[MuxN.scala 41:18:@95877.4]
  assign MuxN_io_ins_1_wstrb_61 = io_in_bits_1_wstrb_61; // @[MuxN.scala 41:18:@95878.4]
  assign MuxN_io_ins_1_wstrb_62 = io_in_bits_1_wstrb_62; // @[MuxN.scala 41:18:@95879.4]
  assign MuxN_io_ins_1_wstrb_63 = io_in_bits_1_wstrb_63; // @[MuxN.scala 41:18:@95880.4]
  assign MuxN_io_sel = io_sel; // @[MuxN.scala 44:18:@95890.4]
endmodule
module ElementCounter( // @[:@95967.2]
  input         clock, // @[:@95968.4]
  input         reset, // @[:@95969.4]
  input         io_reset, // @[:@95970.4]
  input         io_enable, // @[:@95970.4]
  output [31:0] io_out // @[:@95970.4]
);
  reg [31:0] count; // @[Counter.scala 37:22:@95972.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_14; // @[Counter.scala 39:24:@95973.4]
  wire [31:0] newCount; // @[Counter.scala 39:24:@95974.4]
  wire [31:0] _GEN_0; // @[Counter.scala 43:26:@95979.6]
  wire [31:0] _GEN_1; // @[Counter.scala 41:18:@95975.4]
  assign _T_14 = count + 32'h1; // @[Counter.scala 39:24:@95973.4]
  assign newCount = count + 32'h1; // @[Counter.scala 39:24:@95974.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 43:26:@95979.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 41:18:@95975.4]
  assign io_out = count; // @[Counter.scala 47:10:@95982.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module StreamArbiter( // @[:@95984.2]
  input         clock, // @[:@95985.4]
  input         reset, // @[:@95986.4]
  output        io_app_0_cmd_ready, // @[:@95987.4]
  input         io_app_0_cmd_valid, // @[:@95987.4]
  input  [63:0] io_app_0_cmd_bits_addr, // @[:@95987.4]
  input  [31:0] io_app_0_cmd_bits_size, // @[:@95987.4]
  input         io_app_0_cmd_bits_isWr, // @[:@95987.4]
  input  [31:0] io_app_0_cmd_bits_tag, // @[:@95987.4]
  input         io_app_0_wdata_valid, // @[:@95987.4]
  input  [63:0] io_app_0_wdata_bits_wdata_0, // @[:@95987.4]
  input  [63:0] io_app_0_wdata_bits_wdata_1, // @[:@95987.4]
  input  [63:0] io_app_0_wdata_bits_wdata_2, // @[:@95987.4]
  input  [63:0] io_app_0_wdata_bits_wdata_3, // @[:@95987.4]
  input  [63:0] io_app_0_wdata_bits_wdata_4, // @[:@95987.4]
  input  [63:0] io_app_0_wdata_bits_wdata_5, // @[:@95987.4]
  input  [63:0] io_app_0_wdata_bits_wdata_6, // @[:@95987.4]
  input  [63:0] io_app_0_wdata_bits_wdata_7, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_0, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_1, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_2, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_3, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_4, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_5, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_6, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_7, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_8, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_9, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_10, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_11, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_12, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_13, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_14, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_15, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_16, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_17, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_18, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_19, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_20, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_21, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_22, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_23, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_24, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_25, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_26, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_27, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_28, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_29, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_30, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_31, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_32, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_33, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_34, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_35, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_36, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_37, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_38, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_39, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_40, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_41, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_42, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_43, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_44, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_45, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_46, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_47, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_48, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_49, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_50, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_51, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_52, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_53, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_54, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_55, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_56, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_57, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_58, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_59, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_60, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_61, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_62, // @[:@95987.4]
  input         io_app_0_wdata_bits_wstrb_63, // @[:@95987.4]
  input         io_app_0_rresp_ready, // @[:@95987.4]
  output        io_app_0_rresp_valid, // @[:@95987.4]
  output [63:0] io_app_0_rresp_bits_rdata_0, // @[:@95987.4]
  output [63:0] io_app_0_rresp_bits_rdata_1, // @[:@95987.4]
  output [63:0] io_app_0_rresp_bits_rdata_2, // @[:@95987.4]
  output [63:0] io_app_0_rresp_bits_rdata_3, // @[:@95987.4]
  output [63:0] io_app_0_rresp_bits_rdata_4, // @[:@95987.4]
  output [63:0] io_app_0_rresp_bits_rdata_5, // @[:@95987.4]
  output [63:0] io_app_0_rresp_bits_rdata_6, // @[:@95987.4]
  output [63:0] io_app_0_rresp_bits_rdata_7, // @[:@95987.4]
  input         io_app_0_wresp_ready, // @[:@95987.4]
  output        io_app_1_cmd_ready, // @[:@95987.4]
  input         io_app_1_cmd_valid, // @[:@95987.4]
  input  [63:0] io_app_1_cmd_bits_addr, // @[:@95987.4]
  input  [31:0] io_app_1_cmd_bits_size, // @[:@95987.4]
  input         io_app_1_cmd_bits_isWr, // @[:@95987.4]
  input  [31:0] io_app_1_cmd_bits_tag, // @[:@95987.4]
  output        io_app_1_wdata_ready, // @[:@95987.4]
  input         io_app_1_wdata_valid, // @[:@95987.4]
  input  [63:0] io_app_1_wdata_bits_wdata_0, // @[:@95987.4]
  input  [63:0] io_app_1_wdata_bits_wdata_1, // @[:@95987.4]
  input  [63:0] io_app_1_wdata_bits_wdata_2, // @[:@95987.4]
  input  [63:0] io_app_1_wdata_bits_wdata_3, // @[:@95987.4]
  input  [63:0] io_app_1_wdata_bits_wdata_4, // @[:@95987.4]
  input  [63:0] io_app_1_wdata_bits_wdata_5, // @[:@95987.4]
  input  [63:0] io_app_1_wdata_bits_wdata_6, // @[:@95987.4]
  input  [63:0] io_app_1_wdata_bits_wdata_7, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_0, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_1, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_2, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_3, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_4, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_5, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_6, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_7, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_8, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_9, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_10, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_11, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_12, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_13, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_14, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_15, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_16, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_17, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_18, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_19, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_20, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_21, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_22, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_23, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_24, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_25, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_26, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_27, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_28, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_29, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_30, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_31, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_32, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_33, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_34, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_35, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_36, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_37, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_38, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_39, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_40, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_41, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_42, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_43, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_44, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_45, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_46, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_47, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_48, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_49, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_50, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_51, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_52, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_53, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_54, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_55, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_56, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_57, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_58, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_59, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_60, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_61, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_62, // @[:@95987.4]
  input         io_app_1_wdata_bits_wstrb_63, // @[:@95987.4]
  input         io_app_1_rresp_ready, // @[:@95987.4]
  input         io_app_1_wresp_ready, // @[:@95987.4]
  output        io_app_1_wresp_valid, // @[:@95987.4]
  input         io_dram_cmd_ready, // @[:@95987.4]
  output        io_dram_cmd_valid, // @[:@95987.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@95987.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@95987.4]
  output        io_dram_cmd_bits_isWr, // @[:@95987.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@95987.4]
  input         io_dram_wdata_ready, // @[:@95987.4]
  output        io_dram_wdata_valid, // @[:@95987.4]
  output [63:0] io_dram_wdata_bits_wdata_0, // @[:@95987.4]
  output [63:0] io_dram_wdata_bits_wdata_1, // @[:@95987.4]
  output [63:0] io_dram_wdata_bits_wdata_2, // @[:@95987.4]
  output [63:0] io_dram_wdata_bits_wdata_3, // @[:@95987.4]
  output [63:0] io_dram_wdata_bits_wdata_4, // @[:@95987.4]
  output [63:0] io_dram_wdata_bits_wdata_5, // @[:@95987.4]
  output [63:0] io_dram_wdata_bits_wdata_6, // @[:@95987.4]
  output [63:0] io_dram_wdata_bits_wdata_7, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@95987.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@95987.4]
  output        io_dram_rresp_ready, // @[:@95987.4]
  input         io_dram_rresp_valid, // @[:@95987.4]
  input  [63:0] io_dram_rresp_bits_rdata_0, // @[:@95987.4]
  input  [63:0] io_dram_rresp_bits_rdata_1, // @[:@95987.4]
  input  [63:0] io_dram_rresp_bits_rdata_2, // @[:@95987.4]
  input  [63:0] io_dram_rresp_bits_rdata_3, // @[:@95987.4]
  input  [63:0] io_dram_rresp_bits_rdata_4, // @[:@95987.4]
  input  [63:0] io_dram_rresp_bits_rdata_5, // @[:@95987.4]
  input  [63:0] io_dram_rresp_bits_rdata_6, // @[:@95987.4]
  input  [63:0] io_dram_rresp_bits_rdata_7, // @[:@95987.4]
  input  [31:0] io_dram_rresp_bits_tag, // @[:@95987.4]
  output        io_dram_wresp_ready, // @[:@95987.4]
  input         io_dram_wresp_valid, // @[:@95987.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@95987.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@96282.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@96282.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@96282.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@96282.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@96282.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@96289.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@96289.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@96289.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@96289.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@96289.4]
  wire  cmdMux_io_in_ready; // @[StreamArbiter.scala 25:22:@96299.4]
  wire  cmdMux_io_in_valid; // @[StreamArbiter.scala 25:22:@96299.4]
  wire [63:0] cmdMux_io_in_bits_0_addr; // @[StreamArbiter.scala 25:22:@96299.4]
  wire [31:0] cmdMux_io_in_bits_0_size; // @[StreamArbiter.scala 25:22:@96299.4]
  wire  cmdMux_io_in_bits_0_isWr; // @[StreamArbiter.scala 25:22:@96299.4]
  wire [31:0] cmdMux_io_in_bits_0_tag; // @[StreamArbiter.scala 25:22:@96299.4]
  wire [63:0] cmdMux_io_in_bits_1_addr; // @[StreamArbiter.scala 25:22:@96299.4]
  wire [31:0] cmdMux_io_in_bits_1_size; // @[StreamArbiter.scala 25:22:@96299.4]
  wire  cmdMux_io_in_bits_1_isWr; // @[StreamArbiter.scala 25:22:@96299.4]
  wire [31:0] cmdMux_io_in_bits_1_tag; // @[StreamArbiter.scala 25:22:@96299.4]
  wire  cmdMux_io_sel; // @[StreamArbiter.scala 25:22:@96299.4]
  wire  cmdMux_io_out_ready; // @[StreamArbiter.scala 25:22:@96299.4]
  wire  cmdMux_io_out_valid; // @[StreamArbiter.scala 25:22:@96299.4]
  wire [63:0] cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 25:22:@96299.4]
  wire [31:0] cmdMux_io_out_bits_size; // @[StreamArbiter.scala 25:22:@96299.4]
  wire  cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 25:22:@96299.4]
  wire [31:0] cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 25:22:@96299.4]
  wire  wdataMux_io_in_ready; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_valid; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_in_bits_0_wdata_0; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_in_bits_0_wdata_1; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_in_bits_0_wdata_2; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_in_bits_0_wdata_3; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_in_bits_0_wdata_4; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_in_bits_0_wdata_5; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_in_bits_0_wdata_6; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_in_bits_0_wdata_7; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_0; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_1; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_2; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_3; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_4; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_5; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_6; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_7; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_8; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_9; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_10; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_11; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_12; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_13; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_14; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_15; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_16; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_17; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_18; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_19; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_20; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_21; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_22; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_23; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_24; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_25; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_26; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_27; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_28; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_29; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_30; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_31; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_32; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_33; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_34; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_35; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_36; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_37; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_38; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_39; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_40; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_41; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_42; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_43; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_44; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_45; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_46; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_47; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_48; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_49; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_50; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_51; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_52; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_53; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_54; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_55; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_56; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_57; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_58; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_59; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_60; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_61; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_62; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_0_wstrb_63; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_in_bits_1_wdata_0; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_in_bits_1_wdata_1; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_in_bits_1_wdata_2; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_in_bits_1_wdata_3; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_in_bits_1_wdata_4; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_in_bits_1_wdata_5; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_in_bits_1_wdata_6; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_in_bits_1_wdata_7; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_0; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_1; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_2; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_3; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_4; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_5; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_6; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_7; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_8; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_9; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_10; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_11; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_12; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_13; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_14; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_15; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_16; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_17; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_18; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_19; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_20; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_21; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_22; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_23; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_24; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_25; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_26; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_27; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_28; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_29; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_30; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_31; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_32; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_33; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_34; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_35; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_36; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_37; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_38; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_39; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_40; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_41; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_42; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_43; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_44; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_45; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_46; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_47; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_48; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_49; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_50; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_51; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_52; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_53; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_54; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_55; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_56; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_57; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_58; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_59; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_60; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_61; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_62; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_in_bits_1_wstrb_63; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_sel; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_ready; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_valid; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 35:24:@96341.4]
  wire [63:0] wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 35:24:@96341.4]
  wire  elementCtr_clock; // @[StreamArbiter.scala 36:26:@96344.4]
  wire  elementCtr_reset; // @[StreamArbiter.scala 36:26:@96344.4]
  wire  elementCtr_io_reset; // @[StreamArbiter.scala 36:26:@96344.4]
  wire  elementCtr_io_enable; // @[StreamArbiter.scala 36:26:@96344.4]
  wire [31:0] elementCtr_io_out; // @[StreamArbiter.scala 36:26:@96344.4]
  wire  priorityActive; // @[Mux.scala 31:69:@96277.4]
  wire  _T_408; // @[package.scala 96:25:@96287.4 package.scala 96:25:@96288.4]
  wire  _GEN_1; // @[StreamArbiter.scala 21:16:@96296.4]
  wire  _T_412; // @[package.scala 96:25:@96294.4 package.scala 96:25:@96295.4]
  wire  cmdIdx; // @[StreamArbiter.scala 21:16:@96296.4]
  wire [1:0] cmdInDecoder; // @[OneHot.scala 45:35:@96298.4]
  wire  _T_422; // @[FringeBundles.scala 114:28:@96315.4]
  wire [22:0] _T_423; // @[FringeBundles.scala 114:28:@96317.4]
  wire [23:0] _T_425; // @[FringeBundles.scala 115:37:@96320.4]
  wire  _T_433; // @[FringeBundles.scala 114:28:@96333.4]
  wire [22:0] _T_434; // @[FringeBundles.scala 114:28:@96335.4]
  wire [23:0] _T_436; // @[FringeBundles.scala 115:37:@96338.4]
  wire  _T_438; // @[StreamArbiter.scala 37:49:@96347.4]
  wire [31:0] _T_443; // @[:@96351.4 :@96352.4]
  wire [7:0] _T_444; // @[FringeBundles.scala 114:28:@96353.4]
  wire [255:0] cmdOutDecoder; // @[OneHot.scala 45:35:@96359.4]
  wire  _T_457; // @[:@96363.4]
  wire  _GEN_3; // @[StreamArbiter.scala 42:78:@96364.4]
  wire  _T_458; // @[StreamArbiter.scala 42:78:@96364.4]
  wire  _T_459; // @[StreamArbiter.scala 42:121:@96365.4]
  wire [7:0] _T_466; // @[FringeBundles.scala 132:28:@96600.4]
  wire [7:0] _T_474; // @[FringeBundles.scala 140:28:@96609.4]
  wire [255:0] rrespDecoder; // @[OneHot.scala 45:35:@96615.4]
  wire [255:0] wrespDecoder; // @[OneHot.scala 45:35:@96616.4]
  wire  _T_479; // @[StreamArbiter.scala 61:55:@96621.4]
  wire  _T_486; // @[StreamArbiter.scala 64:58:@96630.4]
  wire  _T_490; // @[StreamArbiter.scala 61:55:@96646.4]
  wire  _T_493; // @[StreamArbiter.scala 62:85:@96650.4]
  wire  _T_494; // @[StreamArbiter.scala 62:70:@96651.4]
  wire  _T_499; // @[StreamArbiter.scala 67:58:@96667.4]
  wire  _T_510; // @[:@96674.4]
  wire  _T_520; // @[:@96679.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@96282.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@96289.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  MuxPipe cmdMux ( // @[StreamArbiter.scala 25:22:@96299.4]
    .io_in_ready(cmdMux_io_in_ready),
    .io_in_valid(cmdMux_io_in_valid),
    .io_in_bits_0_addr(cmdMux_io_in_bits_0_addr),
    .io_in_bits_0_size(cmdMux_io_in_bits_0_size),
    .io_in_bits_0_isWr(cmdMux_io_in_bits_0_isWr),
    .io_in_bits_0_tag(cmdMux_io_in_bits_0_tag),
    .io_in_bits_1_addr(cmdMux_io_in_bits_1_addr),
    .io_in_bits_1_size(cmdMux_io_in_bits_1_size),
    .io_in_bits_1_isWr(cmdMux_io_in_bits_1_isWr),
    .io_in_bits_1_tag(cmdMux_io_in_bits_1_tag),
    .io_sel(cmdMux_io_sel),
    .io_out_ready(cmdMux_io_out_ready),
    .io_out_valid(cmdMux_io_out_valid),
    .io_out_bits_addr(cmdMux_io_out_bits_addr),
    .io_out_bits_size(cmdMux_io_out_bits_size),
    .io_out_bits_isWr(cmdMux_io_out_bits_isWr),
    .io_out_bits_tag(cmdMux_io_out_bits_tag)
  );
  MuxPipe_1 wdataMux ( // @[StreamArbiter.scala 35:24:@96341.4]
    .io_in_ready(wdataMux_io_in_ready),
    .io_in_valid(wdataMux_io_in_valid),
    .io_in_bits_0_wdata_0(wdataMux_io_in_bits_0_wdata_0),
    .io_in_bits_0_wdata_1(wdataMux_io_in_bits_0_wdata_1),
    .io_in_bits_0_wdata_2(wdataMux_io_in_bits_0_wdata_2),
    .io_in_bits_0_wdata_3(wdataMux_io_in_bits_0_wdata_3),
    .io_in_bits_0_wdata_4(wdataMux_io_in_bits_0_wdata_4),
    .io_in_bits_0_wdata_5(wdataMux_io_in_bits_0_wdata_5),
    .io_in_bits_0_wdata_6(wdataMux_io_in_bits_0_wdata_6),
    .io_in_bits_0_wdata_7(wdataMux_io_in_bits_0_wdata_7),
    .io_in_bits_0_wstrb_0(wdataMux_io_in_bits_0_wstrb_0),
    .io_in_bits_0_wstrb_1(wdataMux_io_in_bits_0_wstrb_1),
    .io_in_bits_0_wstrb_2(wdataMux_io_in_bits_0_wstrb_2),
    .io_in_bits_0_wstrb_3(wdataMux_io_in_bits_0_wstrb_3),
    .io_in_bits_0_wstrb_4(wdataMux_io_in_bits_0_wstrb_4),
    .io_in_bits_0_wstrb_5(wdataMux_io_in_bits_0_wstrb_5),
    .io_in_bits_0_wstrb_6(wdataMux_io_in_bits_0_wstrb_6),
    .io_in_bits_0_wstrb_7(wdataMux_io_in_bits_0_wstrb_7),
    .io_in_bits_0_wstrb_8(wdataMux_io_in_bits_0_wstrb_8),
    .io_in_bits_0_wstrb_9(wdataMux_io_in_bits_0_wstrb_9),
    .io_in_bits_0_wstrb_10(wdataMux_io_in_bits_0_wstrb_10),
    .io_in_bits_0_wstrb_11(wdataMux_io_in_bits_0_wstrb_11),
    .io_in_bits_0_wstrb_12(wdataMux_io_in_bits_0_wstrb_12),
    .io_in_bits_0_wstrb_13(wdataMux_io_in_bits_0_wstrb_13),
    .io_in_bits_0_wstrb_14(wdataMux_io_in_bits_0_wstrb_14),
    .io_in_bits_0_wstrb_15(wdataMux_io_in_bits_0_wstrb_15),
    .io_in_bits_0_wstrb_16(wdataMux_io_in_bits_0_wstrb_16),
    .io_in_bits_0_wstrb_17(wdataMux_io_in_bits_0_wstrb_17),
    .io_in_bits_0_wstrb_18(wdataMux_io_in_bits_0_wstrb_18),
    .io_in_bits_0_wstrb_19(wdataMux_io_in_bits_0_wstrb_19),
    .io_in_bits_0_wstrb_20(wdataMux_io_in_bits_0_wstrb_20),
    .io_in_bits_0_wstrb_21(wdataMux_io_in_bits_0_wstrb_21),
    .io_in_bits_0_wstrb_22(wdataMux_io_in_bits_0_wstrb_22),
    .io_in_bits_0_wstrb_23(wdataMux_io_in_bits_0_wstrb_23),
    .io_in_bits_0_wstrb_24(wdataMux_io_in_bits_0_wstrb_24),
    .io_in_bits_0_wstrb_25(wdataMux_io_in_bits_0_wstrb_25),
    .io_in_bits_0_wstrb_26(wdataMux_io_in_bits_0_wstrb_26),
    .io_in_bits_0_wstrb_27(wdataMux_io_in_bits_0_wstrb_27),
    .io_in_bits_0_wstrb_28(wdataMux_io_in_bits_0_wstrb_28),
    .io_in_bits_0_wstrb_29(wdataMux_io_in_bits_0_wstrb_29),
    .io_in_bits_0_wstrb_30(wdataMux_io_in_bits_0_wstrb_30),
    .io_in_bits_0_wstrb_31(wdataMux_io_in_bits_0_wstrb_31),
    .io_in_bits_0_wstrb_32(wdataMux_io_in_bits_0_wstrb_32),
    .io_in_bits_0_wstrb_33(wdataMux_io_in_bits_0_wstrb_33),
    .io_in_bits_0_wstrb_34(wdataMux_io_in_bits_0_wstrb_34),
    .io_in_bits_0_wstrb_35(wdataMux_io_in_bits_0_wstrb_35),
    .io_in_bits_0_wstrb_36(wdataMux_io_in_bits_0_wstrb_36),
    .io_in_bits_0_wstrb_37(wdataMux_io_in_bits_0_wstrb_37),
    .io_in_bits_0_wstrb_38(wdataMux_io_in_bits_0_wstrb_38),
    .io_in_bits_0_wstrb_39(wdataMux_io_in_bits_0_wstrb_39),
    .io_in_bits_0_wstrb_40(wdataMux_io_in_bits_0_wstrb_40),
    .io_in_bits_0_wstrb_41(wdataMux_io_in_bits_0_wstrb_41),
    .io_in_bits_0_wstrb_42(wdataMux_io_in_bits_0_wstrb_42),
    .io_in_bits_0_wstrb_43(wdataMux_io_in_bits_0_wstrb_43),
    .io_in_bits_0_wstrb_44(wdataMux_io_in_bits_0_wstrb_44),
    .io_in_bits_0_wstrb_45(wdataMux_io_in_bits_0_wstrb_45),
    .io_in_bits_0_wstrb_46(wdataMux_io_in_bits_0_wstrb_46),
    .io_in_bits_0_wstrb_47(wdataMux_io_in_bits_0_wstrb_47),
    .io_in_bits_0_wstrb_48(wdataMux_io_in_bits_0_wstrb_48),
    .io_in_bits_0_wstrb_49(wdataMux_io_in_bits_0_wstrb_49),
    .io_in_bits_0_wstrb_50(wdataMux_io_in_bits_0_wstrb_50),
    .io_in_bits_0_wstrb_51(wdataMux_io_in_bits_0_wstrb_51),
    .io_in_bits_0_wstrb_52(wdataMux_io_in_bits_0_wstrb_52),
    .io_in_bits_0_wstrb_53(wdataMux_io_in_bits_0_wstrb_53),
    .io_in_bits_0_wstrb_54(wdataMux_io_in_bits_0_wstrb_54),
    .io_in_bits_0_wstrb_55(wdataMux_io_in_bits_0_wstrb_55),
    .io_in_bits_0_wstrb_56(wdataMux_io_in_bits_0_wstrb_56),
    .io_in_bits_0_wstrb_57(wdataMux_io_in_bits_0_wstrb_57),
    .io_in_bits_0_wstrb_58(wdataMux_io_in_bits_0_wstrb_58),
    .io_in_bits_0_wstrb_59(wdataMux_io_in_bits_0_wstrb_59),
    .io_in_bits_0_wstrb_60(wdataMux_io_in_bits_0_wstrb_60),
    .io_in_bits_0_wstrb_61(wdataMux_io_in_bits_0_wstrb_61),
    .io_in_bits_0_wstrb_62(wdataMux_io_in_bits_0_wstrb_62),
    .io_in_bits_0_wstrb_63(wdataMux_io_in_bits_0_wstrb_63),
    .io_in_bits_1_wdata_0(wdataMux_io_in_bits_1_wdata_0),
    .io_in_bits_1_wdata_1(wdataMux_io_in_bits_1_wdata_1),
    .io_in_bits_1_wdata_2(wdataMux_io_in_bits_1_wdata_2),
    .io_in_bits_1_wdata_3(wdataMux_io_in_bits_1_wdata_3),
    .io_in_bits_1_wdata_4(wdataMux_io_in_bits_1_wdata_4),
    .io_in_bits_1_wdata_5(wdataMux_io_in_bits_1_wdata_5),
    .io_in_bits_1_wdata_6(wdataMux_io_in_bits_1_wdata_6),
    .io_in_bits_1_wdata_7(wdataMux_io_in_bits_1_wdata_7),
    .io_in_bits_1_wstrb_0(wdataMux_io_in_bits_1_wstrb_0),
    .io_in_bits_1_wstrb_1(wdataMux_io_in_bits_1_wstrb_1),
    .io_in_bits_1_wstrb_2(wdataMux_io_in_bits_1_wstrb_2),
    .io_in_bits_1_wstrb_3(wdataMux_io_in_bits_1_wstrb_3),
    .io_in_bits_1_wstrb_4(wdataMux_io_in_bits_1_wstrb_4),
    .io_in_bits_1_wstrb_5(wdataMux_io_in_bits_1_wstrb_5),
    .io_in_bits_1_wstrb_6(wdataMux_io_in_bits_1_wstrb_6),
    .io_in_bits_1_wstrb_7(wdataMux_io_in_bits_1_wstrb_7),
    .io_in_bits_1_wstrb_8(wdataMux_io_in_bits_1_wstrb_8),
    .io_in_bits_1_wstrb_9(wdataMux_io_in_bits_1_wstrb_9),
    .io_in_bits_1_wstrb_10(wdataMux_io_in_bits_1_wstrb_10),
    .io_in_bits_1_wstrb_11(wdataMux_io_in_bits_1_wstrb_11),
    .io_in_bits_1_wstrb_12(wdataMux_io_in_bits_1_wstrb_12),
    .io_in_bits_1_wstrb_13(wdataMux_io_in_bits_1_wstrb_13),
    .io_in_bits_1_wstrb_14(wdataMux_io_in_bits_1_wstrb_14),
    .io_in_bits_1_wstrb_15(wdataMux_io_in_bits_1_wstrb_15),
    .io_in_bits_1_wstrb_16(wdataMux_io_in_bits_1_wstrb_16),
    .io_in_bits_1_wstrb_17(wdataMux_io_in_bits_1_wstrb_17),
    .io_in_bits_1_wstrb_18(wdataMux_io_in_bits_1_wstrb_18),
    .io_in_bits_1_wstrb_19(wdataMux_io_in_bits_1_wstrb_19),
    .io_in_bits_1_wstrb_20(wdataMux_io_in_bits_1_wstrb_20),
    .io_in_bits_1_wstrb_21(wdataMux_io_in_bits_1_wstrb_21),
    .io_in_bits_1_wstrb_22(wdataMux_io_in_bits_1_wstrb_22),
    .io_in_bits_1_wstrb_23(wdataMux_io_in_bits_1_wstrb_23),
    .io_in_bits_1_wstrb_24(wdataMux_io_in_bits_1_wstrb_24),
    .io_in_bits_1_wstrb_25(wdataMux_io_in_bits_1_wstrb_25),
    .io_in_bits_1_wstrb_26(wdataMux_io_in_bits_1_wstrb_26),
    .io_in_bits_1_wstrb_27(wdataMux_io_in_bits_1_wstrb_27),
    .io_in_bits_1_wstrb_28(wdataMux_io_in_bits_1_wstrb_28),
    .io_in_bits_1_wstrb_29(wdataMux_io_in_bits_1_wstrb_29),
    .io_in_bits_1_wstrb_30(wdataMux_io_in_bits_1_wstrb_30),
    .io_in_bits_1_wstrb_31(wdataMux_io_in_bits_1_wstrb_31),
    .io_in_bits_1_wstrb_32(wdataMux_io_in_bits_1_wstrb_32),
    .io_in_bits_1_wstrb_33(wdataMux_io_in_bits_1_wstrb_33),
    .io_in_bits_1_wstrb_34(wdataMux_io_in_bits_1_wstrb_34),
    .io_in_bits_1_wstrb_35(wdataMux_io_in_bits_1_wstrb_35),
    .io_in_bits_1_wstrb_36(wdataMux_io_in_bits_1_wstrb_36),
    .io_in_bits_1_wstrb_37(wdataMux_io_in_bits_1_wstrb_37),
    .io_in_bits_1_wstrb_38(wdataMux_io_in_bits_1_wstrb_38),
    .io_in_bits_1_wstrb_39(wdataMux_io_in_bits_1_wstrb_39),
    .io_in_bits_1_wstrb_40(wdataMux_io_in_bits_1_wstrb_40),
    .io_in_bits_1_wstrb_41(wdataMux_io_in_bits_1_wstrb_41),
    .io_in_bits_1_wstrb_42(wdataMux_io_in_bits_1_wstrb_42),
    .io_in_bits_1_wstrb_43(wdataMux_io_in_bits_1_wstrb_43),
    .io_in_bits_1_wstrb_44(wdataMux_io_in_bits_1_wstrb_44),
    .io_in_bits_1_wstrb_45(wdataMux_io_in_bits_1_wstrb_45),
    .io_in_bits_1_wstrb_46(wdataMux_io_in_bits_1_wstrb_46),
    .io_in_bits_1_wstrb_47(wdataMux_io_in_bits_1_wstrb_47),
    .io_in_bits_1_wstrb_48(wdataMux_io_in_bits_1_wstrb_48),
    .io_in_bits_1_wstrb_49(wdataMux_io_in_bits_1_wstrb_49),
    .io_in_bits_1_wstrb_50(wdataMux_io_in_bits_1_wstrb_50),
    .io_in_bits_1_wstrb_51(wdataMux_io_in_bits_1_wstrb_51),
    .io_in_bits_1_wstrb_52(wdataMux_io_in_bits_1_wstrb_52),
    .io_in_bits_1_wstrb_53(wdataMux_io_in_bits_1_wstrb_53),
    .io_in_bits_1_wstrb_54(wdataMux_io_in_bits_1_wstrb_54),
    .io_in_bits_1_wstrb_55(wdataMux_io_in_bits_1_wstrb_55),
    .io_in_bits_1_wstrb_56(wdataMux_io_in_bits_1_wstrb_56),
    .io_in_bits_1_wstrb_57(wdataMux_io_in_bits_1_wstrb_57),
    .io_in_bits_1_wstrb_58(wdataMux_io_in_bits_1_wstrb_58),
    .io_in_bits_1_wstrb_59(wdataMux_io_in_bits_1_wstrb_59),
    .io_in_bits_1_wstrb_60(wdataMux_io_in_bits_1_wstrb_60),
    .io_in_bits_1_wstrb_61(wdataMux_io_in_bits_1_wstrb_61),
    .io_in_bits_1_wstrb_62(wdataMux_io_in_bits_1_wstrb_62),
    .io_in_bits_1_wstrb_63(wdataMux_io_in_bits_1_wstrb_63),
    .io_sel(wdataMux_io_sel),
    .io_out_ready(wdataMux_io_out_ready),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wstrb_0(wdataMux_io_out_bits_wstrb_0),
    .io_out_bits_wstrb_1(wdataMux_io_out_bits_wstrb_1),
    .io_out_bits_wstrb_2(wdataMux_io_out_bits_wstrb_2),
    .io_out_bits_wstrb_3(wdataMux_io_out_bits_wstrb_3),
    .io_out_bits_wstrb_4(wdataMux_io_out_bits_wstrb_4),
    .io_out_bits_wstrb_5(wdataMux_io_out_bits_wstrb_5),
    .io_out_bits_wstrb_6(wdataMux_io_out_bits_wstrb_6),
    .io_out_bits_wstrb_7(wdataMux_io_out_bits_wstrb_7),
    .io_out_bits_wstrb_8(wdataMux_io_out_bits_wstrb_8),
    .io_out_bits_wstrb_9(wdataMux_io_out_bits_wstrb_9),
    .io_out_bits_wstrb_10(wdataMux_io_out_bits_wstrb_10),
    .io_out_bits_wstrb_11(wdataMux_io_out_bits_wstrb_11),
    .io_out_bits_wstrb_12(wdataMux_io_out_bits_wstrb_12),
    .io_out_bits_wstrb_13(wdataMux_io_out_bits_wstrb_13),
    .io_out_bits_wstrb_14(wdataMux_io_out_bits_wstrb_14),
    .io_out_bits_wstrb_15(wdataMux_io_out_bits_wstrb_15),
    .io_out_bits_wstrb_16(wdataMux_io_out_bits_wstrb_16),
    .io_out_bits_wstrb_17(wdataMux_io_out_bits_wstrb_17),
    .io_out_bits_wstrb_18(wdataMux_io_out_bits_wstrb_18),
    .io_out_bits_wstrb_19(wdataMux_io_out_bits_wstrb_19),
    .io_out_bits_wstrb_20(wdataMux_io_out_bits_wstrb_20),
    .io_out_bits_wstrb_21(wdataMux_io_out_bits_wstrb_21),
    .io_out_bits_wstrb_22(wdataMux_io_out_bits_wstrb_22),
    .io_out_bits_wstrb_23(wdataMux_io_out_bits_wstrb_23),
    .io_out_bits_wstrb_24(wdataMux_io_out_bits_wstrb_24),
    .io_out_bits_wstrb_25(wdataMux_io_out_bits_wstrb_25),
    .io_out_bits_wstrb_26(wdataMux_io_out_bits_wstrb_26),
    .io_out_bits_wstrb_27(wdataMux_io_out_bits_wstrb_27),
    .io_out_bits_wstrb_28(wdataMux_io_out_bits_wstrb_28),
    .io_out_bits_wstrb_29(wdataMux_io_out_bits_wstrb_29),
    .io_out_bits_wstrb_30(wdataMux_io_out_bits_wstrb_30),
    .io_out_bits_wstrb_31(wdataMux_io_out_bits_wstrb_31),
    .io_out_bits_wstrb_32(wdataMux_io_out_bits_wstrb_32),
    .io_out_bits_wstrb_33(wdataMux_io_out_bits_wstrb_33),
    .io_out_bits_wstrb_34(wdataMux_io_out_bits_wstrb_34),
    .io_out_bits_wstrb_35(wdataMux_io_out_bits_wstrb_35),
    .io_out_bits_wstrb_36(wdataMux_io_out_bits_wstrb_36),
    .io_out_bits_wstrb_37(wdataMux_io_out_bits_wstrb_37),
    .io_out_bits_wstrb_38(wdataMux_io_out_bits_wstrb_38),
    .io_out_bits_wstrb_39(wdataMux_io_out_bits_wstrb_39),
    .io_out_bits_wstrb_40(wdataMux_io_out_bits_wstrb_40),
    .io_out_bits_wstrb_41(wdataMux_io_out_bits_wstrb_41),
    .io_out_bits_wstrb_42(wdataMux_io_out_bits_wstrb_42),
    .io_out_bits_wstrb_43(wdataMux_io_out_bits_wstrb_43),
    .io_out_bits_wstrb_44(wdataMux_io_out_bits_wstrb_44),
    .io_out_bits_wstrb_45(wdataMux_io_out_bits_wstrb_45),
    .io_out_bits_wstrb_46(wdataMux_io_out_bits_wstrb_46),
    .io_out_bits_wstrb_47(wdataMux_io_out_bits_wstrb_47),
    .io_out_bits_wstrb_48(wdataMux_io_out_bits_wstrb_48),
    .io_out_bits_wstrb_49(wdataMux_io_out_bits_wstrb_49),
    .io_out_bits_wstrb_50(wdataMux_io_out_bits_wstrb_50),
    .io_out_bits_wstrb_51(wdataMux_io_out_bits_wstrb_51),
    .io_out_bits_wstrb_52(wdataMux_io_out_bits_wstrb_52),
    .io_out_bits_wstrb_53(wdataMux_io_out_bits_wstrb_53),
    .io_out_bits_wstrb_54(wdataMux_io_out_bits_wstrb_54),
    .io_out_bits_wstrb_55(wdataMux_io_out_bits_wstrb_55),
    .io_out_bits_wstrb_56(wdataMux_io_out_bits_wstrb_56),
    .io_out_bits_wstrb_57(wdataMux_io_out_bits_wstrb_57),
    .io_out_bits_wstrb_58(wdataMux_io_out_bits_wstrb_58),
    .io_out_bits_wstrb_59(wdataMux_io_out_bits_wstrb_59),
    .io_out_bits_wstrb_60(wdataMux_io_out_bits_wstrb_60),
    .io_out_bits_wstrb_61(wdataMux_io_out_bits_wstrb_61),
    .io_out_bits_wstrb_62(wdataMux_io_out_bits_wstrb_62),
    .io_out_bits_wstrb_63(wdataMux_io_out_bits_wstrb_63)
  );
  ElementCounter elementCtr ( // @[StreamArbiter.scala 36:26:@96344.4]
    .clock(elementCtr_clock),
    .reset(elementCtr_reset),
    .io_reset(elementCtr_io_reset),
    .io_enable(elementCtr_io_enable),
    .io_out(elementCtr_io_out)
  );
  assign priorityActive = io_app_0_cmd_valid ? 1'h0 : 1'h1; // @[Mux.scala 31:69:@96277.4]
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@96287.4 package.scala 96:25:@96288.4]
  assign _GEN_1 = _T_408 ? io_app_1_cmd_valid : io_app_0_cmd_valid; // @[StreamArbiter.scala 21:16:@96296.4]
  assign _T_412 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@96294.4 package.scala 96:25:@96295.4]
  assign cmdIdx = _GEN_1 ? _T_412 : priorityActive; // @[StreamArbiter.scala 21:16:@96296.4]
  assign cmdInDecoder = 2'h1 << cmdIdx; // @[OneHot.scala 45:35:@96298.4]
  assign _T_422 = io_app_0_cmd_bits_tag[8]; // @[FringeBundles.scala 114:28:@96315.4]
  assign _T_423 = io_app_0_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@96317.4]
  assign _T_425 = {_T_423,_T_422}; // @[FringeBundles.scala 115:37:@96320.4]
  assign _T_433 = io_app_1_cmd_bits_tag[8]; // @[FringeBundles.scala 114:28:@96333.4]
  assign _T_434 = io_app_1_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@96335.4]
  assign _T_436 = {_T_434,_T_433}; // @[FringeBundles.scala 115:37:@96338.4]
  assign _T_438 = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:49:@96347.4]
  assign _T_443 = cmdMux_io_out_bits_tag; // @[:@96351.4 :@96352.4]
  assign _T_444 = _T_443[7:0]; // @[FringeBundles.scala 114:28:@96353.4]
  assign cmdOutDecoder = 256'h1 << _T_444; // @[OneHot.scala 45:35:@96359.4]
  assign _T_457 = _T_444[0]; // @[:@96363.4]
  assign _GEN_3 = _T_457 ? io_app_1_wdata_valid : io_app_0_wdata_valid; // @[StreamArbiter.scala 42:78:@96364.4]
  assign _T_458 = _GEN_3 & cmdMux_io_out_valid; // @[StreamArbiter.scala 42:78:@96364.4]
  assign _T_459 = elementCtr_io_out < cmdMux_io_out_bits_size; // @[StreamArbiter.scala 42:121:@96365.4]
  assign _T_466 = io_dram_rresp_bits_tag[7:0]; // @[FringeBundles.scala 132:28:@96600.4]
  assign _T_474 = io_dram_wresp_bits_tag[7:0]; // @[FringeBundles.scala 140:28:@96609.4]
  assign rrespDecoder = 256'h1 << _T_466; // @[OneHot.scala 45:35:@96615.4]
  assign wrespDecoder = 256'h1 << _T_474; // @[OneHot.scala 45:35:@96616.4]
  assign _T_479 = cmdInDecoder[0]; // @[StreamArbiter.scala 61:55:@96621.4]
  assign _T_486 = rrespDecoder[0]; // @[StreamArbiter.scala 64:58:@96630.4]
  assign _T_490 = cmdInDecoder[1]; // @[StreamArbiter.scala 61:55:@96646.4]
  assign _T_493 = cmdOutDecoder[1]; // @[StreamArbiter.scala 62:85:@96650.4]
  assign _T_494 = _T_438 & _T_493; // @[StreamArbiter.scala 62:70:@96651.4]
  assign _T_499 = wrespDecoder[1]; // @[StreamArbiter.scala 67:58:@96667.4]
  assign _T_510 = _T_466[0]; // @[:@96674.4]
  assign _T_520 = _T_474[0]; // @[:@96679.4]
  assign io_app_0_cmd_ready = cmdMux_io_in_ready & _T_479; // @[StreamArbiter.scala 61:19:@96623.4]
  assign io_app_0_rresp_valid = io_dram_rresp_valid & _T_486; // @[StreamArbiter.scala 64:21:@96632.4]
  assign io_app_0_rresp_bits_rdata_0 = io_dram_rresp_bits_rdata_0; // @[StreamArbiter.scala 65:20:@96634.4]
  assign io_app_0_rresp_bits_rdata_1 = io_dram_rresp_bits_rdata_1; // @[StreamArbiter.scala 65:20:@96635.4]
  assign io_app_0_rresp_bits_rdata_2 = io_dram_rresp_bits_rdata_2; // @[StreamArbiter.scala 65:20:@96636.4]
  assign io_app_0_rresp_bits_rdata_3 = io_dram_rresp_bits_rdata_3; // @[StreamArbiter.scala 65:20:@96637.4]
  assign io_app_0_rresp_bits_rdata_4 = io_dram_rresp_bits_rdata_4; // @[StreamArbiter.scala 65:20:@96638.4]
  assign io_app_0_rresp_bits_rdata_5 = io_dram_rresp_bits_rdata_5; // @[StreamArbiter.scala 65:20:@96639.4]
  assign io_app_0_rresp_bits_rdata_6 = io_dram_rresp_bits_rdata_6; // @[StreamArbiter.scala 65:20:@96640.4]
  assign io_app_0_rresp_bits_rdata_7 = io_dram_rresp_bits_rdata_7; // @[StreamArbiter.scala 65:20:@96641.4]
  assign io_app_1_cmd_ready = cmdMux_io_in_ready & _T_490; // @[StreamArbiter.scala 61:19:@96648.4]
  assign io_app_1_wdata_ready = _T_494 & _T_459; // @[StreamArbiter.scala 62:21:@96654.4]
  assign io_app_1_wresp_valid = io_dram_wresp_valid & _T_499; // @[StreamArbiter.scala 67:21:@96669.4]
  assign io_dram_cmd_valid = cmdMux_io_out_valid; // @[StreamArbiter.scala 46:15:@96520.4]
  assign io_dram_cmd_bits_addr = cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 46:15:@96519.4]
  assign io_dram_cmd_bits_size = cmdMux_io_out_bits_size; // @[StreamArbiter.scala 46:15:@96518.4]
  assign io_dram_cmd_bits_isWr = cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 46:15:@96516.4]
  assign io_dram_cmd_bits_tag = cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 46:15:@96515.4]
  assign io_dram_wdata_valid = wdataMux_io_out_valid; // @[StreamArbiter.scala 47:17:@96595.4]
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 47:17:@96587.4]
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 47:17:@96588.4]
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 47:17:@96589.4]
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 47:17:@96590.4]
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 47:17:@96591.4]
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 47:17:@96592.4]
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 47:17:@96593.4]
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 47:17:@96594.4]
  assign io_dram_wdata_bits_wstrb_0 = wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 47:17:@96523.4]
  assign io_dram_wdata_bits_wstrb_1 = wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 47:17:@96524.4]
  assign io_dram_wdata_bits_wstrb_2 = wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 47:17:@96525.4]
  assign io_dram_wdata_bits_wstrb_3 = wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 47:17:@96526.4]
  assign io_dram_wdata_bits_wstrb_4 = wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 47:17:@96527.4]
  assign io_dram_wdata_bits_wstrb_5 = wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 47:17:@96528.4]
  assign io_dram_wdata_bits_wstrb_6 = wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 47:17:@96529.4]
  assign io_dram_wdata_bits_wstrb_7 = wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 47:17:@96530.4]
  assign io_dram_wdata_bits_wstrb_8 = wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 47:17:@96531.4]
  assign io_dram_wdata_bits_wstrb_9 = wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 47:17:@96532.4]
  assign io_dram_wdata_bits_wstrb_10 = wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 47:17:@96533.4]
  assign io_dram_wdata_bits_wstrb_11 = wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 47:17:@96534.4]
  assign io_dram_wdata_bits_wstrb_12 = wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 47:17:@96535.4]
  assign io_dram_wdata_bits_wstrb_13 = wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 47:17:@96536.4]
  assign io_dram_wdata_bits_wstrb_14 = wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 47:17:@96537.4]
  assign io_dram_wdata_bits_wstrb_15 = wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 47:17:@96538.4]
  assign io_dram_wdata_bits_wstrb_16 = wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 47:17:@96539.4]
  assign io_dram_wdata_bits_wstrb_17 = wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 47:17:@96540.4]
  assign io_dram_wdata_bits_wstrb_18 = wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 47:17:@96541.4]
  assign io_dram_wdata_bits_wstrb_19 = wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 47:17:@96542.4]
  assign io_dram_wdata_bits_wstrb_20 = wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 47:17:@96543.4]
  assign io_dram_wdata_bits_wstrb_21 = wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 47:17:@96544.4]
  assign io_dram_wdata_bits_wstrb_22 = wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 47:17:@96545.4]
  assign io_dram_wdata_bits_wstrb_23 = wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 47:17:@96546.4]
  assign io_dram_wdata_bits_wstrb_24 = wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 47:17:@96547.4]
  assign io_dram_wdata_bits_wstrb_25 = wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 47:17:@96548.4]
  assign io_dram_wdata_bits_wstrb_26 = wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 47:17:@96549.4]
  assign io_dram_wdata_bits_wstrb_27 = wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 47:17:@96550.4]
  assign io_dram_wdata_bits_wstrb_28 = wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 47:17:@96551.4]
  assign io_dram_wdata_bits_wstrb_29 = wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 47:17:@96552.4]
  assign io_dram_wdata_bits_wstrb_30 = wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 47:17:@96553.4]
  assign io_dram_wdata_bits_wstrb_31 = wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 47:17:@96554.4]
  assign io_dram_wdata_bits_wstrb_32 = wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 47:17:@96555.4]
  assign io_dram_wdata_bits_wstrb_33 = wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 47:17:@96556.4]
  assign io_dram_wdata_bits_wstrb_34 = wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 47:17:@96557.4]
  assign io_dram_wdata_bits_wstrb_35 = wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 47:17:@96558.4]
  assign io_dram_wdata_bits_wstrb_36 = wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 47:17:@96559.4]
  assign io_dram_wdata_bits_wstrb_37 = wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 47:17:@96560.4]
  assign io_dram_wdata_bits_wstrb_38 = wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 47:17:@96561.4]
  assign io_dram_wdata_bits_wstrb_39 = wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 47:17:@96562.4]
  assign io_dram_wdata_bits_wstrb_40 = wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 47:17:@96563.4]
  assign io_dram_wdata_bits_wstrb_41 = wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 47:17:@96564.4]
  assign io_dram_wdata_bits_wstrb_42 = wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 47:17:@96565.4]
  assign io_dram_wdata_bits_wstrb_43 = wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 47:17:@96566.4]
  assign io_dram_wdata_bits_wstrb_44 = wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 47:17:@96567.4]
  assign io_dram_wdata_bits_wstrb_45 = wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 47:17:@96568.4]
  assign io_dram_wdata_bits_wstrb_46 = wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 47:17:@96569.4]
  assign io_dram_wdata_bits_wstrb_47 = wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 47:17:@96570.4]
  assign io_dram_wdata_bits_wstrb_48 = wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 47:17:@96571.4]
  assign io_dram_wdata_bits_wstrb_49 = wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 47:17:@96572.4]
  assign io_dram_wdata_bits_wstrb_50 = wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 47:17:@96573.4]
  assign io_dram_wdata_bits_wstrb_51 = wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 47:17:@96574.4]
  assign io_dram_wdata_bits_wstrb_52 = wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 47:17:@96575.4]
  assign io_dram_wdata_bits_wstrb_53 = wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 47:17:@96576.4]
  assign io_dram_wdata_bits_wstrb_54 = wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 47:17:@96577.4]
  assign io_dram_wdata_bits_wstrb_55 = wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 47:17:@96578.4]
  assign io_dram_wdata_bits_wstrb_56 = wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 47:17:@96579.4]
  assign io_dram_wdata_bits_wstrb_57 = wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 47:17:@96580.4]
  assign io_dram_wdata_bits_wstrb_58 = wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 47:17:@96581.4]
  assign io_dram_wdata_bits_wstrb_59 = wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 47:17:@96582.4]
  assign io_dram_wdata_bits_wstrb_60 = wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 47:17:@96583.4]
  assign io_dram_wdata_bits_wstrb_61 = wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 47:17:@96584.4]
  assign io_dram_wdata_bits_wstrb_62 = wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 47:17:@96585.4]
  assign io_dram_wdata_bits_wstrb_63 = wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 47:17:@96586.4]
  assign io_dram_rresp_ready = _T_510 ? io_app_1_rresp_ready : io_app_0_rresp_ready; // @[StreamArbiter.scala 72:23:@96675.4]
  assign io_dram_wresp_ready = _T_520 ? io_app_1_wresp_ready : io_app_0_wresp_ready; // @[StreamArbiter.scala 73:23:@96680.4]
  assign RetimeWrapper_clock = clock; // @[:@96283.4]
  assign RetimeWrapper_reset = reset; // @[:@96284.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@96286.4]
  assign RetimeWrapper_io_in = _GEN_1 ? _T_412 : priorityActive; // @[package.scala 94:16:@96285.4]
  assign RetimeWrapper_1_clock = clock; // @[:@96290.4]
  assign RetimeWrapper_1_reset = reset; // @[:@96291.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@96293.4]
  assign RetimeWrapper_1_io_in = _GEN_1 ? _T_412 : priorityActive; // @[package.scala 94:16:@96292.4]
  assign cmdMux_io_in_valid = io_app_0_cmd_valid | io_app_1_cmd_valid; // @[StreamArbiter.scala 26:22:@96303.4]
  assign cmdMux_io_in_bits_0_addr = io_app_0_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@96309.4]
  assign cmdMux_io_in_bits_0_size = io_app_0_cmd_bits_size; // @[StreamArbiter.scala 29:9:@96308.4]
  assign cmdMux_io_in_bits_0_isWr = io_app_0_cmd_bits_isWr; // @[StreamArbiter.scala 29:9:@96306.4]
  assign cmdMux_io_in_bits_0_tag = {_T_425,8'h0}; // @[StreamArbiter.scala 29:9:@96305.4 FringeBundles.scala 115:32:@96322.4]
  assign cmdMux_io_in_bits_1_addr = io_app_1_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@96327.4]
  assign cmdMux_io_in_bits_1_size = io_app_1_cmd_bits_size; // @[StreamArbiter.scala 29:9:@96326.4]
  assign cmdMux_io_in_bits_1_isWr = io_app_1_cmd_bits_isWr; // @[StreamArbiter.scala 29:9:@96324.4]
  assign cmdMux_io_in_bits_1_tag = {_T_436,8'h1}; // @[StreamArbiter.scala 29:9:@96323.4 FringeBundles.scala 115:32:@96340.4]
  assign cmdMux_io_sel = _GEN_1 ? _T_412 : priorityActive; // @[StreamArbiter.scala 27:17:@96304.4]
  assign cmdMux_io_out_ready = io_dram_cmd_valid & io_dram_cmd_ready; // @[StreamArbiter.scala 46:15:@96521.4 StreamArbiter.scala 57:23:@96619.4]
  assign wdataMux_io_in_valid = _T_458 & _T_459; // @[StreamArbiter.scala 42:24:@96367.4]
  assign wdataMux_io_in_bits_0_wdata_0 = io_app_0_wdata_bits_wdata_0; // @[StreamArbiter.scala 44:23:@96434.4]
  assign wdataMux_io_in_bits_0_wdata_1 = io_app_0_wdata_bits_wdata_1; // @[StreamArbiter.scala 44:23:@96435.4]
  assign wdataMux_io_in_bits_0_wdata_2 = io_app_0_wdata_bits_wdata_2; // @[StreamArbiter.scala 44:23:@96436.4]
  assign wdataMux_io_in_bits_0_wdata_3 = io_app_0_wdata_bits_wdata_3; // @[StreamArbiter.scala 44:23:@96437.4]
  assign wdataMux_io_in_bits_0_wdata_4 = io_app_0_wdata_bits_wdata_4; // @[StreamArbiter.scala 44:23:@96438.4]
  assign wdataMux_io_in_bits_0_wdata_5 = io_app_0_wdata_bits_wdata_5; // @[StreamArbiter.scala 44:23:@96439.4]
  assign wdataMux_io_in_bits_0_wdata_6 = io_app_0_wdata_bits_wdata_6; // @[StreamArbiter.scala 44:23:@96440.4]
  assign wdataMux_io_in_bits_0_wdata_7 = io_app_0_wdata_bits_wdata_7; // @[StreamArbiter.scala 44:23:@96441.4]
  assign wdataMux_io_in_bits_0_wstrb_0 = io_app_0_wdata_bits_wstrb_0; // @[StreamArbiter.scala 44:23:@96370.4]
  assign wdataMux_io_in_bits_0_wstrb_1 = io_app_0_wdata_bits_wstrb_1; // @[StreamArbiter.scala 44:23:@96371.4]
  assign wdataMux_io_in_bits_0_wstrb_2 = io_app_0_wdata_bits_wstrb_2; // @[StreamArbiter.scala 44:23:@96372.4]
  assign wdataMux_io_in_bits_0_wstrb_3 = io_app_0_wdata_bits_wstrb_3; // @[StreamArbiter.scala 44:23:@96373.4]
  assign wdataMux_io_in_bits_0_wstrb_4 = io_app_0_wdata_bits_wstrb_4; // @[StreamArbiter.scala 44:23:@96374.4]
  assign wdataMux_io_in_bits_0_wstrb_5 = io_app_0_wdata_bits_wstrb_5; // @[StreamArbiter.scala 44:23:@96375.4]
  assign wdataMux_io_in_bits_0_wstrb_6 = io_app_0_wdata_bits_wstrb_6; // @[StreamArbiter.scala 44:23:@96376.4]
  assign wdataMux_io_in_bits_0_wstrb_7 = io_app_0_wdata_bits_wstrb_7; // @[StreamArbiter.scala 44:23:@96377.4]
  assign wdataMux_io_in_bits_0_wstrb_8 = io_app_0_wdata_bits_wstrb_8; // @[StreamArbiter.scala 44:23:@96378.4]
  assign wdataMux_io_in_bits_0_wstrb_9 = io_app_0_wdata_bits_wstrb_9; // @[StreamArbiter.scala 44:23:@96379.4]
  assign wdataMux_io_in_bits_0_wstrb_10 = io_app_0_wdata_bits_wstrb_10; // @[StreamArbiter.scala 44:23:@96380.4]
  assign wdataMux_io_in_bits_0_wstrb_11 = io_app_0_wdata_bits_wstrb_11; // @[StreamArbiter.scala 44:23:@96381.4]
  assign wdataMux_io_in_bits_0_wstrb_12 = io_app_0_wdata_bits_wstrb_12; // @[StreamArbiter.scala 44:23:@96382.4]
  assign wdataMux_io_in_bits_0_wstrb_13 = io_app_0_wdata_bits_wstrb_13; // @[StreamArbiter.scala 44:23:@96383.4]
  assign wdataMux_io_in_bits_0_wstrb_14 = io_app_0_wdata_bits_wstrb_14; // @[StreamArbiter.scala 44:23:@96384.4]
  assign wdataMux_io_in_bits_0_wstrb_15 = io_app_0_wdata_bits_wstrb_15; // @[StreamArbiter.scala 44:23:@96385.4]
  assign wdataMux_io_in_bits_0_wstrb_16 = io_app_0_wdata_bits_wstrb_16; // @[StreamArbiter.scala 44:23:@96386.4]
  assign wdataMux_io_in_bits_0_wstrb_17 = io_app_0_wdata_bits_wstrb_17; // @[StreamArbiter.scala 44:23:@96387.4]
  assign wdataMux_io_in_bits_0_wstrb_18 = io_app_0_wdata_bits_wstrb_18; // @[StreamArbiter.scala 44:23:@96388.4]
  assign wdataMux_io_in_bits_0_wstrb_19 = io_app_0_wdata_bits_wstrb_19; // @[StreamArbiter.scala 44:23:@96389.4]
  assign wdataMux_io_in_bits_0_wstrb_20 = io_app_0_wdata_bits_wstrb_20; // @[StreamArbiter.scala 44:23:@96390.4]
  assign wdataMux_io_in_bits_0_wstrb_21 = io_app_0_wdata_bits_wstrb_21; // @[StreamArbiter.scala 44:23:@96391.4]
  assign wdataMux_io_in_bits_0_wstrb_22 = io_app_0_wdata_bits_wstrb_22; // @[StreamArbiter.scala 44:23:@96392.4]
  assign wdataMux_io_in_bits_0_wstrb_23 = io_app_0_wdata_bits_wstrb_23; // @[StreamArbiter.scala 44:23:@96393.4]
  assign wdataMux_io_in_bits_0_wstrb_24 = io_app_0_wdata_bits_wstrb_24; // @[StreamArbiter.scala 44:23:@96394.4]
  assign wdataMux_io_in_bits_0_wstrb_25 = io_app_0_wdata_bits_wstrb_25; // @[StreamArbiter.scala 44:23:@96395.4]
  assign wdataMux_io_in_bits_0_wstrb_26 = io_app_0_wdata_bits_wstrb_26; // @[StreamArbiter.scala 44:23:@96396.4]
  assign wdataMux_io_in_bits_0_wstrb_27 = io_app_0_wdata_bits_wstrb_27; // @[StreamArbiter.scala 44:23:@96397.4]
  assign wdataMux_io_in_bits_0_wstrb_28 = io_app_0_wdata_bits_wstrb_28; // @[StreamArbiter.scala 44:23:@96398.4]
  assign wdataMux_io_in_bits_0_wstrb_29 = io_app_0_wdata_bits_wstrb_29; // @[StreamArbiter.scala 44:23:@96399.4]
  assign wdataMux_io_in_bits_0_wstrb_30 = io_app_0_wdata_bits_wstrb_30; // @[StreamArbiter.scala 44:23:@96400.4]
  assign wdataMux_io_in_bits_0_wstrb_31 = io_app_0_wdata_bits_wstrb_31; // @[StreamArbiter.scala 44:23:@96401.4]
  assign wdataMux_io_in_bits_0_wstrb_32 = io_app_0_wdata_bits_wstrb_32; // @[StreamArbiter.scala 44:23:@96402.4]
  assign wdataMux_io_in_bits_0_wstrb_33 = io_app_0_wdata_bits_wstrb_33; // @[StreamArbiter.scala 44:23:@96403.4]
  assign wdataMux_io_in_bits_0_wstrb_34 = io_app_0_wdata_bits_wstrb_34; // @[StreamArbiter.scala 44:23:@96404.4]
  assign wdataMux_io_in_bits_0_wstrb_35 = io_app_0_wdata_bits_wstrb_35; // @[StreamArbiter.scala 44:23:@96405.4]
  assign wdataMux_io_in_bits_0_wstrb_36 = io_app_0_wdata_bits_wstrb_36; // @[StreamArbiter.scala 44:23:@96406.4]
  assign wdataMux_io_in_bits_0_wstrb_37 = io_app_0_wdata_bits_wstrb_37; // @[StreamArbiter.scala 44:23:@96407.4]
  assign wdataMux_io_in_bits_0_wstrb_38 = io_app_0_wdata_bits_wstrb_38; // @[StreamArbiter.scala 44:23:@96408.4]
  assign wdataMux_io_in_bits_0_wstrb_39 = io_app_0_wdata_bits_wstrb_39; // @[StreamArbiter.scala 44:23:@96409.4]
  assign wdataMux_io_in_bits_0_wstrb_40 = io_app_0_wdata_bits_wstrb_40; // @[StreamArbiter.scala 44:23:@96410.4]
  assign wdataMux_io_in_bits_0_wstrb_41 = io_app_0_wdata_bits_wstrb_41; // @[StreamArbiter.scala 44:23:@96411.4]
  assign wdataMux_io_in_bits_0_wstrb_42 = io_app_0_wdata_bits_wstrb_42; // @[StreamArbiter.scala 44:23:@96412.4]
  assign wdataMux_io_in_bits_0_wstrb_43 = io_app_0_wdata_bits_wstrb_43; // @[StreamArbiter.scala 44:23:@96413.4]
  assign wdataMux_io_in_bits_0_wstrb_44 = io_app_0_wdata_bits_wstrb_44; // @[StreamArbiter.scala 44:23:@96414.4]
  assign wdataMux_io_in_bits_0_wstrb_45 = io_app_0_wdata_bits_wstrb_45; // @[StreamArbiter.scala 44:23:@96415.4]
  assign wdataMux_io_in_bits_0_wstrb_46 = io_app_0_wdata_bits_wstrb_46; // @[StreamArbiter.scala 44:23:@96416.4]
  assign wdataMux_io_in_bits_0_wstrb_47 = io_app_0_wdata_bits_wstrb_47; // @[StreamArbiter.scala 44:23:@96417.4]
  assign wdataMux_io_in_bits_0_wstrb_48 = io_app_0_wdata_bits_wstrb_48; // @[StreamArbiter.scala 44:23:@96418.4]
  assign wdataMux_io_in_bits_0_wstrb_49 = io_app_0_wdata_bits_wstrb_49; // @[StreamArbiter.scala 44:23:@96419.4]
  assign wdataMux_io_in_bits_0_wstrb_50 = io_app_0_wdata_bits_wstrb_50; // @[StreamArbiter.scala 44:23:@96420.4]
  assign wdataMux_io_in_bits_0_wstrb_51 = io_app_0_wdata_bits_wstrb_51; // @[StreamArbiter.scala 44:23:@96421.4]
  assign wdataMux_io_in_bits_0_wstrb_52 = io_app_0_wdata_bits_wstrb_52; // @[StreamArbiter.scala 44:23:@96422.4]
  assign wdataMux_io_in_bits_0_wstrb_53 = io_app_0_wdata_bits_wstrb_53; // @[StreamArbiter.scala 44:23:@96423.4]
  assign wdataMux_io_in_bits_0_wstrb_54 = io_app_0_wdata_bits_wstrb_54; // @[StreamArbiter.scala 44:23:@96424.4]
  assign wdataMux_io_in_bits_0_wstrb_55 = io_app_0_wdata_bits_wstrb_55; // @[StreamArbiter.scala 44:23:@96425.4]
  assign wdataMux_io_in_bits_0_wstrb_56 = io_app_0_wdata_bits_wstrb_56; // @[StreamArbiter.scala 44:23:@96426.4]
  assign wdataMux_io_in_bits_0_wstrb_57 = io_app_0_wdata_bits_wstrb_57; // @[StreamArbiter.scala 44:23:@96427.4]
  assign wdataMux_io_in_bits_0_wstrb_58 = io_app_0_wdata_bits_wstrb_58; // @[StreamArbiter.scala 44:23:@96428.4]
  assign wdataMux_io_in_bits_0_wstrb_59 = io_app_0_wdata_bits_wstrb_59; // @[StreamArbiter.scala 44:23:@96429.4]
  assign wdataMux_io_in_bits_0_wstrb_60 = io_app_0_wdata_bits_wstrb_60; // @[StreamArbiter.scala 44:23:@96430.4]
  assign wdataMux_io_in_bits_0_wstrb_61 = io_app_0_wdata_bits_wstrb_61; // @[StreamArbiter.scala 44:23:@96431.4]
  assign wdataMux_io_in_bits_0_wstrb_62 = io_app_0_wdata_bits_wstrb_62; // @[StreamArbiter.scala 44:23:@96432.4]
  assign wdataMux_io_in_bits_0_wstrb_63 = io_app_0_wdata_bits_wstrb_63; // @[StreamArbiter.scala 44:23:@96433.4]
  assign wdataMux_io_in_bits_1_wdata_0 = io_app_1_wdata_bits_wdata_0; // @[StreamArbiter.scala 44:23:@96507.4]
  assign wdataMux_io_in_bits_1_wdata_1 = io_app_1_wdata_bits_wdata_1; // @[StreamArbiter.scala 44:23:@96508.4]
  assign wdataMux_io_in_bits_1_wdata_2 = io_app_1_wdata_bits_wdata_2; // @[StreamArbiter.scala 44:23:@96509.4]
  assign wdataMux_io_in_bits_1_wdata_3 = io_app_1_wdata_bits_wdata_3; // @[StreamArbiter.scala 44:23:@96510.4]
  assign wdataMux_io_in_bits_1_wdata_4 = io_app_1_wdata_bits_wdata_4; // @[StreamArbiter.scala 44:23:@96511.4]
  assign wdataMux_io_in_bits_1_wdata_5 = io_app_1_wdata_bits_wdata_5; // @[StreamArbiter.scala 44:23:@96512.4]
  assign wdataMux_io_in_bits_1_wdata_6 = io_app_1_wdata_bits_wdata_6; // @[StreamArbiter.scala 44:23:@96513.4]
  assign wdataMux_io_in_bits_1_wdata_7 = io_app_1_wdata_bits_wdata_7; // @[StreamArbiter.scala 44:23:@96514.4]
  assign wdataMux_io_in_bits_1_wstrb_0 = io_app_1_wdata_bits_wstrb_0; // @[StreamArbiter.scala 44:23:@96443.4]
  assign wdataMux_io_in_bits_1_wstrb_1 = io_app_1_wdata_bits_wstrb_1; // @[StreamArbiter.scala 44:23:@96444.4]
  assign wdataMux_io_in_bits_1_wstrb_2 = io_app_1_wdata_bits_wstrb_2; // @[StreamArbiter.scala 44:23:@96445.4]
  assign wdataMux_io_in_bits_1_wstrb_3 = io_app_1_wdata_bits_wstrb_3; // @[StreamArbiter.scala 44:23:@96446.4]
  assign wdataMux_io_in_bits_1_wstrb_4 = io_app_1_wdata_bits_wstrb_4; // @[StreamArbiter.scala 44:23:@96447.4]
  assign wdataMux_io_in_bits_1_wstrb_5 = io_app_1_wdata_bits_wstrb_5; // @[StreamArbiter.scala 44:23:@96448.4]
  assign wdataMux_io_in_bits_1_wstrb_6 = io_app_1_wdata_bits_wstrb_6; // @[StreamArbiter.scala 44:23:@96449.4]
  assign wdataMux_io_in_bits_1_wstrb_7 = io_app_1_wdata_bits_wstrb_7; // @[StreamArbiter.scala 44:23:@96450.4]
  assign wdataMux_io_in_bits_1_wstrb_8 = io_app_1_wdata_bits_wstrb_8; // @[StreamArbiter.scala 44:23:@96451.4]
  assign wdataMux_io_in_bits_1_wstrb_9 = io_app_1_wdata_bits_wstrb_9; // @[StreamArbiter.scala 44:23:@96452.4]
  assign wdataMux_io_in_bits_1_wstrb_10 = io_app_1_wdata_bits_wstrb_10; // @[StreamArbiter.scala 44:23:@96453.4]
  assign wdataMux_io_in_bits_1_wstrb_11 = io_app_1_wdata_bits_wstrb_11; // @[StreamArbiter.scala 44:23:@96454.4]
  assign wdataMux_io_in_bits_1_wstrb_12 = io_app_1_wdata_bits_wstrb_12; // @[StreamArbiter.scala 44:23:@96455.4]
  assign wdataMux_io_in_bits_1_wstrb_13 = io_app_1_wdata_bits_wstrb_13; // @[StreamArbiter.scala 44:23:@96456.4]
  assign wdataMux_io_in_bits_1_wstrb_14 = io_app_1_wdata_bits_wstrb_14; // @[StreamArbiter.scala 44:23:@96457.4]
  assign wdataMux_io_in_bits_1_wstrb_15 = io_app_1_wdata_bits_wstrb_15; // @[StreamArbiter.scala 44:23:@96458.4]
  assign wdataMux_io_in_bits_1_wstrb_16 = io_app_1_wdata_bits_wstrb_16; // @[StreamArbiter.scala 44:23:@96459.4]
  assign wdataMux_io_in_bits_1_wstrb_17 = io_app_1_wdata_bits_wstrb_17; // @[StreamArbiter.scala 44:23:@96460.4]
  assign wdataMux_io_in_bits_1_wstrb_18 = io_app_1_wdata_bits_wstrb_18; // @[StreamArbiter.scala 44:23:@96461.4]
  assign wdataMux_io_in_bits_1_wstrb_19 = io_app_1_wdata_bits_wstrb_19; // @[StreamArbiter.scala 44:23:@96462.4]
  assign wdataMux_io_in_bits_1_wstrb_20 = io_app_1_wdata_bits_wstrb_20; // @[StreamArbiter.scala 44:23:@96463.4]
  assign wdataMux_io_in_bits_1_wstrb_21 = io_app_1_wdata_bits_wstrb_21; // @[StreamArbiter.scala 44:23:@96464.4]
  assign wdataMux_io_in_bits_1_wstrb_22 = io_app_1_wdata_bits_wstrb_22; // @[StreamArbiter.scala 44:23:@96465.4]
  assign wdataMux_io_in_bits_1_wstrb_23 = io_app_1_wdata_bits_wstrb_23; // @[StreamArbiter.scala 44:23:@96466.4]
  assign wdataMux_io_in_bits_1_wstrb_24 = io_app_1_wdata_bits_wstrb_24; // @[StreamArbiter.scala 44:23:@96467.4]
  assign wdataMux_io_in_bits_1_wstrb_25 = io_app_1_wdata_bits_wstrb_25; // @[StreamArbiter.scala 44:23:@96468.4]
  assign wdataMux_io_in_bits_1_wstrb_26 = io_app_1_wdata_bits_wstrb_26; // @[StreamArbiter.scala 44:23:@96469.4]
  assign wdataMux_io_in_bits_1_wstrb_27 = io_app_1_wdata_bits_wstrb_27; // @[StreamArbiter.scala 44:23:@96470.4]
  assign wdataMux_io_in_bits_1_wstrb_28 = io_app_1_wdata_bits_wstrb_28; // @[StreamArbiter.scala 44:23:@96471.4]
  assign wdataMux_io_in_bits_1_wstrb_29 = io_app_1_wdata_bits_wstrb_29; // @[StreamArbiter.scala 44:23:@96472.4]
  assign wdataMux_io_in_bits_1_wstrb_30 = io_app_1_wdata_bits_wstrb_30; // @[StreamArbiter.scala 44:23:@96473.4]
  assign wdataMux_io_in_bits_1_wstrb_31 = io_app_1_wdata_bits_wstrb_31; // @[StreamArbiter.scala 44:23:@96474.4]
  assign wdataMux_io_in_bits_1_wstrb_32 = io_app_1_wdata_bits_wstrb_32; // @[StreamArbiter.scala 44:23:@96475.4]
  assign wdataMux_io_in_bits_1_wstrb_33 = io_app_1_wdata_bits_wstrb_33; // @[StreamArbiter.scala 44:23:@96476.4]
  assign wdataMux_io_in_bits_1_wstrb_34 = io_app_1_wdata_bits_wstrb_34; // @[StreamArbiter.scala 44:23:@96477.4]
  assign wdataMux_io_in_bits_1_wstrb_35 = io_app_1_wdata_bits_wstrb_35; // @[StreamArbiter.scala 44:23:@96478.4]
  assign wdataMux_io_in_bits_1_wstrb_36 = io_app_1_wdata_bits_wstrb_36; // @[StreamArbiter.scala 44:23:@96479.4]
  assign wdataMux_io_in_bits_1_wstrb_37 = io_app_1_wdata_bits_wstrb_37; // @[StreamArbiter.scala 44:23:@96480.4]
  assign wdataMux_io_in_bits_1_wstrb_38 = io_app_1_wdata_bits_wstrb_38; // @[StreamArbiter.scala 44:23:@96481.4]
  assign wdataMux_io_in_bits_1_wstrb_39 = io_app_1_wdata_bits_wstrb_39; // @[StreamArbiter.scala 44:23:@96482.4]
  assign wdataMux_io_in_bits_1_wstrb_40 = io_app_1_wdata_bits_wstrb_40; // @[StreamArbiter.scala 44:23:@96483.4]
  assign wdataMux_io_in_bits_1_wstrb_41 = io_app_1_wdata_bits_wstrb_41; // @[StreamArbiter.scala 44:23:@96484.4]
  assign wdataMux_io_in_bits_1_wstrb_42 = io_app_1_wdata_bits_wstrb_42; // @[StreamArbiter.scala 44:23:@96485.4]
  assign wdataMux_io_in_bits_1_wstrb_43 = io_app_1_wdata_bits_wstrb_43; // @[StreamArbiter.scala 44:23:@96486.4]
  assign wdataMux_io_in_bits_1_wstrb_44 = io_app_1_wdata_bits_wstrb_44; // @[StreamArbiter.scala 44:23:@96487.4]
  assign wdataMux_io_in_bits_1_wstrb_45 = io_app_1_wdata_bits_wstrb_45; // @[StreamArbiter.scala 44:23:@96488.4]
  assign wdataMux_io_in_bits_1_wstrb_46 = io_app_1_wdata_bits_wstrb_46; // @[StreamArbiter.scala 44:23:@96489.4]
  assign wdataMux_io_in_bits_1_wstrb_47 = io_app_1_wdata_bits_wstrb_47; // @[StreamArbiter.scala 44:23:@96490.4]
  assign wdataMux_io_in_bits_1_wstrb_48 = io_app_1_wdata_bits_wstrb_48; // @[StreamArbiter.scala 44:23:@96491.4]
  assign wdataMux_io_in_bits_1_wstrb_49 = io_app_1_wdata_bits_wstrb_49; // @[StreamArbiter.scala 44:23:@96492.4]
  assign wdataMux_io_in_bits_1_wstrb_50 = io_app_1_wdata_bits_wstrb_50; // @[StreamArbiter.scala 44:23:@96493.4]
  assign wdataMux_io_in_bits_1_wstrb_51 = io_app_1_wdata_bits_wstrb_51; // @[StreamArbiter.scala 44:23:@96494.4]
  assign wdataMux_io_in_bits_1_wstrb_52 = io_app_1_wdata_bits_wstrb_52; // @[StreamArbiter.scala 44:23:@96495.4]
  assign wdataMux_io_in_bits_1_wstrb_53 = io_app_1_wdata_bits_wstrb_53; // @[StreamArbiter.scala 44:23:@96496.4]
  assign wdataMux_io_in_bits_1_wstrb_54 = io_app_1_wdata_bits_wstrb_54; // @[StreamArbiter.scala 44:23:@96497.4]
  assign wdataMux_io_in_bits_1_wstrb_55 = io_app_1_wdata_bits_wstrb_55; // @[StreamArbiter.scala 44:23:@96498.4]
  assign wdataMux_io_in_bits_1_wstrb_56 = io_app_1_wdata_bits_wstrb_56; // @[StreamArbiter.scala 44:23:@96499.4]
  assign wdataMux_io_in_bits_1_wstrb_57 = io_app_1_wdata_bits_wstrb_57; // @[StreamArbiter.scala 44:23:@96500.4]
  assign wdataMux_io_in_bits_1_wstrb_58 = io_app_1_wdata_bits_wstrb_58; // @[StreamArbiter.scala 44:23:@96501.4]
  assign wdataMux_io_in_bits_1_wstrb_59 = io_app_1_wdata_bits_wstrb_59; // @[StreamArbiter.scala 44:23:@96502.4]
  assign wdataMux_io_in_bits_1_wstrb_60 = io_app_1_wdata_bits_wstrb_60; // @[StreamArbiter.scala 44:23:@96503.4]
  assign wdataMux_io_in_bits_1_wstrb_61 = io_app_1_wdata_bits_wstrb_61; // @[StreamArbiter.scala 44:23:@96504.4]
  assign wdataMux_io_in_bits_1_wstrb_62 = io_app_1_wdata_bits_wstrb_62; // @[StreamArbiter.scala 44:23:@96505.4]
  assign wdataMux_io_in_bits_1_wstrb_63 = io_app_1_wdata_bits_wstrb_63; // @[StreamArbiter.scala 44:23:@96506.4]
  assign wdataMux_io_sel = _T_444[0]; // @[StreamArbiter.scala 43:19:@96368.4]
  assign wdataMux_io_out_ready = io_dram_wdata_valid & io_dram_wdata_ready; // @[StreamArbiter.scala 47:17:@96596.4 StreamArbiter.scala 58:25:@96620.4]
  assign elementCtr_clock = clock; // @[:@96345.4]
  assign elementCtr_reset = reset; // @[:@96346.4]
  assign elementCtr_io_reset = cmdMux_io_out_ready; // @[StreamArbiter.scala 38:23:@96349.4]
  assign elementCtr_io_enable = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:24:@96348.4]
endmodule
module Counter_112( // @[:@96682.2]
  input         clock, // @[:@96683.4]
  input         reset, // @[:@96684.4]
  input         io_reset, // @[:@96685.4]
  input         io_enable, // @[:@96685.4]
  input  [31:0] io_stride, // @[:@96685.4]
  output [31:0] io_out, // @[:@96685.4]
  output [31:0] io_next // @[:@96685.4]
);
  reg [31:0] count; // @[Counter.scala 15:22:@96687.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_17; // @[Counter.scala 17:24:@96688.4]
  wire [31:0] newCount; // @[Counter.scala 17:24:@96689.4]
  wire [31:0] _GEN_0; // @[Counter.scala 21:26:@96694.6]
  wire [31:0] _GEN_1; // @[Counter.scala 19:18:@96690.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@96688.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@96689.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@96694.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 19:18:@96690.4]
  assign io_out = count; // @[Counter.scala 25:10:@96697.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@96698.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module AXICmdSplit( // @[:@96700.2]
  input         clock, // @[:@96701.4]
  input         reset, // @[:@96702.4]
  output        io_in_cmd_ready, // @[:@96703.4]
  input         io_in_cmd_valid, // @[:@96703.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@96703.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@96703.4]
  input         io_in_cmd_bits_isWr, // @[:@96703.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@96703.4]
  output        io_in_wdata_ready, // @[:@96703.4]
  input         io_in_wdata_valid, // @[:@96703.4]
  input  [63:0] io_in_wdata_bits_wdata_0, // @[:@96703.4]
  input  [63:0] io_in_wdata_bits_wdata_1, // @[:@96703.4]
  input  [63:0] io_in_wdata_bits_wdata_2, // @[:@96703.4]
  input  [63:0] io_in_wdata_bits_wdata_3, // @[:@96703.4]
  input  [63:0] io_in_wdata_bits_wdata_4, // @[:@96703.4]
  input  [63:0] io_in_wdata_bits_wdata_5, // @[:@96703.4]
  input  [63:0] io_in_wdata_bits_wdata_6, // @[:@96703.4]
  input  [63:0] io_in_wdata_bits_wdata_7, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@96703.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@96703.4]
  input         io_in_rresp_ready, // @[:@96703.4]
  output        io_in_rresp_valid, // @[:@96703.4]
  output [63:0] io_in_rresp_bits_rdata_0, // @[:@96703.4]
  output [63:0] io_in_rresp_bits_rdata_1, // @[:@96703.4]
  output [63:0] io_in_rresp_bits_rdata_2, // @[:@96703.4]
  output [63:0] io_in_rresp_bits_rdata_3, // @[:@96703.4]
  output [63:0] io_in_rresp_bits_rdata_4, // @[:@96703.4]
  output [63:0] io_in_rresp_bits_rdata_5, // @[:@96703.4]
  output [63:0] io_in_rresp_bits_rdata_6, // @[:@96703.4]
  output [63:0] io_in_rresp_bits_rdata_7, // @[:@96703.4]
  output [31:0] io_in_rresp_bits_tag, // @[:@96703.4]
  input         io_in_wresp_ready, // @[:@96703.4]
  output        io_in_wresp_valid, // @[:@96703.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@96703.4]
  input         io_out_cmd_ready, // @[:@96703.4]
  output        io_out_cmd_valid, // @[:@96703.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@96703.4]
  output [31:0] io_out_cmd_bits_size, // @[:@96703.4]
  output        io_out_cmd_bits_isWr, // @[:@96703.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@96703.4]
  input         io_out_wdata_ready, // @[:@96703.4]
  output        io_out_wdata_valid, // @[:@96703.4]
  output [63:0] io_out_wdata_bits_wdata_0, // @[:@96703.4]
  output [63:0] io_out_wdata_bits_wdata_1, // @[:@96703.4]
  output [63:0] io_out_wdata_bits_wdata_2, // @[:@96703.4]
  output [63:0] io_out_wdata_bits_wdata_3, // @[:@96703.4]
  output [63:0] io_out_wdata_bits_wdata_4, // @[:@96703.4]
  output [63:0] io_out_wdata_bits_wdata_5, // @[:@96703.4]
  output [63:0] io_out_wdata_bits_wdata_6, // @[:@96703.4]
  output [63:0] io_out_wdata_bits_wdata_7, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@96703.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@96703.4]
  output        io_out_rresp_ready, // @[:@96703.4]
  input         io_out_rresp_valid, // @[:@96703.4]
  input  [63:0] io_out_rresp_bits_rdata_0, // @[:@96703.4]
  input  [63:0] io_out_rresp_bits_rdata_1, // @[:@96703.4]
  input  [63:0] io_out_rresp_bits_rdata_2, // @[:@96703.4]
  input  [63:0] io_out_rresp_bits_rdata_3, // @[:@96703.4]
  input  [63:0] io_out_rresp_bits_rdata_4, // @[:@96703.4]
  input  [63:0] io_out_rresp_bits_rdata_5, // @[:@96703.4]
  input  [63:0] io_out_rresp_bits_rdata_6, // @[:@96703.4]
  input  [63:0] io_out_rresp_bits_rdata_7, // @[:@96703.4]
  input  [31:0] io_out_rresp_bits_tag, // @[:@96703.4]
  output        io_out_wresp_ready, // @[:@96703.4]
  input         io_out_wresp_valid, // @[:@96703.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@96703.4]
);
  wire  cmdSizeCounter_clock; // @[AXIProtocol.scala 18:30:@96801.4]
  wire  cmdSizeCounter_reset; // @[AXIProtocol.scala 18:30:@96801.4]
  wire  cmdSizeCounter_io_reset; // @[AXIProtocol.scala 18:30:@96801.4]
  wire  cmdSizeCounter_io_enable; // @[AXIProtocol.scala 18:30:@96801.4]
  wire [31:0] cmdSizeCounter_io_stride; // @[AXIProtocol.scala 18:30:@96801.4]
  wire [31:0] cmdSizeCounter_io_out; // @[AXIProtocol.scala 18:30:@96801.4]
  wire [31:0] cmdSizeCounter_io_next; // @[AXIProtocol.scala 18:30:@96801.4]
  wire [32:0] _T_199; // @[AXIProtocol.scala 20:46:@96804.4]
  wire [32:0] _T_200; // @[AXIProtocol.scala 20:46:@96805.4]
  wire [31:0] cmdSizeRemaining; // @[AXIProtocol.scala 20:46:@96806.4]
  wire  lastCmd; // @[AXIProtocol.scala 23:35:@96807.4]
  wire [37:0] _GEN_0; // @[AXIProtocol.scala 27:47:@96810.4]
  wire [37:0] addrOffsetBytes; // @[AXIProtocol.scala 27:47:@96810.4]
  wire [63:0] _GEN_1; // @[AXIProtocol.scala 28:49:@96811.4]
  wire [64:0] _T_201; // @[AXIProtocol.scala 28:49:@96811.4]
  wire [63:0] cmdAddr_bits; // @[AXIProtocol.scala 28:49:@96812.4]
  wire [57:0] _T_204; // @[FringeBundles.scala 158:22:@96815.4]
  wire [7:0] cmdTag_streamID; // @[FringeBundles.scala 114:28:@96822.4]
  wire [22:0] cmdTag_uid; // @[FringeBundles.scala 114:28:@96826.4]
  wire [23:0] _T_214; // @[FringeBundles.scala 115:37:@96829.4]
  wire  cmdIssue; // @[AXIProtocol.scala 36:35:@96832.4]
  wire  _T_223; // @[FringeBundles.scala 140:28:@96843.4]
  Counter_112 cmdSizeCounter ( // @[AXIProtocol.scala 18:30:@96801.4]
    .clock(cmdSizeCounter_clock),
    .reset(cmdSizeCounter_reset),
    .io_reset(cmdSizeCounter_io_reset),
    .io_enable(cmdSizeCounter_io_enable),
    .io_stride(cmdSizeCounter_io_stride),
    .io_out(cmdSizeCounter_io_out),
    .io_next(cmdSizeCounter_io_next)
  );
  assign _T_199 = io_in_cmd_bits_size - cmdSizeCounter_io_out; // @[AXIProtocol.scala 20:46:@96804.4]
  assign _T_200 = $unsigned(_T_199); // @[AXIProtocol.scala 20:46:@96805.4]
  assign cmdSizeRemaining = _T_200[31:0]; // @[AXIProtocol.scala 20:46:@96806.4]
  assign lastCmd = cmdSizeRemaining <= 32'h100; // @[AXIProtocol.scala 23:35:@96807.4]
  assign _GEN_0 = {{6'd0}, cmdSizeCounter_io_out}; // @[AXIProtocol.scala 27:47:@96810.4]
  assign addrOffsetBytes = _GEN_0 << 6; // @[AXIProtocol.scala 27:47:@96810.4]
  assign _GEN_1 = {{26'd0}, addrOffsetBytes}; // @[AXIProtocol.scala 28:49:@96811.4]
  assign _T_201 = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@96811.4]
  assign cmdAddr_bits = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@96812.4]
  assign _T_204 = cmdAddr_bits[63:6]; // @[FringeBundles.scala 158:22:@96815.4]
  assign cmdTag_streamID = io_in_cmd_bits_tag[7:0]; // @[FringeBundles.scala 114:28:@96822.4]
  assign cmdTag_uid = io_in_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@96826.4]
  assign _T_214 = {cmdTag_uid,lastCmd}; // @[FringeBundles.scala 115:37:@96829.4]
  assign cmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 36:35:@96832.4]
  assign _T_223 = io_out_wresp_bits_tag[8]; // @[FringeBundles.scala 140:28:@96843.4]
  assign io_in_cmd_ready = lastCmd & cmdIssue; // @[AXIProtocol.scala 15:10:@96800.4 AXIProtocol.scala 38:19:@96834.4]
  assign io_in_wdata_ready = io_out_wdata_ready; // @[AXIProtocol.scala 15:10:@96793.4]
  assign io_in_rresp_valid = io_out_rresp_valid; // @[AXIProtocol.scala 15:10:@96717.4]
  assign io_in_rresp_bits_rdata_0 = io_out_rresp_bits_rdata_0; // @[AXIProtocol.scala 15:10:@96709.4]
  assign io_in_rresp_bits_rdata_1 = io_out_rresp_bits_rdata_1; // @[AXIProtocol.scala 15:10:@96710.4]
  assign io_in_rresp_bits_rdata_2 = io_out_rresp_bits_rdata_2; // @[AXIProtocol.scala 15:10:@96711.4]
  assign io_in_rresp_bits_rdata_3 = io_out_rresp_bits_rdata_3; // @[AXIProtocol.scala 15:10:@96712.4]
  assign io_in_rresp_bits_rdata_4 = io_out_rresp_bits_rdata_4; // @[AXIProtocol.scala 15:10:@96713.4]
  assign io_in_rresp_bits_rdata_5 = io_out_rresp_bits_rdata_5; // @[AXIProtocol.scala 15:10:@96714.4]
  assign io_in_rresp_bits_rdata_6 = io_out_rresp_bits_rdata_6; // @[AXIProtocol.scala 15:10:@96715.4]
  assign io_in_rresp_bits_rdata_7 = io_out_rresp_bits_rdata_7; // @[AXIProtocol.scala 15:10:@96716.4]
  assign io_in_rresp_bits_tag = io_out_rresp_bits_tag; // @[AXIProtocol.scala 15:10:@96708.4]
  assign io_in_wresp_valid = io_out_wresp_valid & _T_223; // @[AXIProtocol.scala 15:10:@96706.4 AXIProtocol.scala 46:21:@96848.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 15:10:@96705.4]
  assign io_out_cmd_valid = io_in_cmd_valid; // @[AXIProtocol.scala 15:10:@96799.4]
  assign io_out_cmd_bits_addr = {_T_204,6'h0}; // @[AXIProtocol.scala 15:10:@96798.4 AXIProtocol.scala 29:24:@96817.4]
  assign io_out_cmd_bits_size = lastCmd ? cmdSizeRemaining : 32'h100; // @[AXIProtocol.scala 15:10:@96797.4 AXIProtocol.scala 25:24:@96809.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 15:10:@96795.4]
  assign io_out_cmd_bits_tag = {_T_214,cmdTag_streamID}; // @[AXIProtocol.scala 15:10:@96794.4 FringeBundles.scala 115:32:@96831.4]
  assign io_out_wdata_valid = io_in_wdata_valid; // @[AXIProtocol.scala 15:10:@96792.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 15:10:@96784.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 15:10:@96785.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 15:10:@96786.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 15:10:@96787.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 15:10:@96788.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 15:10:@96789.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 15:10:@96790.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 15:10:@96791.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 15:10:@96720.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 15:10:@96721.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 15:10:@96722.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 15:10:@96723.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 15:10:@96724.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 15:10:@96725.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 15:10:@96726.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 15:10:@96727.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 15:10:@96728.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 15:10:@96729.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 15:10:@96730.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 15:10:@96731.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 15:10:@96732.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 15:10:@96733.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 15:10:@96734.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 15:10:@96735.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 15:10:@96736.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 15:10:@96737.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 15:10:@96738.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 15:10:@96739.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 15:10:@96740.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 15:10:@96741.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 15:10:@96742.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 15:10:@96743.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 15:10:@96744.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 15:10:@96745.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 15:10:@96746.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 15:10:@96747.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 15:10:@96748.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 15:10:@96749.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 15:10:@96750.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 15:10:@96751.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 15:10:@96752.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 15:10:@96753.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 15:10:@96754.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 15:10:@96755.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 15:10:@96756.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 15:10:@96757.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 15:10:@96758.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 15:10:@96759.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 15:10:@96760.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 15:10:@96761.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 15:10:@96762.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 15:10:@96763.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 15:10:@96764.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 15:10:@96765.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 15:10:@96766.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 15:10:@96767.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 15:10:@96768.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 15:10:@96769.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 15:10:@96770.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 15:10:@96771.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 15:10:@96772.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 15:10:@96773.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 15:10:@96774.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 15:10:@96775.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 15:10:@96776.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 15:10:@96777.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 15:10:@96778.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 15:10:@96779.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 15:10:@96780.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 15:10:@96781.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 15:10:@96782.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 15:10:@96783.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 15:10:@96718.4]
  assign io_out_wresp_ready = _T_223 ? io_in_wresp_ready : 1'h1; // @[AXIProtocol.scala 15:10:@96707.4 AXIProtocol.scala 47:22:@96850.4]
  assign cmdSizeCounter_clock = clock; // @[:@96802.4]
  assign cmdSizeCounter_reset = reset; // @[:@96803.4]
  assign cmdSizeCounter_io_reset = lastCmd & cmdIssue; // @[AXIProtocol.scala 40:27:@96835.4]
  assign cmdSizeCounter_io_enable = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 41:28:@96836.4]
  assign cmdSizeCounter_io_stride = 32'h100; // @[AXIProtocol.scala 42:28:@96837.4]
endmodule
module AXICmdIssue( // @[:@96870.2]
  input         clock, // @[:@96871.4]
  input         reset, // @[:@96872.4]
  output        io_in_cmd_ready, // @[:@96873.4]
  input         io_in_cmd_valid, // @[:@96873.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@96873.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@96873.4]
  input         io_in_cmd_bits_isWr, // @[:@96873.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@96873.4]
  output        io_in_wdata_ready, // @[:@96873.4]
  input         io_in_wdata_valid, // @[:@96873.4]
  input  [63:0] io_in_wdata_bits_wdata_0, // @[:@96873.4]
  input  [63:0] io_in_wdata_bits_wdata_1, // @[:@96873.4]
  input  [63:0] io_in_wdata_bits_wdata_2, // @[:@96873.4]
  input  [63:0] io_in_wdata_bits_wdata_3, // @[:@96873.4]
  input  [63:0] io_in_wdata_bits_wdata_4, // @[:@96873.4]
  input  [63:0] io_in_wdata_bits_wdata_5, // @[:@96873.4]
  input  [63:0] io_in_wdata_bits_wdata_6, // @[:@96873.4]
  input  [63:0] io_in_wdata_bits_wdata_7, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@96873.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@96873.4]
  input         io_in_rresp_ready, // @[:@96873.4]
  output        io_in_rresp_valid, // @[:@96873.4]
  output [63:0] io_in_rresp_bits_rdata_0, // @[:@96873.4]
  output [63:0] io_in_rresp_bits_rdata_1, // @[:@96873.4]
  output [63:0] io_in_rresp_bits_rdata_2, // @[:@96873.4]
  output [63:0] io_in_rresp_bits_rdata_3, // @[:@96873.4]
  output [63:0] io_in_rresp_bits_rdata_4, // @[:@96873.4]
  output [63:0] io_in_rresp_bits_rdata_5, // @[:@96873.4]
  output [63:0] io_in_rresp_bits_rdata_6, // @[:@96873.4]
  output [63:0] io_in_rresp_bits_rdata_7, // @[:@96873.4]
  output [31:0] io_in_rresp_bits_tag, // @[:@96873.4]
  input         io_in_wresp_ready, // @[:@96873.4]
  output        io_in_wresp_valid, // @[:@96873.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@96873.4]
  input         io_out_cmd_ready, // @[:@96873.4]
  output        io_out_cmd_valid, // @[:@96873.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@96873.4]
  output [31:0] io_out_cmd_bits_size, // @[:@96873.4]
  output        io_out_cmd_bits_isWr, // @[:@96873.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@96873.4]
  input         io_out_wdata_ready, // @[:@96873.4]
  output        io_out_wdata_valid, // @[:@96873.4]
  output [63:0] io_out_wdata_bits_wdata_0, // @[:@96873.4]
  output [63:0] io_out_wdata_bits_wdata_1, // @[:@96873.4]
  output [63:0] io_out_wdata_bits_wdata_2, // @[:@96873.4]
  output [63:0] io_out_wdata_bits_wdata_3, // @[:@96873.4]
  output [63:0] io_out_wdata_bits_wdata_4, // @[:@96873.4]
  output [63:0] io_out_wdata_bits_wdata_5, // @[:@96873.4]
  output [63:0] io_out_wdata_bits_wdata_6, // @[:@96873.4]
  output [63:0] io_out_wdata_bits_wdata_7, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@96873.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@96873.4]
  output        io_out_wdata_bits_wlast, // @[:@96873.4]
  output        io_out_rresp_ready, // @[:@96873.4]
  input         io_out_rresp_valid, // @[:@96873.4]
  input  [63:0] io_out_rresp_bits_rdata_0, // @[:@96873.4]
  input  [63:0] io_out_rresp_bits_rdata_1, // @[:@96873.4]
  input  [63:0] io_out_rresp_bits_rdata_2, // @[:@96873.4]
  input  [63:0] io_out_rresp_bits_rdata_3, // @[:@96873.4]
  input  [63:0] io_out_rresp_bits_rdata_4, // @[:@96873.4]
  input  [63:0] io_out_rresp_bits_rdata_5, // @[:@96873.4]
  input  [63:0] io_out_rresp_bits_rdata_6, // @[:@96873.4]
  input  [63:0] io_out_rresp_bits_rdata_7, // @[:@96873.4]
  input  [31:0] io_out_rresp_bits_tag, // @[:@96873.4]
  output        io_out_wresp_ready, // @[:@96873.4]
  input         io_out_wresp_valid, // @[:@96873.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@96873.4]
);
  wire  wdataCounter_clock; // @[AXIProtocol.scala 59:28:@96971.4]
  wire  wdataCounter_reset; // @[AXIProtocol.scala 59:28:@96971.4]
  wire  wdataCounter_io_reset; // @[AXIProtocol.scala 59:28:@96971.4]
  wire  wdataCounter_io_enable; // @[AXIProtocol.scala 59:28:@96971.4]
  wire [31:0] wdataCounter_io_stride; // @[AXIProtocol.scala 59:28:@96971.4]
  wire [31:0] wdataCounter_io_out; // @[AXIProtocol.scala 59:28:@96971.4]
  wire [31:0] wdataCounter_io_next; // @[AXIProtocol.scala 59:28:@96971.4]
  reg  writeIssued; // @[AXIProtocol.scala 61:28:@96974.4]
  reg [31:0] _RAND_0;
  wire  dramCmdIssue; // @[AXIProtocol.scala 63:39:@96975.4]
  wire  dramWriteIssue; // @[AXIProtocol.scala 64:43:@96976.4]
  wire  _T_201; // @[AXIProtocol.scala 68:54:@96977.4]
  wire  wlast; // @[AXIProtocol.scala 68:30:@96978.4]
  wire  _T_203; // @[AXIProtocol.scala 72:28:@96984.6]
  wire  _GEN_0; // @[AXIProtocol.scala 72:40:@96985.6]
  wire  _GEN_1; // @[AXIProtocol.scala 70:15:@96980.4]
  wire  _T_208; // @[AXIProtocol.scala 84:55:@96994.4]
  wire  _T_210; // @[AXIProtocol.scala 84:44:@96995.4]
  Counter_112 wdataCounter ( // @[AXIProtocol.scala 59:28:@96971.4]
    .clock(wdataCounter_clock),
    .reset(wdataCounter_reset),
    .io_reset(wdataCounter_io_reset),
    .io_enable(wdataCounter_io_enable),
    .io_stride(wdataCounter_io_stride),
    .io_out(wdataCounter_io_out),
    .io_next(wdataCounter_io_next)
  );
  assign dramCmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 63:39:@96975.4]
  assign dramWriteIssue = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 64:43:@96976.4]
  assign _T_201 = wdataCounter_io_next == io_in_cmd_bits_size; // @[AXIProtocol.scala 68:54:@96977.4]
  assign wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 68:30:@96978.4]
  assign _T_203 = dramCmdIssue & io_in_cmd_bits_isWr; // @[AXIProtocol.scala 72:28:@96984.6]
  assign _GEN_0 = _T_203 ? 1'h1 : writeIssued; // @[AXIProtocol.scala 72:40:@96985.6]
  assign _GEN_1 = wlast ? 1'h0 : _GEN_0; // @[AXIProtocol.scala 70:15:@96980.4]
  assign _T_208 = writeIssued == 1'h0; // @[AXIProtocol.scala 84:55:@96994.4]
  assign _T_210 = io_in_cmd_bits_isWr ? _T_208 : 1'h1; // @[AXIProtocol.scala 84:44:@96995.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? wlast : dramCmdIssue; // @[AXIProtocol.scala 56:10:@96970.4 AXIProtocol.scala 81:19:@96992.4]
  assign io_in_wdata_ready = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 56:10:@96963.4 AXIProtocol.scala 82:21:@96993.4]
  assign io_in_rresp_valid = io_out_rresp_valid; // @[AXIProtocol.scala 56:10:@96887.4]
  assign io_in_rresp_bits_rdata_0 = io_out_rresp_bits_rdata_0; // @[AXIProtocol.scala 56:10:@96879.4]
  assign io_in_rresp_bits_rdata_1 = io_out_rresp_bits_rdata_1; // @[AXIProtocol.scala 56:10:@96880.4]
  assign io_in_rresp_bits_rdata_2 = io_out_rresp_bits_rdata_2; // @[AXIProtocol.scala 56:10:@96881.4]
  assign io_in_rresp_bits_rdata_3 = io_out_rresp_bits_rdata_3; // @[AXIProtocol.scala 56:10:@96882.4]
  assign io_in_rresp_bits_rdata_4 = io_out_rresp_bits_rdata_4; // @[AXIProtocol.scala 56:10:@96883.4]
  assign io_in_rresp_bits_rdata_5 = io_out_rresp_bits_rdata_5; // @[AXIProtocol.scala 56:10:@96884.4]
  assign io_in_rresp_bits_rdata_6 = io_out_rresp_bits_rdata_6; // @[AXIProtocol.scala 56:10:@96885.4]
  assign io_in_rresp_bits_rdata_7 = io_out_rresp_bits_rdata_7; // @[AXIProtocol.scala 56:10:@96886.4]
  assign io_in_rresp_bits_tag = io_out_rresp_bits_tag; // @[AXIProtocol.scala 56:10:@96878.4]
  assign io_in_wresp_valid = io_out_wresp_valid; // @[AXIProtocol.scala 56:10:@96876.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 56:10:@96875.4]
  assign io_out_cmd_valid = io_in_cmd_valid & _T_210; // @[AXIProtocol.scala 56:10:@96969.4 AXIProtocol.scala 84:20:@96997.4]
  assign io_out_cmd_bits_addr = io_in_cmd_bits_addr; // @[AXIProtocol.scala 56:10:@96968.4]
  assign io_out_cmd_bits_size = io_in_cmd_bits_size; // @[AXIProtocol.scala 56:10:@96967.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 56:10:@96965.4]
  assign io_out_cmd_bits_tag = io_in_cmd_bits_tag; // @[AXIProtocol.scala 56:10:@96964.4]
  assign io_out_wdata_valid = io_in_wdata_valid & writeIssued; // @[AXIProtocol.scala 56:10:@96962.4 AXIProtocol.scala 86:22:@96999.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 56:10:@96954.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 56:10:@96955.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 56:10:@96956.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 56:10:@96957.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 56:10:@96958.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 56:10:@96959.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 56:10:@96960.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 56:10:@96961.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 56:10:@96890.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 56:10:@96891.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 56:10:@96892.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 56:10:@96893.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 56:10:@96894.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 56:10:@96895.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 56:10:@96896.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 56:10:@96897.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 56:10:@96898.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 56:10:@96899.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 56:10:@96900.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 56:10:@96901.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 56:10:@96902.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 56:10:@96903.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 56:10:@96904.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 56:10:@96905.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 56:10:@96906.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 56:10:@96907.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 56:10:@96908.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 56:10:@96909.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 56:10:@96910.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 56:10:@96911.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 56:10:@96912.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 56:10:@96913.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 56:10:@96914.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 56:10:@96915.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 56:10:@96916.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 56:10:@96917.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 56:10:@96918.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 56:10:@96919.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 56:10:@96920.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 56:10:@96921.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 56:10:@96922.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 56:10:@96923.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 56:10:@96924.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 56:10:@96925.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 56:10:@96926.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 56:10:@96927.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 56:10:@96928.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 56:10:@96929.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 56:10:@96930.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 56:10:@96931.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 56:10:@96932.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 56:10:@96933.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 56:10:@96934.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 56:10:@96935.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 56:10:@96936.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 56:10:@96937.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 56:10:@96938.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 56:10:@96939.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 56:10:@96940.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 56:10:@96941.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 56:10:@96942.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 56:10:@96943.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 56:10:@96944.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 56:10:@96945.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 56:10:@96946.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 56:10:@96947.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 56:10:@96948.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 56:10:@96949.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 56:10:@96950.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 56:10:@96951.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 56:10:@96952.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 56:10:@96953.4]
  assign io_out_wdata_bits_wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 56:10:@96889.4 AXIProtocol.scala 87:27:@97000.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 56:10:@96888.4]
  assign io_out_wresp_ready = io_in_wresp_ready; // @[AXIProtocol.scala 56:10:@96877.4]
  assign wdataCounter_clock = clock; // @[:@96972.4]
  assign wdataCounter_reset = reset; // @[:@96973.4]
  assign wdataCounter_io_reset = dramWriteIssue & _T_201; // @[AXIProtocol.scala 76:25:@96988.4]
  assign wdataCounter_io_enable = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 77:26:@96989.4]
  assign wdataCounter_io_stride = 32'h1; // @[AXIProtocol.scala 78:26:@96990.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeIssued = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      writeIssued <= 1'h0;
    end else begin
      if (wlast) begin
        writeIssued <= 1'h0;
      end else begin
        if (_T_203) begin
          writeIssued <= 1'h1;
        end
      end
    end
  end
endmodule
module DRAMArbiter( // @[:@97002.2]
  input         clock, // @[:@97003.4]
  input         reset, // @[:@97004.4]
  input         io_enable, // @[:@97005.4]
  output        io_app_loads_0_cmd_ready, // @[:@97005.4]
  input         io_app_loads_0_cmd_valid, // @[:@97005.4]
  input  [63:0] io_app_loads_0_cmd_bits_addr, // @[:@97005.4]
  input  [31:0] io_app_loads_0_cmd_bits_size, // @[:@97005.4]
  input         io_app_loads_0_data_ready, // @[:@97005.4]
  output        io_app_loads_0_data_valid, // @[:@97005.4]
  output [31:0] io_app_loads_0_data_bits_rdata_0, // @[:@97005.4]
  output        io_app_stores_0_cmd_ready, // @[:@97005.4]
  input         io_app_stores_0_cmd_valid, // @[:@97005.4]
  input  [63:0] io_app_stores_0_cmd_bits_addr, // @[:@97005.4]
  input  [31:0] io_app_stores_0_cmd_bits_size, // @[:@97005.4]
  output        io_app_stores_0_data_ready, // @[:@97005.4]
  input         io_app_stores_0_data_valid, // @[:@97005.4]
  input  [31:0] io_app_stores_0_data_bits_wdata_0, // @[:@97005.4]
  input         io_app_stores_0_data_bits_wstrb, // @[:@97005.4]
  input         io_app_stores_0_wresp_ready, // @[:@97005.4]
  output        io_app_stores_0_wresp_valid, // @[:@97005.4]
  output        io_app_stores_0_wresp_bits, // @[:@97005.4]
  input         io_dram_cmd_ready, // @[:@97005.4]
  output        io_dram_cmd_valid, // @[:@97005.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@97005.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@97005.4]
  output        io_dram_cmd_bits_isWr, // @[:@97005.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@97005.4]
  input         io_dram_wdata_ready, // @[:@97005.4]
  output        io_dram_wdata_valid, // @[:@97005.4]
  output [63:0] io_dram_wdata_bits_wdata_0, // @[:@97005.4]
  output [63:0] io_dram_wdata_bits_wdata_1, // @[:@97005.4]
  output [63:0] io_dram_wdata_bits_wdata_2, // @[:@97005.4]
  output [63:0] io_dram_wdata_bits_wdata_3, // @[:@97005.4]
  output [63:0] io_dram_wdata_bits_wdata_4, // @[:@97005.4]
  output [63:0] io_dram_wdata_bits_wdata_5, // @[:@97005.4]
  output [63:0] io_dram_wdata_bits_wdata_6, // @[:@97005.4]
  output [63:0] io_dram_wdata_bits_wdata_7, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@97005.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@97005.4]
  output        io_dram_wdata_bits_wlast, // @[:@97005.4]
  output        io_dram_rresp_ready, // @[:@97005.4]
  input         io_dram_rresp_valid, // @[:@97005.4]
  input  [63:0] io_dram_rresp_bits_rdata_0, // @[:@97005.4]
  input  [63:0] io_dram_rresp_bits_rdata_1, // @[:@97005.4]
  input  [63:0] io_dram_rresp_bits_rdata_2, // @[:@97005.4]
  input  [63:0] io_dram_rresp_bits_rdata_3, // @[:@97005.4]
  input  [63:0] io_dram_rresp_bits_rdata_4, // @[:@97005.4]
  input  [63:0] io_dram_rresp_bits_rdata_5, // @[:@97005.4]
  input  [63:0] io_dram_rresp_bits_rdata_6, // @[:@97005.4]
  input  [63:0] io_dram_rresp_bits_rdata_7, // @[:@97005.4]
  input  [31:0] io_dram_rresp_bits_tag, // @[:@97005.4]
  output        io_dram_wresp_ready, // @[:@97005.4]
  input         io_dram_wresp_valid, // @[:@97005.4]
  input  [31:0] io_dram_wresp_bits_tag, // @[:@97005.4]
  output [31:0] io_debugSignals_0, // @[:@97005.4]
  output [31:0] io_debugSignals_1, // @[:@97005.4]
  output [31:0] io_debugSignals_2, // @[:@97005.4]
  output [31:0] io_debugSignals_3, // @[:@97005.4]
  output [31:0] io_debugSignals_4, // @[:@97005.4]
  output [31:0] io_debugSignals_5, // @[:@97005.4]
  output [31:0] io_debugSignals_6, // @[:@97005.4]
  output [31:0] io_debugSignals_7, // @[:@97005.4]
  output [31:0] io_debugSignals_8, // @[:@97005.4]
  output [31:0] io_debugSignals_9, // @[:@97005.4]
  output [31:0] io_debugSignals_10, // @[:@97005.4]
  output [31:0] io_debugSignals_11, // @[:@97005.4]
  output [31:0] io_debugSignals_12, // @[:@97005.4]
  output [31:0] io_debugSignals_13, // @[:@97005.4]
  output [31:0] io_debugSignals_14, // @[:@97005.4]
  output [31:0] io_debugSignals_15, // @[:@97005.4]
  output [31:0] io_debugSignals_16, // @[:@97005.4]
  output [31:0] io_debugSignals_17, // @[:@97005.4]
  output [31:0] io_debugSignals_18, // @[:@97005.4]
  output [31:0] io_debugSignals_19, // @[:@97005.4]
  output [31:0] io_debugSignals_20, // @[:@97005.4]
  output [31:0] io_debugSignals_21, // @[:@97005.4]
  output [31:0] io_debugSignals_22, // @[:@97005.4]
  output [31:0] io_debugSignals_23, // @[:@97005.4]
  output [31:0] io_debugSignals_24, // @[:@97005.4]
  output [31:0] io_debugSignals_25, // @[:@97005.4]
  output [31:0] io_debugSignals_26, // @[:@97005.4]
  output [31:0] io_debugSignals_27, // @[:@97005.4]
  output [31:0] io_debugSignals_28, // @[:@97005.4]
  output [31:0] io_debugSignals_29, // @[:@97005.4]
  output [31:0] io_debugSignals_30, // @[:@97005.4]
  output [31:0] io_debugSignals_41 // @[:@97005.4]
);
  wire  StreamControllerLoad_clock; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire  StreamControllerLoad_reset; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire  StreamControllerLoad_io_dram_cmd_ready; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire  StreamControllerLoad_io_dram_cmd_valid; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire [63:0] StreamControllerLoad_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire [31:0] StreamControllerLoad_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire  StreamControllerLoad_io_dram_rresp_ready; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire  StreamControllerLoad_io_dram_rresp_valid; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire [63:0] StreamControllerLoad_io_dram_rresp_bits_rdata_0; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire [63:0] StreamControllerLoad_io_dram_rresp_bits_rdata_1; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire [63:0] StreamControllerLoad_io_dram_rresp_bits_rdata_2; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire [63:0] StreamControllerLoad_io_dram_rresp_bits_rdata_3; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire [63:0] StreamControllerLoad_io_dram_rresp_bits_rdata_4; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire [63:0] StreamControllerLoad_io_dram_rresp_bits_rdata_5; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire [63:0] StreamControllerLoad_io_dram_rresp_bits_rdata_6; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire [63:0] StreamControllerLoad_io_dram_rresp_bits_rdata_7; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire  StreamControllerLoad_io_load_cmd_ready; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire  StreamControllerLoad_io_load_cmd_valid; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire [63:0] StreamControllerLoad_io_load_cmd_bits_addr; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire [31:0] StreamControllerLoad_io_load_cmd_bits_size; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire  StreamControllerLoad_io_load_data_ready; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire  StreamControllerLoad_io_load_data_valid; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire [31:0] StreamControllerLoad_io_load_data_bits_rdata_0; // @[DRAMArbiter.scala 60:21:@97828.4]
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire [63:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire [63:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire [63:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire [63:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire [63:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire [63:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire [63:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire [63:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@97838.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_rresp_valid; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_rresp_bits_rdata_0; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_rresp_bits_rdata_1; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_rresp_bits_rdata_2; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_rresp_bits_rdata_3; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_rresp_bits_rdata_4; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_rresp_bits_rdata_5; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_rresp_bits_rdata_6; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_0_rresp_bits_rdata_7; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_cmd_ready; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_cmd_valid; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_1_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [31:0] StreamArbiter_io_app_1_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [31:0] StreamArbiter_io_app_1_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_ready; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_valid; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_1_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_1_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_1_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_1_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_1_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_1_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_1_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_app_1_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_rresp_ready; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wresp_ready; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_app_1_wresp_valid; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_rresp_valid; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_rresp_bits_rdata_0; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_rresp_bits_rdata_1; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_rresp_bits_rdata_2; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_rresp_bits_rdata_3; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_rresp_bits_rdata_4; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_rresp_bits_rdata_5; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_rresp_bits_rdata_6; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [63:0] StreamArbiter_io_dram_rresp_bits_rdata_7; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [31:0] StreamArbiter_io_dram_rresp_bits_tag; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@97852.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_rresp_valid; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_rresp_bits_rdata_0; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_rresp_bits_rdata_1; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_rresp_bits_rdata_2; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_rresp_bits_rdata_3; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_rresp_bits_rdata_4; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_rresp_bits_rdata_5; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_rresp_bits_rdata_6; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_in_rresp_bits_rdata_7; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [31:0] AXICmdSplit_io_in_rresp_bits_tag; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_rresp_valid; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_rresp_bits_rdata_0; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_rresp_bits_rdata_1; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_rresp_bits_rdata_2; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_rresp_bits_rdata_3; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_rresp_bits_rdata_4; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_rresp_bits_rdata_5; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_rresp_bits_rdata_6; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [63:0] AXICmdSplit_io_out_rresp_bits_rdata_7; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [31:0] AXICmdSplit_io_out_rresp_bits_tag; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@98240.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_rresp_valid; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_rresp_bits_rdata_0; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_rresp_bits_rdata_1; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_rresp_bits_rdata_2; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_rresp_bits_rdata_3; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_rresp_bits_rdata_4; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_rresp_bits_rdata_5; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_rresp_bits_rdata_6; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_in_rresp_bits_rdata_7; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [31:0] AXICmdIssue_io_in_rresp_bits_tag; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_rresp_valid; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_rresp_bits_rdata_0; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_rresp_bits_rdata_1; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_rresp_bits_rdata_2; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_rresp_bits_rdata_3; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_rresp_bits_rdata_4; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_rresp_bits_rdata_5; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_rresp_bits_rdata_6; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [63:0] AXICmdIssue_io_out_rresp_bits_rdata_7; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [31:0] AXICmdIssue_io_out_rresp_bits_tag; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@98339.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@98339.4]
  reg [63:0] _T_1916; // @[DRAMArbiter.scala 121:24:@98538.4]
  reg [63:0] _RAND_0;
  wire [64:0] _T_1918; // @[DRAMArbiter.scala 123:18:@98540.6]
  wire [63:0] _T_1919; // @[DRAMArbiter.scala 123:18:@98541.6]
  wire [63:0] _GEN_0; // @[DRAMArbiter.scala 122:19:@98539.4]
  wire  _T_1920; // @[DRAMArbiter.scala 139:60:@98545.4]
  wire  _T_1927; // @[DRAMArbiter.scala 140:57:@98552.4]
  reg [63:0] _T_1930; // @[DRAMArbiter.scala 121:24:@98553.4]
  reg [63:0] _RAND_1;
  wire [64:0] _T_1932; // @[DRAMArbiter.scala 123:18:@98555.6]
  wire [63:0] _T_1933; // @[DRAMArbiter.scala 123:18:@98556.6]
  wire [63:0] _GEN_2; // @[DRAMArbiter.scala 122:19:@98554.4]
  wire  _T_1934; // @[DRAMArbiter.scala 141:70:@98559.4]
  reg [63:0] _T_1937; // @[DRAMArbiter.scala 121:24:@98560.4]
  reg [63:0] _RAND_2;
  wire [64:0] _T_1939; // @[DRAMArbiter.scala 123:18:@98562.6]
  wire [63:0] _T_1940; // @[DRAMArbiter.scala 123:18:@98563.6]
  wire [63:0] _GEN_3; // @[DRAMArbiter.scala 122:19:@98561.4]
  wire  _T_1941; // @[DRAMArbiter.scala 144:52:@98567.4]
  reg [63:0] _T_1944; // @[DRAMArbiter.scala 121:24:@98568.4]
  reg [63:0] _RAND_3;
  wire [64:0] _T_1946; // @[DRAMArbiter.scala 123:18:@98570.6]
  wire [63:0] _T_1947; // @[DRAMArbiter.scala 123:18:@98571.6]
  wire [63:0] _GEN_4; // @[DRAMArbiter.scala 122:19:@98569.4]
  wire  _T_1950; // @[DRAMArbiter.scala 145:74:@98576.4]
  wire  _T_1951; // @[DRAMArbiter.scala 145:72:@98577.4]
  reg [63:0] _T_1954; // @[DRAMArbiter.scala 121:24:@98578.4]
  reg [63:0] _RAND_4;
  wire [64:0] _T_1956; // @[DRAMArbiter.scala 123:18:@98580.6]
  wire [63:0] _T_1957; // @[DRAMArbiter.scala 123:18:@98581.6]
  wire [63:0] _GEN_5; // @[DRAMArbiter.scala 122:19:@98579.4]
  wire  _T_1959; // @[DRAMArbiter.scala 146:72:@98586.4]
  reg [63:0] _T_1962; // @[DRAMArbiter.scala 121:24:@98587.4]
  reg [63:0] _RAND_5;
  wire [64:0] _T_1964; // @[DRAMArbiter.scala 123:18:@98589.6]
  wire [63:0] _T_1965; // @[DRAMArbiter.scala 123:18:@98590.6]
  wire [63:0] _GEN_6; // @[DRAMArbiter.scala 122:19:@98588.4]
  wire  _T_1966; // @[DRAMArbiter.scala 150:59:@98594.4]
  wire  _T_1967; // @[DRAMArbiter.scala 150:76:@98595.4]
  reg [63:0] _T_1970; // @[DRAMArbiter.scala 121:24:@98596.4]
  reg [63:0] _RAND_6;
  wire [64:0] _T_1972; // @[DRAMArbiter.scala 123:18:@98598.6]
  wire [63:0] _T_1973; // @[DRAMArbiter.scala 123:18:@98599.6]
  wire [63:0] _GEN_7; // @[DRAMArbiter.scala 122:19:@98597.4]
  wire  _T_1974; // @[DRAMArbiter.scala 156:60:@98603.4]
  wire  _T_1975; // @[DRAMArbiter.scala 156:78:@98604.4]
  reg [63:0] _T_1978; // @[DRAMArbiter.scala 121:24:@98605.4]
  reg [63:0] _RAND_7;
  wire [64:0] _T_1980; // @[DRAMArbiter.scala 123:18:@98607.6]
  wire [63:0] _T_1981; // @[DRAMArbiter.scala 123:18:@98608.6]
  wire [63:0] _GEN_8; // @[DRAMArbiter.scala 122:19:@98606.4]
  reg [63:0] _T_1985; // @[DRAMArbiter.scala 121:24:@98613.4]
  reg [63:0] _RAND_8;
  wire [64:0] _T_1987; // @[DRAMArbiter.scala 123:18:@98615.6]
  wire [63:0] _T_1988; // @[DRAMArbiter.scala 123:18:@98616.6]
  wire [63:0] _GEN_9; // @[DRAMArbiter.scala 122:19:@98614.4]
  wire  _T_1990; // @[DRAMArbiter.scala 161:56:@98620.4]
  wire  _T_1991; // @[DRAMArbiter.scala 161:54:@98621.4]
  reg [63:0] _T_1994; // @[DRAMArbiter.scala 121:24:@98622.4]
  reg [63:0] _RAND_9;
  wire [64:0] _T_1996; // @[DRAMArbiter.scala 123:18:@98624.6]
  wire [63:0] _T_1997; // @[DRAMArbiter.scala 123:18:@98625.6]
  wire [63:0] _GEN_10; // @[DRAMArbiter.scala 122:19:@98623.4]
  wire  _T_1999; // @[DRAMArbiter.scala 162:34:@98629.4]
  wire  _T_2000; // @[DRAMArbiter.scala 162:55:@98630.4]
  reg [63:0] _T_2003; // @[DRAMArbiter.scala 121:24:@98631.4]
  reg [63:0] _RAND_10;
  wire [64:0] _T_2005; // @[DRAMArbiter.scala 123:18:@98633.6]
  wire [63:0] _T_2006; // @[DRAMArbiter.scala 123:18:@98634.6]
  wire [63:0] _GEN_11; // @[DRAMArbiter.scala 122:19:@98632.4]
  wire [7:0] _T_2013; // @[FringeBundles.scala 132:28:@98642.4]
  wire  _T_2017; // @[DRAMArbiter.scala 165:116:@98648.4]
  wire  _T_2018; // @[DRAMArbiter.scala 165:78:@98649.4]
  reg [63:0] _T_2021; // @[DRAMArbiter.scala 121:24:@98650.4]
  reg [63:0] _RAND_11;
  wire [64:0] _T_2023; // @[DRAMArbiter.scala 123:18:@98652.6]
  wire [63:0] _T_2024; // @[DRAMArbiter.scala 123:18:@98653.6]
  wire [63:0] _GEN_12; // @[DRAMArbiter.scala 122:19:@98651.4]
  wire  _T_2025; // @[DRAMArbiter.scala 167:54:@98657.4]
  reg [63:0] _T_2028; // @[DRAMArbiter.scala 121:24:@98658.4]
  reg [63:0] _RAND_12;
  wire [64:0] _T_2030; // @[DRAMArbiter.scala 123:18:@98660.6]
  wire [63:0] _T_2031; // @[DRAMArbiter.scala 123:18:@98661.6]
  wire [63:0] _GEN_13; // @[DRAMArbiter.scala 122:19:@98659.4]
  wire  _T_2033; // @[DRAMArbiter.scala 168:56:@98665.4]
  wire  _T_2034; // @[DRAMArbiter.scala 168:54:@98666.4]
  reg [63:0] _T_2037; // @[DRAMArbiter.scala 121:24:@98667.4]
  reg [63:0] _RAND_13;
  wire [64:0] _T_2039; // @[DRAMArbiter.scala 123:18:@98669.6]
  wire [63:0] _T_2040; // @[DRAMArbiter.scala 123:18:@98670.6]
  wire [63:0] _GEN_14; // @[DRAMArbiter.scala 122:19:@98668.4]
  wire  _T_2042; // @[DRAMArbiter.scala 169:34:@98674.4]
  wire  _T_2043; // @[DRAMArbiter.scala 169:55:@98675.4]
  reg [63:0] _T_2046; // @[DRAMArbiter.scala 121:24:@98676.4]
  reg [63:0] _RAND_14;
  wire [64:0] _T_2048; // @[DRAMArbiter.scala 123:18:@98678.6]
  wire [63:0] _T_2049; // @[DRAMArbiter.scala 123:18:@98679.6]
  wire [63:0] _GEN_15; // @[DRAMArbiter.scala 122:19:@98677.4]
  wire [7:0] _T_2056; // @[FringeBundles.scala 140:28:@98687.4]
  wire  _T_2060; // @[DRAMArbiter.scala 172:116:@98693.4]
  wire  _T_2061; // @[DRAMArbiter.scala 172:78:@98694.4]
  reg [63:0] _T_2064; // @[DRAMArbiter.scala 121:24:@98695.4]
  reg [63:0] _RAND_15;
  wire [64:0] _T_2066; // @[DRAMArbiter.scala 123:18:@98697.6]
  wire [63:0] _T_2067; // @[DRAMArbiter.scala 123:18:@98698.6]
  wire [63:0] _GEN_16; // @[DRAMArbiter.scala 122:19:@98696.4]
  wire  _T_2068; // @[DRAMArbiter.scala 176:70:@98702.4]
  reg [63:0] _T_2070; // @[DRAMArbiter.scala 129:25:@98703.4]
  reg [63:0] _RAND_16;
  wire [63:0] _GEN_17; // @[DRAMArbiter.scala 130:19:@98704.4]
  reg [31:0] _T_2073; // @[DRAMArbiter.scala 129:25:@98709.4]
  reg [31:0] _RAND_17;
  wire [31:0] _GEN_18; // @[DRAMArbiter.scala 130:19:@98710.4]
  reg [63:0] _T_2076; // @[DRAMArbiter.scala 129:25:@98715.4]
  reg [63:0] _RAND_18;
  wire [63:0] _GEN_19; // @[DRAMArbiter.scala 130:19:@98716.4]
  reg  _T_2079; // @[DRAMArbiter.scala 129:25:@98721.4]
  reg [31:0] _RAND_19;
  wire  _GEN_20; // @[DRAMArbiter.scala 130:19:@98722.4]
  wire  _T_2082; // @[DRAMArbiter.scala 180:115:@98727.4]
  wire  _T_2083; // @[DRAMArbiter.scala 180:102:@98728.4]
  reg [63:0] _T_2085; // @[DRAMArbiter.scala 129:25:@98729.4]
  reg [63:0] _RAND_20;
  wire [63:0] _GEN_21; // @[DRAMArbiter.scala 130:19:@98730.4]
  reg  _T_2091; // @[DRAMArbiter.scala 129:25:@98737.4]
  reg [31:0] _RAND_21;
  wire  _GEN_22; // @[DRAMArbiter.scala 130:19:@98738.4]
  wire  _T_2094; // @[DRAMArbiter.scala 182:115:@98743.4]
  wire  _T_2095; // @[DRAMArbiter.scala 182:102:@98744.4]
  reg [63:0] _T_2097; // @[DRAMArbiter.scala 129:25:@98745.4]
  reg [63:0] _RAND_22;
  wire [63:0] _GEN_23; // @[DRAMArbiter.scala 130:19:@98746.4]
  reg  _T_2103; // @[DRAMArbiter.scala 129:25:@98753.4]
  reg [31:0] _RAND_23;
  wire  _GEN_24; // @[DRAMArbiter.scala 130:19:@98754.4]
  wire  _T_2104; // @[DRAMArbiter.scala 184:92:@98758.4]
  reg [63:0] _T_2106; // @[DRAMArbiter.scala 129:25:@98759.4]
  reg [63:0] _RAND_24;
  wire [63:0] _GEN_25; // @[DRAMArbiter.scala 130:19:@98760.4]
  reg [31:0] _T_2109; // @[DRAMArbiter.scala 129:25:@98765.4]
  reg [31:0] _RAND_25;
  wire [31:0] _GEN_26; // @[DRAMArbiter.scala 130:19:@98766.4]
  reg [31:0] _T_2112; // @[DRAMArbiter.scala 129:25:@98771.4]
  reg [31:0] _RAND_26;
  wire [31:0] _GEN_27; // @[DRAMArbiter.scala 130:19:@98772.4]
  reg  _T_2115; // @[DRAMArbiter.scala 129:25:@98777.4]
  reg [31:0] _RAND_27;
  wire  _GEN_28; // @[DRAMArbiter.scala 130:19:@98778.4]
  wire  _T_2118; // @[DRAMArbiter.scala 188:148:@98783.4]
  wire  _T_2119; // @[DRAMArbiter.scala 188:132:@98784.4]
  reg [31:0] _T_2121; // @[DRAMArbiter.scala 129:25:@98785.4]
  reg [31:0] _RAND_28;
  wire [31:0] _GEN_29; // @[DRAMArbiter.scala 130:19:@98786.4]
  reg  _T_2127; // @[DRAMArbiter.scala 129:25:@98793.4]
  reg [31:0] _RAND_29;
  wire  _GEN_30; // @[DRAMArbiter.scala 130:19:@98794.4]
  wire  _T_2130; // @[DRAMArbiter.scala 190:148:@98799.4]
  wire  _T_2131; // @[DRAMArbiter.scala 190:132:@98800.4]
  reg [31:0] _T_2133; // @[DRAMArbiter.scala 129:25:@98801.4]
  reg [31:0] _RAND_30;
  wire [31:0] _GEN_31; // @[DRAMArbiter.scala 130:19:@98802.4]
  reg  _T_2139; // @[DRAMArbiter.scala 129:25:@98809.4]
  reg [31:0] _RAND_31;
  wire  _GEN_32; // @[DRAMArbiter.scala 130:19:@98810.4]
  reg [63:0] _T_2211; // @[DRAMArbiter.scala 121:24:@98891.4]
  reg [63:0] _RAND_32;
  wire [64:0] _T_2213; // @[DRAMArbiter.scala 123:18:@98893.6]
  wire [63:0] _T_2214; // @[DRAMArbiter.scala 123:18:@98894.6]
  StreamControllerLoad StreamControllerLoad ( // @[DRAMArbiter.scala 60:21:@97828.4]
    .clock(StreamControllerLoad_clock),
    .reset(StreamControllerLoad_reset),
    .io_dram_cmd_ready(StreamControllerLoad_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerLoad_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerLoad_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerLoad_io_dram_cmd_bits_size),
    .io_dram_rresp_ready(StreamControllerLoad_io_dram_rresp_ready),
    .io_dram_rresp_valid(StreamControllerLoad_io_dram_rresp_valid),
    .io_dram_rresp_bits_rdata_0(StreamControllerLoad_io_dram_rresp_bits_rdata_0),
    .io_dram_rresp_bits_rdata_1(StreamControllerLoad_io_dram_rresp_bits_rdata_1),
    .io_dram_rresp_bits_rdata_2(StreamControllerLoad_io_dram_rresp_bits_rdata_2),
    .io_dram_rresp_bits_rdata_3(StreamControllerLoad_io_dram_rresp_bits_rdata_3),
    .io_dram_rresp_bits_rdata_4(StreamControllerLoad_io_dram_rresp_bits_rdata_4),
    .io_dram_rresp_bits_rdata_5(StreamControllerLoad_io_dram_rresp_bits_rdata_5),
    .io_dram_rresp_bits_rdata_6(StreamControllerLoad_io_dram_rresp_bits_rdata_6),
    .io_dram_rresp_bits_rdata_7(StreamControllerLoad_io_dram_rresp_bits_rdata_7),
    .io_load_cmd_ready(StreamControllerLoad_io_load_cmd_ready),
    .io_load_cmd_valid(StreamControllerLoad_io_load_cmd_valid),
    .io_load_cmd_bits_addr(StreamControllerLoad_io_load_cmd_bits_addr),
    .io_load_cmd_bits_size(StreamControllerLoad_io_load_cmd_bits_size),
    .io_load_data_ready(StreamControllerLoad_io_load_data_ready),
    .io_load_data_valid(StreamControllerLoad_io_load_data_valid),
    .io_load_data_bits_rdata_0(StreamControllerLoad_io_load_data_bits_rdata_0)
  );
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@97838.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@97852.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_rresp_valid(StreamArbiter_io_app_0_rresp_valid),
    .io_app_0_rresp_bits_rdata_0(StreamArbiter_io_app_0_rresp_bits_rdata_0),
    .io_app_0_rresp_bits_rdata_1(StreamArbiter_io_app_0_rresp_bits_rdata_1),
    .io_app_0_rresp_bits_rdata_2(StreamArbiter_io_app_0_rresp_bits_rdata_2),
    .io_app_0_rresp_bits_rdata_3(StreamArbiter_io_app_0_rresp_bits_rdata_3),
    .io_app_0_rresp_bits_rdata_4(StreamArbiter_io_app_0_rresp_bits_rdata_4),
    .io_app_0_rresp_bits_rdata_5(StreamArbiter_io_app_0_rresp_bits_rdata_5),
    .io_app_0_rresp_bits_rdata_6(StreamArbiter_io_app_0_rresp_bits_rdata_6),
    .io_app_0_rresp_bits_rdata_7(StreamArbiter_io_app_0_rresp_bits_rdata_7),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_1_cmd_ready(StreamArbiter_io_app_1_cmd_ready),
    .io_app_1_cmd_valid(StreamArbiter_io_app_1_cmd_valid),
    .io_app_1_cmd_bits_addr(StreamArbiter_io_app_1_cmd_bits_addr),
    .io_app_1_cmd_bits_size(StreamArbiter_io_app_1_cmd_bits_size),
    .io_app_1_cmd_bits_isWr(StreamArbiter_io_app_1_cmd_bits_isWr),
    .io_app_1_cmd_bits_tag(StreamArbiter_io_app_1_cmd_bits_tag),
    .io_app_1_wdata_ready(StreamArbiter_io_app_1_wdata_ready),
    .io_app_1_wdata_valid(StreamArbiter_io_app_1_wdata_valid),
    .io_app_1_wdata_bits_wdata_0(StreamArbiter_io_app_1_wdata_bits_wdata_0),
    .io_app_1_wdata_bits_wdata_1(StreamArbiter_io_app_1_wdata_bits_wdata_1),
    .io_app_1_wdata_bits_wdata_2(StreamArbiter_io_app_1_wdata_bits_wdata_2),
    .io_app_1_wdata_bits_wdata_3(StreamArbiter_io_app_1_wdata_bits_wdata_3),
    .io_app_1_wdata_bits_wdata_4(StreamArbiter_io_app_1_wdata_bits_wdata_4),
    .io_app_1_wdata_bits_wdata_5(StreamArbiter_io_app_1_wdata_bits_wdata_5),
    .io_app_1_wdata_bits_wdata_6(StreamArbiter_io_app_1_wdata_bits_wdata_6),
    .io_app_1_wdata_bits_wdata_7(StreamArbiter_io_app_1_wdata_bits_wdata_7),
    .io_app_1_wdata_bits_wstrb_0(StreamArbiter_io_app_1_wdata_bits_wstrb_0),
    .io_app_1_wdata_bits_wstrb_1(StreamArbiter_io_app_1_wdata_bits_wstrb_1),
    .io_app_1_wdata_bits_wstrb_2(StreamArbiter_io_app_1_wdata_bits_wstrb_2),
    .io_app_1_wdata_bits_wstrb_3(StreamArbiter_io_app_1_wdata_bits_wstrb_3),
    .io_app_1_wdata_bits_wstrb_4(StreamArbiter_io_app_1_wdata_bits_wstrb_4),
    .io_app_1_wdata_bits_wstrb_5(StreamArbiter_io_app_1_wdata_bits_wstrb_5),
    .io_app_1_wdata_bits_wstrb_6(StreamArbiter_io_app_1_wdata_bits_wstrb_6),
    .io_app_1_wdata_bits_wstrb_7(StreamArbiter_io_app_1_wdata_bits_wstrb_7),
    .io_app_1_wdata_bits_wstrb_8(StreamArbiter_io_app_1_wdata_bits_wstrb_8),
    .io_app_1_wdata_bits_wstrb_9(StreamArbiter_io_app_1_wdata_bits_wstrb_9),
    .io_app_1_wdata_bits_wstrb_10(StreamArbiter_io_app_1_wdata_bits_wstrb_10),
    .io_app_1_wdata_bits_wstrb_11(StreamArbiter_io_app_1_wdata_bits_wstrb_11),
    .io_app_1_wdata_bits_wstrb_12(StreamArbiter_io_app_1_wdata_bits_wstrb_12),
    .io_app_1_wdata_bits_wstrb_13(StreamArbiter_io_app_1_wdata_bits_wstrb_13),
    .io_app_1_wdata_bits_wstrb_14(StreamArbiter_io_app_1_wdata_bits_wstrb_14),
    .io_app_1_wdata_bits_wstrb_15(StreamArbiter_io_app_1_wdata_bits_wstrb_15),
    .io_app_1_wdata_bits_wstrb_16(StreamArbiter_io_app_1_wdata_bits_wstrb_16),
    .io_app_1_wdata_bits_wstrb_17(StreamArbiter_io_app_1_wdata_bits_wstrb_17),
    .io_app_1_wdata_bits_wstrb_18(StreamArbiter_io_app_1_wdata_bits_wstrb_18),
    .io_app_1_wdata_bits_wstrb_19(StreamArbiter_io_app_1_wdata_bits_wstrb_19),
    .io_app_1_wdata_bits_wstrb_20(StreamArbiter_io_app_1_wdata_bits_wstrb_20),
    .io_app_1_wdata_bits_wstrb_21(StreamArbiter_io_app_1_wdata_bits_wstrb_21),
    .io_app_1_wdata_bits_wstrb_22(StreamArbiter_io_app_1_wdata_bits_wstrb_22),
    .io_app_1_wdata_bits_wstrb_23(StreamArbiter_io_app_1_wdata_bits_wstrb_23),
    .io_app_1_wdata_bits_wstrb_24(StreamArbiter_io_app_1_wdata_bits_wstrb_24),
    .io_app_1_wdata_bits_wstrb_25(StreamArbiter_io_app_1_wdata_bits_wstrb_25),
    .io_app_1_wdata_bits_wstrb_26(StreamArbiter_io_app_1_wdata_bits_wstrb_26),
    .io_app_1_wdata_bits_wstrb_27(StreamArbiter_io_app_1_wdata_bits_wstrb_27),
    .io_app_1_wdata_bits_wstrb_28(StreamArbiter_io_app_1_wdata_bits_wstrb_28),
    .io_app_1_wdata_bits_wstrb_29(StreamArbiter_io_app_1_wdata_bits_wstrb_29),
    .io_app_1_wdata_bits_wstrb_30(StreamArbiter_io_app_1_wdata_bits_wstrb_30),
    .io_app_1_wdata_bits_wstrb_31(StreamArbiter_io_app_1_wdata_bits_wstrb_31),
    .io_app_1_wdata_bits_wstrb_32(StreamArbiter_io_app_1_wdata_bits_wstrb_32),
    .io_app_1_wdata_bits_wstrb_33(StreamArbiter_io_app_1_wdata_bits_wstrb_33),
    .io_app_1_wdata_bits_wstrb_34(StreamArbiter_io_app_1_wdata_bits_wstrb_34),
    .io_app_1_wdata_bits_wstrb_35(StreamArbiter_io_app_1_wdata_bits_wstrb_35),
    .io_app_1_wdata_bits_wstrb_36(StreamArbiter_io_app_1_wdata_bits_wstrb_36),
    .io_app_1_wdata_bits_wstrb_37(StreamArbiter_io_app_1_wdata_bits_wstrb_37),
    .io_app_1_wdata_bits_wstrb_38(StreamArbiter_io_app_1_wdata_bits_wstrb_38),
    .io_app_1_wdata_bits_wstrb_39(StreamArbiter_io_app_1_wdata_bits_wstrb_39),
    .io_app_1_wdata_bits_wstrb_40(StreamArbiter_io_app_1_wdata_bits_wstrb_40),
    .io_app_1_wdata_bits_wstrb_41(StreamArbiter_io_app_1_wdata_bits_wstrb_41),
    .io_app_1_wdata_bits_wstrb_42(StreamArbiter_io_app_1_wdata_bits_wstrb_42),
    .io_app_1_wdata_bits_wstrb_43(StreamArbiter_io_app_1_wdata_bits_wstrb_43),
    .io_app_1_wdata_bits_wstrb_44(StreamArbiter_io_app_1_wdata_bits_wstrb_44),
    .io_app_1_wdata_bits_wstrb_45(StreamArbiter_io_app_1_wdata_bits_wstrb_45),
    .io_app_1_wdata_bits_wstrb_46(StreamArbiter_io_app_1_wdata_bits_wstrb_46),
    .io_app_1_wdata_bits_wstrb_47(StreamArbiter_io_app_1_wdata_bits_wstrb_47),
    .io_app_1_wdata_bits_wstrb_48(StreamArbiter_io_app_1_wdata_bits_wstrb_48),
    .io_app_1_wdata_bits_wstrb_49(StreamArbiter_io_app_1_wdata_bits_wstrb_49),
    .io_app_1_wdata_bits_wstrb_50(StreamArbiter_io_app_1_wdata_bits_wstrb_50),
    .io_app_1_wdata_bits_wstrb_51(StreamArbiter_io_app_1_wdata_bits_wstrb_51),
    .io_app_1_wdata_bits_wstrb_52(StreamArbiter_io_app_1_wdata_bits_wstrb_52),
    .io_app_1_wdata_bits_wstrb_53(StreamArbiter_io_app_1_wdata_bits_wstrb_53),
    .io_app_1_wdata_bits_wstrb_54(StreamArbiter_io_app_1_wdata_bits_wstrb_54),
    .io_app_1_wdata_bits_wstrb_55(StreamArbiter_io_app_1_wdata_bits_wstrb_55),
    .io_app_1_wdata_bits_wstrb_56(StreamArbiter_io_app_1_wdata_bits_wstrb_56),
    .io_app_1_wdata_bits_wstrb_57(StreamArbiter_io_app_1_wdata_bits_wstrb_57),
    .io_app_1_wdata_bits_wstrb_58(StreamArbiter_io_app_1_wdata_bits_wstrb_58),
    .io_app_1_wdata_bits_wstrb_59(StreamArbiter_io_app_1_wdata_bits_wstrb_59),
    .io_app_1_wdata_bits_wstrb_60(StreamArbiter_io_app_1_wdata_bits_wstrb_60),
    .io_app_1_wdata_bits_wstrb_61(StreamArbiter_io_app_1_wdata_bits_wstrb_61),
    .io_app_1_wdata_bits_wstrb_62(StreamArbiter_io_app_1_wdata_bits_wstrb_62),
    .io_app_1_wdata_bits_wstrb_63(StreamArbiter_io_app_1_wdata_bits_wstrb_63),
    .io_app_1_rresp_ready(StreamArbiter_io_app_1_rresp_ready),
    .io_app_1_wresp_ready(StreamArbiter_io_app_1_wresp_ready),
    .io_app_1_wresp_valid(StreamArbiter_io_app_1_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_rresp_valid(StreamArbiter_io_dram_rresp_valid),
    .io_dram_rresp_bits_rdata_0(StreamArbiter_io_dram_rresp_bits_rdata_0),
    .io_dram_rresp_bits_rdata_1(StreamArbiter_io_dram_rresp_bits_rdata_1),
    .io_dram_rresp_bits_rdata_2(StreamArbiter_io_dram_rresp_bits_rdata_2),
    .io_dram_rresp_bits_rdata_3(StreamArbiter_io_dram_rresp_bits_rdata_3),
    .io_dram_rresp_bits_rdata_4(StreamArbiter_io_dram_rresp_bits_rdata_4),
    .io_dram_rresp_bits_rdata_5(StreamArbiter_io_dram_rresp_bits_rdata_5),
    .io_dram_rresp_bits_rdata_6(StreamArbiter_io_dram_rresp_bits_rdata_6),
    .io_dram_rresp_bits_rdata_7(StreamArbiter_io_dram_rresp_bits_rdata_7),
    .io_dram_rresp_bits_tag(StreamArbiter_io_dram_rresp_bits_tag),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@98240.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_rresp_valid(AXICmdSplit_io_in_rresp_valid),
    .io_in_rresp_bits_rdata_0(AXICmdSplit_io_in_rresp_bits_rdata_0),
    .io_in_rresp_bits_rdata_1(AXICmdSplit_io_in_rresp_bits_rdata_1),
    .io_in_rresp_bits_rdata_2(AXICmdSplit_io_in_rresp_bits_rdata_2),
    .io_in_rresp_bits_rdata_3(AXICmdSplit_io_in_rresp_bits_rdata_3),
    .io_in_rresp_bits_rdata_4(AXICmdSplit_io_in_rresp_bits_rdata_4),
    .io_in_rresp_bits_rdata_5(AXICmdSplit_io_in_rresp_bits_rdata_5),
    .io_in_rresp_bits_rdata_6(AXICmdSplit_io_in_rresp_bits_rdata_6),
    .io_in_rresp_bits_rdata_7(AXICmdSplit_io_in_rresp_bits_rdata_7),
    .io_in_rresp_bits_tag(AXICmdSplit_io_in_rresp_bits_tag),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_rresp_valid(AXICmdSplit_io_out_rresp_valid),
    .io_out_rresp_bits_rdata_0(AXICmdSplit_io_out_rresp_bits_rdata_0),
    .io_out_rresp_bits_rdata_1(AXICmdSplit_io_out_rresp_bits_rdata_1),
    .io_out_rresp_bits_rdata_2(AXICmdSplit_io_out_rresp_bits_rdata_2),
    .io_out_rresp_bits_rdata_3(AXICmdSplit_io_out_rresp_bits_rdata_3),
    .io_out_rresp_bits_rdata_4(AXICmdSplit_io_out_rresp_bits_rdata_4),
    .io_out_rresp_bits_rdata_5(AXICmdSplit_io_out_rresp_bits_rdata_5),
    .io_out_rresp_bits_rdata_6(AXICmdSplit_io_out_rresp_bits_rdata_6),
    .io_out_rresp_bits_rdata_7(AXICmdSplit_io_out_rresp_bits_rdata_7),
    .io_out_rresp_bits_tag(AXICmdSplit_io_out_rresp_bits_tag),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@98339.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_rresp_valid(AXICmdIssue_io_in_rresp_valid),
    .io_in_rresp_bits_rdata_0(AXICmdIssue_io_in_rresp_bits_rdata_0),
    .io_in_rresp_bits_rdata_1(AXICmdIssue_io_in_rresp_bits_rdata_1),
    .io_in_rresp_bits_rdata_2(AXICmdIssue_io_in_rresp_bits_rdata_2),
    .io_in_rresp_bits_rdata_3(AXICmdIssue_io_in_rresp_bits_rdata_3),
    .io_in_rresp_bits_rdata_4(AXICmdIssue_io_in_rresp_bits_rdata_4),
    .io_in_rresp_bits_rdata_5(AXICmdIssue_io_in_rresp_bits_rdata_5),
    .io_in_rresp_bits_rdata_6(AXICmdIssue_io_in_rresp_bits_rdata_6),
    .io_in_rresp_bits_rdata_7(AXICmdIssue_io_in_rresp_bits_rdata_7),
    .io_in_rresp_bits_tag(AXICmdIssue_io_in_rresp_bits_tag),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_rresp_valid(AXICmdIssue_io_out_rresp_valid),
    .io_out_rresp_bits_rdata_0(AXICmdIssue_io_out_rresp_bits_rdata_0),
    .io_out_rresp_bits_rdata_1(AXICmdIssue_io_out_rresp_bits_rdata_1),
    .io_out_rresp_bits_rdata_2(AXICmdIssue_io_out_rresp_bits_rdata_2),
    .io_out_rresp_bits_rdata_3(AXICmdIssue_io_out_rresp_bits_rdata_3),
    .io_out_rresp_bits_rdata_4(AXICmdIssue_io_out_rresp_bits_rdata_4),
    .io_out_rresp_bits_rdata_5(AXICmdIssue_io_out_rresp_bits_rdata_5),
    .io_out_rresp_bits_rdata_6(AXICmdIssue_io_out_rresp_bits_rdata_6),
    .io_out_rresp_bits_rdata_7(AXICmdIssue_io_out_rresp_bits_rdata_7),
    .io_out_rresp_bits_tag(AXICmdIssue_io_out_rresp_bits_tag),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign _T_1918 = _T_1916 + 64'h1; // @[DRAMArbiter.scala 123:18:@98540.6]
  assign _T_1919 = _T_1916 + 64'h1; // @[DRAMArbiter.scala 123:18:@98541.6]
  assign _GEN_0 = io_enable ? _T_1919 : _T_1916; // @[DRAMArbiter.scala 122:19:@98539.4]
  assign _T_1920 = io_dram_rresp_valid & io_dram_rresp_ready; // @[DRAMArbiter.scala 139:60:@98545.4]
  assign _T_1927 = io_dram_wdata_valid & io_dram_wdata_ready; // @[DRAMArbiter.scala 140:57:@98552.4]
  assign _T_1932 = _T_1930 + 64'h1; // @[DRAMArbiter.scala 123:18:@98555.6]
  assign _T_1933 = _T_1930 + 64'h1; // @[DRAMArbiter.scala 123:18:@98556.6]
  assign _GEN_2 = _T_1927 ? _T_1933 : _T_1930; // @[DRAMArbiter.scala 122:19:@98554.4]
  assign _T_1934 = io_app_stores_0_data_valid & io_app_stores_0_data_ready; // @[DRAMArbiter.scala 141:70:@98559.4]
  assign _T_1939 = _T_1937 + 64'h1; // @[DRAMArbiter.scala 123:18:@98562.6]
  assign _T_1940 = _T_1937 + 64'h1; // @[DRAMArbiter.scala 123:18:@98563.6]
  assign _GEN_3 = _T_1934 ? _T_1940 : _T_1937; // @[DRAMArbiter.scala 122:19:@98561.4]
  assign _T_1941 = io_dram_cmd_ready & io_dram_cmd_valid; // @[DRAMArbiter.scala 144:52:@98567.4]
  assign _T_1946 = _T_1944 + 64'h1; // @[DRAMArbiter.scala 123:18:@98570.6]
  assign _T_1947 = _T_1944 + 64'h1; // @[DRAMArbiter.scala 123:18:@98571.6]
  assign _GEN_4 = _T_1941 ? _T_1947 : _T_1944; // @[DRAMArbiter.scala 122:19:@98569.4]
  assign _T_1950 = io_dram_cmd_bits_isWr == 1'h0; // @[DRAMArbiter.scala 145:74:@98576.4]
  assign _T_1951 = _T_1941 & _T_1950; // @[DRAMArbiter.scala 145:72:@98577.4]
  assign _T_1956 = _T_1954 + 64'h1; // @[DRAMArbiter.scala 123:18:@98580.6]
  assign _T_1957 = _T_1954 + 64'h1; // @[DRAMArbiter.scala 123:18:@98581.6]
  assign _GEN_5 = _T_1951 ? _T_1957 : _T_1954; // @[DRAMArbiter.scala 122:19:@98579.4]
  assign _T_1959 = _T_1941 & io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 146:72:@98586.4]
  assign _T_1964 = _T_1962 + 64'h1; // @[DRAMArbiter.scala 123:18:@98589.6]
  assign _T_1965 = _T_1962 + 64'h1; // @[DRAMArbiter.scala 123:18:@98590.6]
  assign _GEN_6 = _T_1959 ? _T_1965 : _T_1962; // @[DRAMArbiter.scala 122:19:@98588.4]
  assign _T_1966 = io_enable & io_app_loads_0_cmd_valid; // @[DRAMArbiter.scala 150:59:@98594.4]
  assign _T_1967 = _T_1966 & io_app_loads_0_cmd_ready; // @[DRAMArbiter.scala 150:76:@98595.4]
  assign _T_1972 = _T_1970 + 64'h1; // @[DRAMArbiter.scala 123:18:@98598.6]
  assign _T_1973 = _T_1970 + 64'h1; // @[DRAMArbiter.scala 123:18:@98599.6]
  assign _GEN_7 = _T_1967 ? _T_1973 : _T_1970; // @[DRAMArbiter.scala 122:19:@98597.4]
  assign _T_1974 = io_enable & io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 156:60:@98603.4]
  assign _T_1975 = _T_1974 & io_app_stores_0_cmd_ready; // @[DRAMArbiter.scala 156:78:@98604.4]
  assign _T_1980 = _T_1978 + 64'h1; // @[DRAMArbiter.scala 123:18:@98607.6]
  assign _T_1981 = _T_1978 + 64'h1; // @[DRAMArbiter.scala 123:18:@98608.6]
  assign _GEN_8 = _T_1975 ? _T_1981 : _T_1978; // @[DRAMArbiter.scala 122:19:@98606.4]
  assign _T_1987 = _T_1985 + 64'h1; // @[DRAMArbiter.scala 123:18:@98615.6]
  assign _T_1988 = _T_1985 + 64'h1; // @[DRAMArbiter.scala 123:18:@98616.6]
  assign _GEN_9 = _T_1920 ? _T_1988 : _T_1985; // @[DRAMArbiter.scala 122:19:@98614.4]
  assign _T_1990 = io_dram_rresp_ready == 1'h0; // @[DRAMArbiter.scala 161:56:@98620.4]
  assign _T_1991 = io_dram_rresp_valid & _T_1990; // @[DRAMArbiter.scala 161:54:@98621.4]
  assign _T_1996 = _T_1994 + 64'h1; // @[DRAMArbiter.scala 123:18:@98624.6]
  assign _T_1997 = _T_1994 + 64'h1; // @[DRAMArbiter.scala 123:18:@98625.6]
  assign _GEN_10 = _T_1991 ? _T_1997 : _T_1994; // @[DRAMArbiter.scala 122:19:@98623.4]
  assign _T_1999 = io_dram_rresp_valid == 1'h0; // @[DRAMArbiter.scala 162:34:@98629.4]
  assign _T_2000 = _T_1999 & io_dram_rresp_ready; // @[DRAMArbiter.scala 162:55:@98630.4]
  assign _T_2005 = _T_2003 + 64'h1; // @[DRAMArbiter.scala 123:18:@98633.6]
  assign _T_2006 = _T_2003 + 64'h1; // @[DRAMArbiter.scala 123:18:@98634.6]
  assign _GEN_11 = _T_2000 ? _T_2006 : _T_2003; // @[DRAMArbiter.scala 122:19:@98632.4]
  assign _T_2013 = io_dram_rresp_bits_tag[7:0]; // @[FringeBundles.scala 132:28:@98642.4]
  assign _T_2017 = _T_2013 == 8'h0; // @[DRAMArbiter.scala 165:116:@98648.4]
  assign _T_2018 = _T_1920 & _T_2017; // @[DRAMArbiter.scala 165:78:@98649.4]
  assign _T_2023 = _T_2021 + 64'h1; // @[DRAMArbiter.scala 123:18:@98652.6]
  assign _T_2024 = _T_2021 + 64'h1; // @[DRAMArbiter.scala 123:18:@98653.6]
  assign _GEN_12 = _T_2018 ? _T_2024 : _T_2021; // @[DRAMArbiter.scala 122:19:@98651.4]
  assign _T_2025 = io_dram_wresp_valid & io_dram_wresp_ready; // @[DRAMArbiter.scala 167:54:@98657.4]
  assign _T_2030 = _T_2028 + 64'h1; // @[DRAMArbiter.scala 123:18:@98660.6]
  assign _T_2031 = _T_2028 + 64'h1; // @[DRAMArbiter.scala 123:18:@98661.6]
  assign _GEN_13 = _T_2025 ? _T_2031 : _T_2028; // @[DRAMArbiter.scala 122:19:@98659.4]
  assign _T_2033 = io_dram_wresp_ready == 1'h0; // @[DRAMArbiter.scala 168:56:@98665.4]
  assign _T_2034 = io_dram_wresp_valid & _T_2033; // @[DRAMArbiter.scala 168:54:@98666.4]
  assign _T_2039 = _T_2037 + 64'h1; // @[DRAMArbiter.scala 123:18:@98669.6]
  assign _T_2040 = _T_2037 + 64'h1; // @[DRAMArbiter.scala 123:18:@98670.6]
  assign _GEN_14 = _T_2034 ? _T_2040 : _T_2037; // @[DRAMArbiter.scala 122:19:@98668.4]
  assign _T_2042 = io_dram_wresp_valid == 1'h0; // @[DRAMArbiter.scala 169:34:@98674.4]
  assign _T_2043 = _T_2042 & io_dram_wresp_ready; // @[DRAMArbiter.scala 169:55:@98675.4]
  assign _T_2048 = _T_2046 + 64'h1; // @[DRAMArbiter.scala 123:18:@98678.6]
  assign _T_2049 = _T_2046 + 64'h1; // @[DRAMArbiter.scala 123:18:@98679.6]
  assign _GEN_15 = _T_2043 ? _T_2049 : _T_2046; // @[DRAMArbiter.scala 122:19:@98677.4]
  assign _T_2056 = io_dram_wresp_bits_tag[7:0]; // @[FringeBundles.scala 140:28:@98687.4]
  assign _T_2060 = _T_2056 == 8'h1; // @[DRAMArbiter.scala 172:116:@98693.4]
  assign _T_2061 = _T_2025 & _T_2060; // @[DRAMArbiter.scala 172:78:@98694.4]
  assign _T_2066 = _T_2064 + 64'h1; // @[DRAMArbiter.scala 123:18:@98697.6]
  assign _T_2067 = _T_2064 + 64'h1; // @[DRAMArbiter.scala 123:18:@98698.6]
  assign _GEN_16 = _T_2061 ? _T_2067 : _T_2064; // @[DRAMArbiter.scala 122:19:@98696.4]
  assign _T_2068 = io_dram_cmd_valid & io_dram_cmd_ready; // @[DRAMArbiter.scala 176:70:@98702.4]
  assign _GEN_17 = _T_2068 ? io_dram_cmd_bits_addr : _T_2070; // @[DRAMArbiter.scala 130:19:@98704.4]
  assign _GEN_18 = _T_2068 ? io_dram_cmd_bits_size : _T_2073; // @[DRAMArbiter.scala 130:19:@98710.4]
  assign _GEN_19 = _T_1927 ? io_dram_wdata_bits_wdata_0 : _T_2076; // @[DRAMArbiter.scala 130:19:@98716.4]
  assign _GEN_20 = _T_1927 ? io_dram_wdata_bits_wstrb_0 : _T_2079; // @[DRAMArbiter.scala 130:19:@98722.4]
  assign _T_2082 = _T_1930 == 64'h0; // @[DRAMArbiter.scala 180:115:@98727.4]
  assign _T_2083 = _T_1927 & _T_2082; // @[DRAMArbiter.scala 180:102:@98728.4]
  assign _GEN_21 = _T_2083 ? io_dram_wdata_bits_wdata_0 : _T_2085; // @[DRAMArbiter.scala 130:19:@98730.4]
  assign _GEN_22 = _T_2083 ? io_dram_wdata_bits_wstrb_0 : _T_2091; // @[DRAMArbiter.scala 130:19:@98738.4]
  assign _T_2094 = _T_1930 == 64'h1; // @[DRAMArbiter.scala 182:115:@98743.4]
  assign _T_2095 = _T_1927 & _T_2094; // @[DRAMArbiter.scala 182:102:@98744.4]
  assign _GEN_23 = _T_2095 ? io_dram_wdata_bits_wdata_0 : _T_2097; // @[DRAMArbiter.scala 130:19:@98746.4]
  assign _GEN_24 = _T_2095 ? io_dram_wdata_bits_wstrb_0 : _T_2103; // @[DRAMArbiter.scala 130:19:@98754.4]
  assign _T_2104 = io_app_stores_0_cmd_valid & io_app_stores_0_cmd_ready; // @[DRAMArbiter.scala 184:92:@98758.4]
  assign _GEN_25 = _T_2104 ? io_app_stores_0_cmd_bits_addr : _T_2106; // @[DRAMArbiter.scala 130:19:@98760.4]
  assign _GEN_26 = _T_2104 ? io_app_stores_0_cmd_bits_size : _T_2109; // @[DRAMArbiter.scala 130:19:@98766.4]
  assign _GEN_27 = _T_1934 ? io_app_stores_0_data_bits_wdata_0 : _T_2112; // @[DRAMArbiter.scala 130:19:@98772.4]
  assign _GEN_28 = _T_1934 ? io_app_stores_0_data_bits_wstrb : _T_2115; // @[DRAMArbiter.scala 130:19:@98778.4]
  assign _T_2118 = _T_1937 == 64'h0; // @[DRAMArbiter.scala 188:148:@98783.4]
  assign _T_2119 = _T_1934 & _T_2118; // @[DRAMArbiter.scala 188:132:@98784.4]
  assign _GEN_29 = _T_2119 ? io_app_stores_0_data_bits_wdata_0 : _T_2121; // @[DRAMArbiter.scala 130:19:@98786.4]
  assign _GEN_30 = _T_2119 ? io_app_stores_0_data_bits_wstrb : _T_2127; // @[DRAMArbiter.scala 130:19:@98794.4]
  assign _T_2130 = _T_1937 == 64'h1; // @[DRAMArbiter.scala 190:148:@98799.4]
  assign _T_2131 = _T_1934 & _T_2130; // @[DRAMArbiter.scala 190:132:@98800.4]
  assign _GEN_31 = _T_2131 ? io_app_stores_0_data_bits_wdata_0 : _T_2133; // @[DRAMArbiter.scala 130:19:@98802.4]
  assign _GEN_32 = _T_2131 ? io_app_stores_0_data_bits_wstrb : _T_2139; // @[DRAMArbiter.scala 130:19:@98810.4]
  assign _T_2213 = _T_2211 + 64'h1; // @[DRAMArbiter.scala 123:18:@98893.6]
  assign _T_2214 = _T_2211 + 64'h1; // @[DRAMArbiter.scala 123:18:@98894.6]
  assign io_app_loads_0_cmd_ready = StreamControllerLoad_io_load_cmd_ready; // @[DRAMArbiter.scala 61:17:@97837.4]
  assign io_app_loads_0_data_valid = StreamControllerLoad_io_load_data_valid; // @[DRAMArbiter.scala 61:17:@97832.4]
  assign io_app_loads_0_data_bits_rdata_0 = StreamControllerLoad_io_load_data_bits_rdata_0; // @[DRAMArbiter.scala 61:17:@97831.4]
  assign io_app_stores_0_cmd_ready = StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 68:18:@97851.4]
  assign io_app_stores_0_data_ready = StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 68:18:@97847.4]
  assign io_app_stores_0_wresp_valid = StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 68:18:@97842.4]
  assign io_app_stores_0_wresp_bits = StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 68:18:@97841.4]
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@98532.4 DRAMArbiter.scala 100:23:@98535.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@98531.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@98530.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@98528.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@98527.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@98525.4 DRAMArbiter.scala 101:25:@98537.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@98517.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@98518.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@98519.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@98520.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@98521.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@98522.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@98523.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@98524.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@98453.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@98454.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@98455.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@98456.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@98457.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@98458.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@98459.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@98460.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@98461.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@98462.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@98463.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@98464.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@98465.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@98466.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@98467.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@98468.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@98469.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@98470.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@98471.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@98472.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@98473.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@98474.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@98475.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@98476.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@98477.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@98478.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@98479.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@98480.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@98481.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@98482.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@98483.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@98484.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@98485.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@98486.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@98487.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@98488.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@98489.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@98490.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@98491.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@98492.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@98493.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@98494.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@98495.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@98496.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@98497.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@98498.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@98499.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@98500.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@98501.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@98502.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@98503.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@98504.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@98505.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@98506.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@98507.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@98508.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@98509.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@98510.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@98511.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@98512.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@98513.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@98514.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@98515.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@98516.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@98452.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@98451.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@98440.4]
  assign io_debugSignals_0 = _T_1916[31:0]; // @[DRAMArbiter.scala 111:39:@98544.4]
  assign io_debugSignals_1 = _T_1930[31:0]; // @[DRAMArbiter.scala 111:39:@98566.4]
  assign io_debugSignals_2 = _T_1944[31:0]; // @[DRAMArbiter.scala 111:39:@98574.4]
  assign io_debugSignals_3 = _T_1954[31:0]; // @[DRAMArbiter.scala 111:39:@98584.4]
  assign io_debugSignals_4 = _T_1962[31:0]; // @[DRAMArbiter.scala 111:39:@98593.4]
  assign io_debugSignals_5 = _T_1970[31:0]; // @[DRAMArbiter.scala 111:39:@98602.4]
  assign io_debugSignals_6 = _T_1978[31:0]; // @[DRAMArbiter.scala 111:39:@98611.4]
  assign io_debugSignals_7 = _T_1985[31:0]; // @[DRAMArbiter.scala 111:39:@98619.4]
  assign io_debugSignals_8 = _T_1994[31:0]; // @[DRAMArbiter.scala 111:39:@98628.4]
  assign io_debugSignals_9 = _T_2003[31:0]; // @[DRAMArbiter.scala 111:39:@98637.4]
  assign io_debugSignals_10 = _T_2021[31:0]; // @[DRAMArbiter.scala 111:39:@98656.4]
  assign io_debugSignals_11 = _T_2028[31:0]; // @[DRAMArbiter.scala 111:39:@98664.4]
  assign io_debugSignals_12 = _T_2037[31:0]; // @[DRAMArbiter.scala 111:39:@98673.4]
  assign io_debugSignals_13 = _T_2046[31:0]; // @[DRAMArbiter.scala 111:39:@98682.4]
  assign io_debugSignals_14 = _T_2064[31:0]; // @[DRAMArbiter.scala 111:39:@98701.4]
  assign io_debugSignals_15 = _T_2070[31:0]; // @[DRAMArbiter.scala 111:39:@98707.4]
  assign io_debugSignals_16 = _T_2073; // @[DRAMArbiter.scala 111:39:@98713.4]
  assign io_debugSignals_17 = _T_2076[31:0]; // @[DRAMArbiter.scala 111:39:@98719.4]
  assign io_debugSignals_18 = {{31'd0}, _T_2079}; // @[DRAMArbiter.scala 111:39:@98725.4]
  assign io_debugSignals_19 = _T_2085[31:0]; // @[DRAMArbiter.scala 111:39:@98733.4]
  assign io_debugSignals_20 = {{31'd0}, _T_2091}; // @[DRAMArbiter.scala 111:39:@98741.4]
  assign io_debugSignals_21 = _T_2097[31:0]; // @[DRAMArbiter.scala 111:39:@98749.4]
  assign io_debugSignals_22 = {{31'd0}, _T_2103}; // @[DRAMArbiter.scala 111:39:@98757.4]
  assign io_debugSignals_23 = _T_2106[31:0]; // @[DRAMArbiter.scala 111:39:@98763.4]
  assign io_debugSignals_24 = _T_2109; // @[DRAMArbiter.scala 111:39:@98769.4]
  assign io_debugSignals_25 = _T_2112; // @[DRAMArbiter.scala 111:39:@98775.4]
  assign io_debugSignals_26 = {{31'd0}, _T_2115}; // @[DRAMArbiter.scala 111:39:@98781.4]
  assign io_debugSignals_27 = _T_2121; // @[DRAMArbiter.scala 111:39:@98789.4]
  assign io_debugSignals_28 = {{31'd0}, _T_2127}; // @[DRAMArbiter.scala 111:39:@98797.4]
  assign io_debugSignals_29 = _T_2133; // @[DRAMArbiter.scala 111:39:@98805.4]
  assign io_debugSignals_30 = {{31'd0}, _T_2139}; // @[DRAMArbiter.scala 111:39:@98813.4]
  assign io_debugSignals_41 = _T_2211[31:0]; // @[DRAMArbiter.scala 111:39:@98897.4]
  assign StreamControllerLoad_clock = clock; // @[:@97829.4]
  assign StreamControllerLoad_reset = reset; // @[:@97830.4]
  assign StreamControllerLoad_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@97951.4]
  assign StreamControllerLoad_io_dram_rresp_valid = StreamArbiter_io_app_0_rresp_valid; // @[DRAMArbiter.scala 87:32:@97868.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_0 = StreamArbiter_io_app_0_rresp_bits_rdata_0; // @[DRAMArbiter.scala 87:32:@97860.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_1 = StreamArbiter_io_app_0_rresp_bits_rdata_1; // @[DRAMArbiter.scala 87:32:@97861.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_2 = StreamArbiter_io_app_0_rresp_bits_rdata_2; // @[DRAMArbiter.scala 87:32:@97862.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_3 = StreamArbiter_io_app_0_rresp_bits_rdata_3; // @[DRAMArbiter.scala 87:32:@97863.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_4 = StreamArbiter_io_app_0_rresp_bits_rdata_4; // @[DRAMArbiter.scala 87:32:@97864.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_5 = StreamArbiter_io_app_0_rresp_bits_rdata_5; // @[DRAMArbiter.scala 87:32:@97865.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_6 = StreamArbiter_io_app_0_rresp_bits_rdata_6; // @[DRAMArbiter.scala 87:32:@97866.4]
  assign StreamControllerLoad_io_dram_rresp_bits_rdata_7 = StreamArbiter_io_app_0_rresp_bits_rdata_7; // @[DRAMArbiter.scala 87:32:@97867.4]
  assign StreamControllerLoad_io_load_cmd_valid = io_app_loads_0_cmd_valid; // @[DRAMArbiter.scala 61:17:@97836.4]
  assign StreamControllerLoad_io_load_cmd_bits_addr = io_app_loads_0_cmd_bits_addr; // @[DRAMArbiter.scala 61:17:@97835.4]
  assign StreamControllerLoad_io_load_cmd_bits_size = io_app_loads_0_cmd_bits_size; // @[DRAMArbiter.scala 61:17:@97834.4]
  assign StreamControllerLoad_io_load_data_ready = io_app_loads_0_data_ready; // @[DRAMArbiter.scala 61:17:@97833.4]
  assign StreamControllerStore_clock = clock; // @[:@97839.4]
  assign StreamControllerStore_reset = reset; // @[:@97840.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_1_cmd_ready; // @[DRAMArbiter.scala 87:32:@98047.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_1_wdata_ready; // @[DRAMArbiter.scala 87:32:@98040.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_1_wresp_valid; // @[DRAMArbiter.scala 87:32:@97953.4]
  assign StreamControllerStore_io_store_cmd_valid = io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 68:18:@97850.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = io_app_stores_0_cmd_bits_addr; // @[DRAMArbiter.scala 68:18:@97849.4]
  assign StreamControllerStore_io_store_cmd_bits_size = io_app_stores_0_cmd_bits_size; // @[DRAMArbiter.scala 68:18:@97848.4]
  assign StreamControllerStore_io_store_data_valid = io_app_stores_0_data_valid; // @[DRAMArbiter.scala 68:18:@97846.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = io_app_stores_0_data_bits_wdata_0; // @[DRAMArbiter.scala 68:18:@97845.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = io_app_stores_0_data_bits_wstrb; // @[DRAMArbiter.scala 68:18:@97844.4]
  assign StreamControllerStore_io_store_wresp_ready = io_app_stores_0_wresp_ready; // @[DRAMArbiter.scala 68:18:@97843.4]
  assign StreamArbiter_clock = clock; // @[:@97853.4]
  assign StreamArbiter_reset = reset; // @[:@97854.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerLoad_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@98142.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerLoad_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@98141.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerLoad_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@98140.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h0; // @[DRAMArbiter.scala 87:22:@98138.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@98137.4]
  assign StreamArbiter_io_app_0_wdata_valid = 1'h0; // @[DRAMArbiter.scala 87:22:@98135.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = 64'h0; // @[DRAMArbiter.scala 87:22:@98127.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = 64'h0; // @[DRAMArbiter.scala 87:22:@98128.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = 64'h0; // @[DRAMArbiter.scala 87:22:@98129.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = 64'h0; // @[DRAMArbiter.scala 87:22:@98130.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = 64'h0; // @[DRAMArbiter.scala 87:22:@98131.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = 64'h0; // @[DRAMArbiter.scala 87:22:@98132.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = 64'h0; // @[DRAMArbiter.scala 87:22:@98133.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = 64'h0; // @[DRAMArbiter.scala 87:22:@98134.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = 1'h0; // @[DRAMArbiter.scala 87:22:@98063.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = 1'h0; // @[DRAMArbiter.scala 87:22:@98064.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = 1'h0; // @[DRAMArbiter.scala 87:22:@98065.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = 1'h0; // @[DRAMArbiter.scala 87:22:@98066.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = 1'h0; // @[DRAMArbiter.scala 87:22:@98067.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = 1'h0; // @[DRAMArbiter.scala 87:22:@98068.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = 1'h0; // @[DRAMArbiter.scala 87:22:@98069.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = 1'h0; // @[DRAMArbiter.scala 87:22:@98070.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = 1'h0; // @[DRAMArbiter.scala 87:22:@98071.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = 1'h0; // @[DRAMArbiter.scala 87:22:@98072.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = 1'h0; // @[DRAMArbiter.scala 87:22:@98073.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = 1'h0; // @[DRAMArbiter.scala 87:22:@98074.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = 1'h0; // @[DRAMArbiter.scala 87:22:@98075.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = 1'h0; // @[DRAMArbiter.scala 87:22:@98076.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = 1'h0; // @[DRAMArbiter.scala 87:22:@98077.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = 1'h0; // @[DRAMArbiter.scala 87:22:@98078.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = 1'h0; // @[DRAMArbiter.scala 87:22:@98079.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = 1'h0; // @[DRAMArbiter.scala 87:22:@98080.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = 1'h0; // @[DRAMArbiter.scala 87:22:@98081.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = 1'h0; // @[DRAMArbiter.scala 87:22:@98082.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = 1'h0; // @[DRAMArbiter.scala 87:22:@98083.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = 1'h0; // @[DRAMArbiter.scala 87:22:@98084.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = 1'h0; // @[DRAMArbiter.scala 87:22:@98085.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = 1'h0; // @[DRAMArbiter.scala 87:22:@98086.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = 1'h0; // @[DRAMArbiter.scala 87:22:@98087.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = 1'h0; // @[DRAMArbiter.scala 87:22:@98088.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = 1'h0; // @[DRAMArbiter.scala 87:22:@98089.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = 1'h0; // @[DRAMArbiter.scala 87:22:@98090.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = 1'h0; // @[DRAMArbiter.scala 87:22:@98091.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = 1'h0; // @[DRAMArbiter.scala 87:22:@98092.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = 1'h0; // @[DRAMArbiter.scala 87:22:@98093.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = 1'h0; // @[DRAMArbiter.scala 87:22:@98094.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = 1'h0; // @[DRAMArbiter.scala 87:22:@98095.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = 1'h0; // @[DRAMArbiter.scala 87:22:@98096.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = 1'h0; // @[DRAMArbiter.scala 87:22:@98097.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = 1'h0; // @[DRAMArbiter.scala 87:22:@98098.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = 1'h0; // @[DRAMArbiter.scala 87:22:@98099.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = 1'h0; // @[DRAMArbiter.scala 87:22:@98100.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = 1'h0; // @[DRAMArbiter.scala 87:22:@98101.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = 1'h0; // @[DRAMArbiter.scala 87:22:@98102.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = 1'h0; // @[DRAMArbiter.scala 87:22:@98103.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = 1'h0; // @[DRAMArbiter.scala 87:22:@98104.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = 1'h0; // @[DRAMArbiter.scala 87:22:@98105.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = 1'h0; // @[DRAMArbiter.scala 87:22:@98106.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = 1'h0; // @[DRAMArbiter.scala 87:22:@98107.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = 1'h0; // @[DRAMArbiter.scala 87:22:@98108.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = 1'h0; // @[DRAMArbiter.scala 87:22:@98109.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = 1'h0; // @[DRAMArbiter.scala 87:22:@98110.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = 1'h0; // @[DRAMArbiter.scala 87:22:@98111.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = 1'h0; // @[DRAMArbiter.scala 87:22:@98112.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = 1'h0; // @[DRAMArbiter.scala 87:22:@98113.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = 1'h0; // @[DRAMArbiter.scala 87:22:@98114.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = 1'h0; // @[DRAMArbiter.scala 87:22:@98115.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = 1'h0; // @[DRAMArbiter.scala 87:22:@98116.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = 1'h0; // @[DRAMArbiter.scala 87:22:@98117.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = 1'h0; // @[DRAMArbiter.scala 87:22:@98118.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = 1'h0; // @[DRAMArbiter.scala 87:22:@98119.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = 1'h0; // @[DRAMArbiter.scala 87:22:@98120.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = 1'h0; // @[DRAMArbiter.scala 87:22:@98121.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = 1'h0; // @[DRAMArbiter.scala 87:22:@98122.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = 1'h0; // @[DRAMArbiter.scala 87:22:@98123.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = 1'h0; // @[DRAMArbiter.scala 87:22:@98124.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = 1'h0; // @[DRAMArbiter.scala 87:22:@98125.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = 1'h0; // @[DRAMArbiter.scala 87:22:@98126.4]
  assign StreamArbiter_io_app_0_rresp_ready = StreamControllerLoad_io_dram_rresp_ready; // @[DRAMArbiter.scala 87:22:@98061.4]
  assign StreamArbiter_io_app_0_wresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@98050.4]
  assign StreamArbiter_io_app_1_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@98238.4]
  assign StreamArbiter_io_app_1_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@98237.4]
  assign StreamArbiter_io_app_1_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@98236.4]
  assign StreamArbiter_io_app_1_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@98234.4]
  assign StreamArbiter_io_app_1_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@98233.4]
  assign StreamArbiter_io_app_1_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@98231.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@98223.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@98224.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@98225.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@98226.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@98227.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@98228.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@98229.4]
  assign StreamArbiter_io_app_1_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@98230.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@98159.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@98160.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@98161.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@98162.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@98163.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@98164.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@98165.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@98166.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@98167.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@98168.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@98169.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@98170.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@98171.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@98172.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@98173.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@98174.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@98175.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@98176.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@98177.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@98178.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@98179.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@98180.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@98181.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@98182.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@98183.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@98184.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@98185.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@98186.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@98187.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@98188.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@98189.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@98190.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@98191.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@98192.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@98193.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@98194.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@98195.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@98196.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@98197.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@98198.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@98199.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@98200.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@98201.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@98202.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@98203.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@98204.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@98205.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@98206.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@98207.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@98208.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@98209.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@98210.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@98211.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@98212.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@98213.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@98214.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@98215.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@98216.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@98217.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@98218.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@98219.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@98220.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@98221.4]
  assign StreamArbiter_io_app_1_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@98222.4]
  assign StreamArbiter_io_app_1_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@98157.4]
  assign StreamArbiter_io_app_1_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@98146.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@98338.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@98331.4]
  assign StreamArbiter_io_dram_rresp_valid = AXICmdSplit_io_in_rresp_valid; // @[DRAMArbiter.scala 95:20:@98255.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_0 = AXICmdSplit_io_in_rresp_bits_rdata_0; // @[DRAMArbiter.scala 95:20:@98247.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_1 = AXICmdSplit_io_in_rresp_bits_rdata_1; // @[DRAMArbiter.scala 95:20:@98248.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_2 = AXICmdSplit_io_in_rresp_bits_rdata_2; // @[DRAMArbiter.scala 95:20:@98249.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_3 = AXICmdSplit_io_in_rresp_bits_rdata_3; // @[DRAMArbiter.scala 95:20:@98250.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_4 = AXICmdSplit_io_in_rresp_bits_rdata_4; // @[DRAMArbiter.scala 95:20:@98251.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_5 = AXICmdSplit_io_in_rresp_bits_rdata_5; // @[DRAMArbiter.scala 95:20:@98252.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_6 = AXICmdSplit_io_in_rresp_bits_rdata_6; // @[DRAMArbiter.scala 95:20:@98253.4]
  assign StreamArbiter_io_dram_rresp_bits_rdata_7 = AXICmdSplit_io_in_rresp_bits_rdata_7; // @[DRAMArbiter.scala 95:20:@98254.4]
  assign StreamArbiter_io_dram_rresp_bits_tag = AXICmdSplit_io_in_rresp_bits_tag; // @[DRAMArbiter.scala 95:20:@98246.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@98244.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@98243.4]
  assign AXICmdSplit_clock = clock; // @[:@98241.4]
  assign AXICmdSplit_reset = reset; // @[:@98242.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@98337.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@98336.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@98335.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@98333.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@98332.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@98330.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@98322.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@98323.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@98324.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@98325.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@98326.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@98327.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@98328.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@98329.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@98258.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@98259.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@98260.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@98261.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@98262.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@98263.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@98264.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@98265.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@98266.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@98267.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@98268.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@98269.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@98270.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@98271.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@98272.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@98273.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@98274.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@98275.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@98276.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@98277.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@98278.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@98279.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@98280.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@98281.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@98282.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@98283.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@98284.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@98285.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@98286.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@98287.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@98288.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@98289.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@98290.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@98291.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@98292.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@98293.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@98294.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@98295.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@98296.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@98297.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@98298.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@98299.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@98300.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@98301.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@98302.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@98303.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@98304.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@98305.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@98306.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@98307.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@98308.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@98309.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@98310.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@98311.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@98312.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@98313.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@98314.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@98315.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@98316.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@98317.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@98318.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@98319.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@98320.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@98321.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@98256.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@98245.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@98437.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@98430.4]
  assign AXICmdSplit_io_out_rresp_valid = AXICmdIssue_io_in_rresp_valid; // @[DRAMArbiter.scala 98:20:@98354.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_0 = AXICmdIssue_io_in_rresp_bits_rdata_0; // @[DRAMArbiter.scala 98:20:@98346.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_1 = AXICmdIssue_io_in_rresp_bits_rdata_1; // @[DRAMArbiter.scala 98:20:@98347.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_2 = AXICmdIssue_io_in_rresp_bits_rdata_2; // @[DRAMArbiter.scala 98:20:@98348.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_3 = AXICmdIssue_io_in_rresp_bits_rdata_3; // @[DRAMArbiter.scala 98:20:@98349.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_4 = AXICmdIssue_io_in_rresp_bits_rdata_4; // @[DRAMArbiter.scala 98:20:@98350.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_5 = AXICmdIssue_io_in_rresp_bits_rdata_5; // @[DRAMArbiter.scala 98:20:@98351.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_6 = AXICmdIssue_io_in_rresp_bits_rdata_6; // @[DRAMArbiter.scala 98:20:@98352.4]
  assign AXICmdSplit_io_out_rresp_bits_rdata_7 = AXICmdIssue_io_in_rresp_bits_rdata_7; // @[DRAMArbiter.scala 98:20:@98353.4]
  assign AXICmdSplit_io_out_rresp_bits_tag = AXICmdIssue_io_in_rresp_bits_tag; // @[DRAMArbiter.scala 98:20:@98345.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@98343.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@98342.4]
  assign AXICmdIssue_clock = clock; // @[:@98340.4]
  assign AXICmdIssue_reset = reset; // @[:@98341.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@98436.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@98435.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@98434.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@98432.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@98431.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@98429.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@98421.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@98422.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@98423.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@98424.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@98425.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@98426.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@98427.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@98428.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@98357.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@98358.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@98359.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@98360.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@98361.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@98362.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@98363.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@98364.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@98365.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@98366.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@98367.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@98368.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@98369.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@98370.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@98371.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@98372.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@98373.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@98374.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@98375.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@98376.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@98377.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@98378.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@98379.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@98380.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@98381.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@98382.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@98383.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@98384.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@98385.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@98386.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@98387.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@98388.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@98389.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@98390.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@98391.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@98392.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@98393.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@98394.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@98395.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@98396.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@98397.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@98398.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@98399.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@98400.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@98401.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@98402.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@98403.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@98404.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@98405.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@98406.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@98407.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@98408.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@98409.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@98410.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@98411.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@98412.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@98413.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@98414.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@98415.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@98416.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@98417.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@98418.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@98419.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@98420.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@98355.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@98344.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@98533.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@98526.4]
  assign AXICmdIssue_io_out_rresp_valid = io_dram_rresp_valid; // @[DRAMArbiter.scala 99:13:@98450.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_0 = io_dram_rresp_bits_rdata_0; // @[DRAMArbiter.scala 99:13:@98442.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_1 = io_dram_rresp_bits_rdata_1; // @[DRAMArbiter.scala 99:13:@98443.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_2 = io_dram_rresp_bits_rdata_2; // @[DRAMArbiter.scala 99:13:@98444.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_3 = io_dram_rresp_bits_rdata_3; // @[DRAMArbiter.scala 99:13:@98445.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_4 = io_dram_rresp_bits_rdata_4; // @[DRAMArbiter.scala 99:13:@98446.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_5 = io_dram_rresp_bits_rdata_5; // @[DRAMArbiter.scala 99:13:@98447.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_6 = io_dram_rresp_bits_rdata_6; // @[DRAMArbiter.scala 99:13:@98448.4]
  assign AXICmdIssue_io_out_rresp_bits_rdata_7 = io_dram_rresp_bits_rdata_7; // @[DRAMArbiter.scala 99:13:@98449.4]
  assign AXICmdIssue_io_out_rresp_bits_tag = io_dram_rresp_bits_tag; // @[DRAMArbiter.scala 99:13:@98441.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@98439.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@98438.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_1916 = _RAND_0[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  _T_1930 = _RAND_1[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  _T_1937 = _RAND_2[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{`RANDOM}};
  _T_1944 = _RAND_3[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  _T_1954 = _RAND_4[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  _T_1962 = _RAND_5[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {2{`RANDOM}};
  _T_1970 = _RAND_6[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {2{`RANDOM}};
  _T_1978 = _RAND_7[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {2{`RANDOM}};
  _T_1985 = _RAND_8[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {2{`RANDOM}};
  _T_1994 = _RAND_9[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  _T_2003 = _RAND_10[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  _T_2021 = _RAND_11[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  _T_2028 = _RAND_12[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  _T_2037 = _RAND_13[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {2{`RANDOM}};
  _T_2046 = _RAND_14[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {2{`RANDOM}};
  _T_2064 = _RAND_15[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {2{`RANDOM}};
  _T_2070 = _RAND_16[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_2073 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {2{`RANDOM}};
  _T_2076 = _RAND_18[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_2079 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  _T_2085 = _RAND_20[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_2091 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  _T_2097 = _RAND_22[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_2103 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {2{`RANDOM}};
  _T_2106 = _RAND_24[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_2109 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_2112 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_2115 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_2121 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_2127 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_2133 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_2139 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {2{`RANDOM}};
  _T_2211 = _RAND_32[63:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1916 <= 64'h0;
    end else begin
      if (io_enable) begin
        _T_1916 <= _T_1919;
      end
    end
    if (reset) begin
      _T_1930 <= 64'h0;
    end else begin
      if (_T_1927) begin
        _T_1930 <= _T_1933;
      end
    end
    if (reset) begin
      _T_1937 <= 64'h0;
    end else begin
      if (_T_1934) begin
        _T_1937 <= _T_1940;
      end
    end
    if (reset) begin
      _T_1944 <= 64'h0;
    end else begin
      if (_T_1941) begin
        _T_1944 <= _T_1947;
      end
    end
    if (reset) begin
      _T_1954 <= 64'h0;
    end else begin
      if (_T_1951) begin
        _T_1954 <= _T_1957;
      end
    end
    if (reset) begin
      _T_1962 <= 64'h0;
    end else begin
      if (_T_1959) begin
        _T_1962 <= _T_1965;
      end
    end
    if (reset) begin
      _T_1970 <= 64'h0;
    end else begin
      if (_T_1967) begin
        _T_1970 <= _T_1973;
      end
    end
    if (reset) begin
      _T_1978 <= 64'h0;
    end else begin
      if (_T_1975) begin
        _T_1978 <= _T_1981;
      end
    end
    if (reset) begin
      _T_1985 <= 64'h0;
    end else begin
      if (_T_1920) begin
        _T_1985 <= _T_1988;
      end
    end
    if (reset) begin
      _T_1994 <= 64'h0;
    end else begin
      if (_T_1991) begin
        _T_1994 <= _T_1997;
      end
    end
    if (reset) begin
      _T_2003 <= 64'h0;
    end else begin
      if (_T_2000) begin
        _T_2003 <= _T_2006;
      end
    end
    if (reset) begin
      _T_2021 <= 64'h0;
    end else begin
      if (_T_2018) begin
        _T_2021 <= _T_2024;
      end
    end
    if (reset) begin
      _T_2028 <= 64'h0;
    end else begin
      if (_T_2025) begin
        _T_2028 <= _T_2031;
      end
    end
    if (reset) begin
      _T_2037 <= 64'h0;
    end else begin
      if (_T_2034) begin
        _T_2037 <= _T_2040;
      end
    end
    if (reset) begin
      _T_2046 <= 64'h0;
    end else begin
      if (_T_2043) begin
        _T_2046 <= _T_2049;
      end
    end
    if (reset) begin
      _T_2064 <= 64'h0;
    end else begin
      if (_T_2061) begin
        _T_2064 <= _T_2067;
      end
    end
    if (reset) begin
      _T_2070 <= io_dram_cmd_bits_addr;
    end else begin
      if (_T_2068) begin
        _T_2070 <= io_dram_cmd_bits_addr;
      end
    end
    if (reset) begin
      _T_2073 <= io_dram_cmd_bits_size;
    end else begin
      if (_T_2068) begin
        _T_2073 <= io_dram_cmd_bits_size;
      end
    end
    if (reset) begin
      _T_2076 <= io_dram_wdata_bits_wdata_0;
    end else begin
      if (_T_1927) begin
        _T_2076 <= io_dram_wdata_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_2079 <= io_dram_wdata_bits_wstrb_0;
    end else begin
      if (_T_1927) begin
        _T_2079 <= io_dram_wdata_bits_wstrb_0;
      end
    end
    if (reset) begin
      _T_2085 <= io_dram_wdata_bits_wdata_0;
    end else begin
      if (_T_2083) begin
        _T_2085 <= io_dram_wdata_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_2091 <= io_dram_wdata_bits_wstrb_0;
    end else begin
      if (_T_2083) begin
        _T_2091 <= io_dram_wdata_bits_wstrb_0;
      end
    end
    if (reset) begin
      _T_2097 <= io_dram_wdata_bits_wdata_0;
    end else begin
      if (_T_2095) begin
        _T_2097 <= io_dram_wdata_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_2103 <= io_dram_wdata_bits_wstrb_0;
    end else begin
      if (_T_2095) begin
        _T_2103 <= io_dram_wdata_bits_wstrb_0;
      end
    end
    if (reset) begin
      _T_2106 <= io_app_stores_0_cmd_bits_addr;
    end else begin
      if (_T_2104) begin
        _T_2106 <= io_app_stores_0_cmd_bits_addr;
      end
    end
    if (reset) begin
      _T_2109 <= io_app_stores_0_cmd_bits_size;
    end else begin
      if (_T_2104) begin
        _T_2109 <= io_app_stores_0_cmd_bits_size;
      end
    end
    if (reset) begin
      _T_2112 <= io_app_stores_0_data_bits_wdata_0;
    end else begin
      if (_T_1934) begin
        _T_2112 <= io_app_stores_0_data_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_2115 <= io_app_stores_0_data_bits_wstrb;
    end else begin
      if (_T_1934) begin
        _T_2115 <= io_app_stores_0_data_bits_wstrb;
      end
    end
    if (reset) begin
      _T_2121 <= io_app_stores_0_data_bits_wdata_0;
    end else begin
      if (_T_2119) begin
        _T_2121 <= io_app_stores_0_data_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_2127 <= io_app_stores_0_data_bits_wstrb;
    end else begin
      if (_T_2119) begin
        _T_2127 <= io_app_stores_0_data_bits_wstrb;
      end
    end
    if (reset) begin
      _T_2133 <= io_app_stores_0_data_bits_wdata_0;
    end else begin
      if (_T_2131) begin
        _T_2133 <= io_app_stores_0_data_bits_wdata_0;
      end
    end
    if (reset) begin
      _T_2139 <= io_app_stores_0_data_bits_wstrb;
    end else begin
      if (_T_2131) begin
        _T_2139 <= io_app_stores_0_data_bits_wstrb;
      end
    end
    if (reset) begin
      _T_2211 <= 64'h0;
    end else begin
      _T_2211 <= _T_2214;
    end
  end
endmodule
module DRAMHeap( // @[:@120779.2]
  input         io_accel_0_req_valid, // @[:@120782.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@120782.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@120782.4]
  output        io_accel_0_resp_valid, // @[:@120782.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@120782.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@120782.4]
  output        io_host_0_req_valid, // @[:@120782.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@120782.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@120782.4]
  input         io_host_0_resp_valid, // @[:@120782.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@120782.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@120782.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@120789.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@120791.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@120790.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@120786.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@120785.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@120784.4]
endmodule
module FringeFF( // @[:@120825.2]
  input         clock, // @[:@120826.4]
  input         reset, // @[:@120827.4]
  input  [63:0] io_in, // @[:@120828.4]
  input         io_reset, // @[:@120828.4]
  output [63:0] io_out, // @[:@120828.4]
  input         io_enable // @[:@120828.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@120831.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@120831.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@120831.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@120831.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@120831.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@120836.4 package.scala 96:25:@120837.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@120842.6]
  RetimeWrapper_37 RetimeWrapper ( // @[package.scala 93:22:@120831.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@120836.4 package.scala 96:25:@120837.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@120842.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@120848.4]
  assign RetimeWrapper_clock = clock; // @[:@120832.4]
  assign RetimeWrapper_reset = reset; // @[:@120833.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@120835.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@120834.4]
endmodule
module MuxN_4( // @[:@149464.2]
  input  [63:0] io_ins_0, // @[:@149467.4]
  input  [63:0] io_ins_1, // @[:@149467.4]
  input  [63:0] io_ins_2, // @[:@149467.4]
  input  [63:0] io_ins_3, // @[:@149467.4]
  input  [63:0] io_ins_4, // @[:@149467.4]
  input  [63:0] io_ins_5, // @[:@149467.4]
  input  [63:0] io_ins_6, // @[:@149467.4]
  input  [63:0] io_ins_7, // @[:@149467.4]
  input  [63:0] io_ins_8, // @[:@149467.4]
  input  [63:0] io_ins_9, // @[:@149467.4]
  input  [63:0] io_ins_10, // @[:@149467.4]
  input  [63:0] io_ins_11, // @[:@149467.4]
  input  [63:0] io_ins_12, // @[:@149467.4]
  input  [63:0] io_ins_13, // @[:@149467.4]
  input  [63:0] io_ins_14, // @[:@149467.4]
  input  [63:0] io_ins_15, // @[:@149467.4]
  input  [63:0] io_ins_16, // @[:@149467.4]
  input  [63:0] io_ins_17, // @[:@149467.4]
  input  [63:0] io_ins_18, // @[:@149467.4]
  input  [63:0] io_ins_19, // @[:@149467.4]
  input  [63:0] io_ins_20, // @[:@149467.4]
  input  [63:0] io_ins_21, // @[:@149467.4]
  input  [63:0] io_ins_22, // @[:@149467.4]
  input  [63:0] io_ins_23, // @[:@149467.4]
  input  [63:0] io_ins_24, // @[:@149467.4]
  input  [63:0] io_ins_25, // @[:@149467.4]
  input  [63:0] io_ins_26, // @[:@149467.4]
  input  [63:0] io_ins_27, // @[:@149467.4]
  input  [63:0] io_ins_28, // @[:@149467.4]
  input  [63:0] io_ins_29, // @[:@149467.4]
  input  [63:0] io_ins_30, // @[:@149467.4]
  input  [63:0] io_ins_31, // @[:@149467.4]
  input  [63:0] io_ins_32, // @[:@149467.4]
  input  [63:0] io_ins_33, // @[:@149467.4]
  input  [63:0] io_ins_34, // @[:@149467.4]
  input  [63:0] io_ins_35, // @[:@149467.4]
  input  [63:0] io_ins_36, // @[:@149467.4]
  input  [63:0] io_ins_37, // @[:@149467.4]
  input  [63:0] io_ins_38, // @[:@149467.4]
  input  [63:0] io_ins_39, // @[:@149467.4]
  input  [63:0] io_ins_40, // @[:@149467.4]
  input  [63:0] io_ins_41, // @[:@149467.4]
  input  [63:0] io_ins_42, // @[:@149467.4]
  input  [63:0] io_ins_43, // @[:@149467.4]
  input  [63:0] io_ins_44, // @[:@149467.4]
  input  [63:0] io_ins_45, // @[:@149467.4]
  input  [63:0] io_ins_46, // @[:@149467.4]
  input  [63:0] io_ins_47, // @[:@149467.4]
  input  [63:0] io_ins_48, // @[:@149467.4]
  input  [63:0] io_ins_49, // @[:@149467.4]
  input  [63:0] io_ins_50, // @[:@149467.4]
  input  [63:0] io_ins_51, // @[:@149467.4]
  input  [63:0] io_ins_52, // @[:@149467.4]
  input  [63:0] io_ins_53, // @[:@149467.4]
  input  [63:0] io_ins_54, // @[:@149467.4]
  input  [63:0] io_ins_55, // @[:@149467.4]
  input  [63:0] io_ins_56, // @[:@149467.4]
  input  [63:0] io_ins_57, // @[:@149467.4]
  input  [63:0] io_ins_58, // @[:@149467.4]
  input  [63:0] io_ins_59, // @[:@149467.4]
  input  [63:0] io_ins_60, // @[:@149467.4]
  input  [63:0] io_ins_61, // @[:@149467.4]
  input  [63:0] io_ins_62, // @[:@149467.4]
  input  [63:0] io_ins_63, // @[:@149467.4]
  input  [63:0] io_ins_64, // @[:@149467.4]
  input  [63:0] io_ins_65, // @[:@149467.4]
  input  [63:0] io_ins_66, // @[:@149467.4]
  input  [63:0] io_ins_67, // @[:@149467.4]
  input  [63:0] io_ins_68, // @[:@149467.4]
  input  [63:0] io_ins_69, // @[:@149467.4]
  input  [63:0] io_ins_70, // @[:@149467.4]
  input  [63:0] io_ins_71, // @[:@149467.4]
  input  [63:0] io_ins_72, // @[:@149467.4]
  input  [63:0] io_ins_73, // @[:@149467.4]
  input  [63:0] io_ins_74, // @[:@149467.4]
  input  [63:0] io_ins_75, // @[:@149467.4]
  input  [63:0] io_ins_76, // @[:@149467.4]
  input  [63:0] io_ins_77, // @[:@149467.4]
  input  [63:0] io_ins_78, // @[:@149467.4]
  input  [63:0] io_ins_79, // @[:@149467.4]
  input  [63:0] io_ins_80, // @[:@149467.4]
  input  [63:0] io_ins_81, // @[:@149467.4]
  input  [63:0] io_ins_82, // @[:@149467.4]
  input  [63:0] io_ins_83, // @[:@149467.4]
  input  [63:0] io_ins_84, // @[:@149467.4]
  input  [63:0] io_ins_85, // @[:@149467.4]
  input  [63:0] io_ins_86, // @[:@149467.4]
  input  [63:0] io_ins_87, // @[:@149467.4]
  input  [63:0] io_ins_88, // @[:@149467.4]
  input  [63:0] io_ins_89, // @[:@149467.4]
  input  [63:0] io_ins_90, // @[:@149467.4]
  input  [63:0] io_ins_91, // @[:@149467.4]
  input  [63:0] io_ins_92, // @[:@149467.4]
  input  [63:0] io_ins_93, // @[:@149467.4]
  input  [63:0] io_ins_94, // @[:@149467.4]
  input  [63:0] io_ins_95, // @[:@149467.4]
  input  [63:0] io_ins_96, // @[:@149467.4]
  input  [63:0] io_ins_97, // @[:@149467.4]
  input  [63:0] io_ins_98, // @[:@149467.4]
  input  [63:0] io_ins_99, // @[:@149467.4]
  input  [63:0] io_ins_100, // @[:@149467.4]
  input  [63:0] io_ins_101, // @[:@149467.4]
  input  [63:0] io_ins_102, // @[:@149467.4]
  input  [63:0] io_ins_103, // @[:@149467.4]
  input  [63:0] io_ins_104, // @[:@149467.4]
  input  [63:0] io_ins_105, // @[:@149467.4]
  input  [63:0] io_ins_106, // @[:@149467.4]
  input  [63:0] io_ins_107, // @[:@149467.4]
  input  [63:0] io_ins_108, // @[:@149467.4]
  input  [63:0] io_ins_109, // @[:@149467.4]
  input  [63:0] io_ins_110, // @[:@149467.4]
  input  [63:0] io_ins_111, // @[:@149467.4]
  input  [63:0] io_ins_112, // @[:@149467.4]
  input  [63:0] io_ins_113, // @[:@149467.4]
  input  [63:0] io_ins_114, // @[:@149467.4]
  input  [63:0] io_ins_115, // @[:@149467.4]
  input  [63:0] io_ins_116, // @[:@149467.4]
  input  [63:0] io_ins_117, // @[:@149467.4]
  input  [63:0] io_ins_118, // @[:@149467.4]
  input  [63:0] io_ins_119, // @[:@149467.4]
  input  [63:0] io_ins_120, // @[:@149467.4]
  input  [63:0] io_ins_121, // @[:@149467.4]
  input  [63:0] io_ins_122, // @[:@149467.4]
  input  [63:0] io_ins_123, // @[:@149467.4]
  input  [63:0] io_ins_124, // @[:@149467.4]
  input  [63:0] io_ins_125, // @[:@149467.4]
  input  [63:0] io_ins_126, // @[:@149467.4]
  input  [63:0] io_ins_127, // @[:@149467.4]
  input  [63:0] io_ins_128, // @[:@149467.4]
  input  [63:0] io_ins_129, // @[:@149467.4]
  input  [63:0] io_ins_130, // @[:@149467.4]
  input  [63:0] io_ins_131, // @[:@149467.4]
  input  [63:0] io_ins_132, // @[:@149467.4]
  input  [63:0] io_ins_133, // @[:@149467.4]
  input  [63:0] io_ins_134, // @[:@149467.4]
  input  [63:0] io_ins_135, // @[:@149467.4]
  input  [63:0] io_ins_136, // @[:@149467.4]
  input  [63:0] io_ins_137, // @[:@149467.4]
  input  [63:0] io_ins_138, // @[:@149467.4]
  input  [63:0] io_ins_139, // @[:@149467.4]
  input  [63:0] io_ins_140, // @[:@149467.4]
  input  [63:0] io_ins_141, // @[:@149467.4]
  input  [63:0] io_ins_142, // @[:@149467.4]
  input  [63:0] io_ins_143, // @[:@149467.4]
  input  [63:0] io_ins_144, // @[:@149467.4]
  input  [63:0] io_ins_145, // @[:@149467.4]
  input  [63:0] io_ins_146, // @[:@149467.4]
  input  [63:0] io_ins_147, // @[:@149467.4]
  input  [63:0] io_ins_148, // @[:@149467.4]
  input  [63:0] io_ins_149, // @[:@149467.4]
  input  [63:0] io_ins_150, // @[:@149467.4]
  input  [63:0] io_ins_151, // @[:@149467.4]
  input  [63:0] io_ins_152, // @[:@149467.4]
  input  [63:0] io_ins_153, // @[:@149467.4]
  input  [63:0] io_ins_154, // @[:@149467.4]
  input  [63:0] io_ins_155, // @[:@149467.4]
  input  [63:0] io_ins_156, // @[:@149467.4]
  input  [63:0] io_ins_157, // @[:@149467.4]
  input  [63:0] io_ins_158, // @[:@149467.4]
  input  [63:0] io_ins_159, // @[:@149467.4]
  input  [63:0] io_ins_160, // @[:@149467.4]
  input  [63:0] io_ins_161, // @[:@149467.4]
  input  [63:0] io_ins_162, // @[:@149467.4]
  input  [63:0] io_ins_163, // @[:@149467.4]
  input  [63:0] io_ins_164, // @[:@149467.4]
  input  [63:0] io_ins_165, // @[:@149467.4]
  input  [63:0] io_ins_166, // @[:@149467.4]
  input  [63:0] io_ins_167, // @[:@149467.4]
  input  [63:0] io_ins_168, // @[:@149467.4]
  input  [63:0] io_ins_169, // @[:@149467.4]
  input  [63:0] io_ins_170, // @[:@149467.4]
  input  [63:0] io_ins_171, // @[:@149467.4]
  input  [63:0] io_ins_172, // @[:@149467.4]
  input  [63:0] io_ins_173, // @[:@149467.4]
  input  [63:0] io_ins_174, // @[:@149467.4]
  input  [63:0] io_ins_175, // @[:@149467.4]
  input  [63:0] io_ins_176, // @[:@149467.4]
  input  [63:0] io_ins_177, // @[:@149467.4]
  input  [63:0] io_ins_178, // @[:@149467.4]
  input  [63:0] io_ins_179, // @[:@149467.4]
  input  [63:0] io_ins_180, // @[:@149467.4]
  input  [63:0] io_ins_181, // @[:@149467.4]
  input  [63:0] io_ins_182, // @[:@149467.4]
  input  [63:0] io_ins_183, // @[:@149467.4]
  input  [63:0] io_ins_184, // @[:@149467.4]
  input  [63:0] io_ins_185, // @[:@149467.4]
  input  [63:0] io_ins_186, // @[:@149467.4]
  input  [63:0] io_ins_187, // @[:@149467.4]
  input  [63:0] io_ins_188, // @[:@149467.4]
  input  [63:0] io_ins_189, // @[:@149467.4]
  input  [63:0] io_ins_190, // @[:@149467.4]
  input  [63:0] io_ins_191, // @[:@149467.4]
  input  [63:0] io_ins_192, // @[:@149467.4]
  input  [63:0] io_ins_193, // @[:@149467.4]
  input  [63:0] io_ins_194, // @[:@149467.4]
  input  [63:0] io_ins_195, // @[:@149467.4]
  input  [63:0] io_ins_196, // @[:@149467.4]
  input  [63:0] io_ins_197, // @[:@149467.4]
  input  [63:0] io_ins_198, // @[:@149467.4]
  input  [63:0] io_ins_199, // @[:@149467.4]
  input  [63:0] io_ins_200, // @[:@149467.4]
  input  [63:0] io_ins_201, // @[:@149467.4]
  input  [63:0] io_ins_202, // @[:@149467.4]
  input  [63:0] io_ins_203, // @[:@149467.4]
  input  [63:0] io_ins_204, // @[:@149467.4]
  input  [63:0] io_ins_205, // @[:@149467.4]
  input  [63:0] io_ins_206, // @[:@149467.4]
  input  [63:0] io_ins_207, // @[:@149467.4]
  input  [63:0] io_ins_208, // @[:@149467.4]
  input  [63:0] io_ins_209, // @[:@149467.4]
  input  [63:0] io_ins_210, // @[:@149467.4]
  input  [63:0] io_ins_211, // @[:@149467.4]
  input  [63:0] io_ins_212, // @[:@149467.4]
  input  [63:0] io_ins_213, // @[:@149467.4]
  input  [63:0] io_ins_214, // @[:@149467.4]
  input  [63:0] io_ins_215, // @[:@149467.4]
  input  [63:0] io_ins_216, // @[:@149467.4]
  input  [63:0] io_ins_217, // @[:@149467.4]
  input  [63:0] io_ins_218, // @[:@149467.4]
  input  [63:0] io_ins_219, // @[:@149467.4]
  input  [63:0] io_ins_220, // @[:@149467.4]
  input  [63:0] io_ins_221, // @[:@149467.4]
  input  [63:0] io_ins_222, // @[:@149467.4]
  input  [63:0] io_ins_223, // @[:@149467.4]
  input  [63:0] io_ins_224, // @[:@149467.4]
  input  [63:0] io_ins_225, // @[:@149467.4]
  input  [63:0] io_ins_226, // @[:@149467.4]
  input  [63:0] io_ins_227, // @[:@149467.4]
  input  [63:0] io_ins_228, // @[:@149467.4]
  input  [63:0] io_ins_229, // @[:@149467.4]
  input  [63:0] io_ins_230, // @[:@149467.4]
  input  [63:0] io_ins_231, // @[:@149467.4]
  input  [63:0] io_ins_232, // @[:@149467.4]
  input  [63:0] io_ins_233, // @[:@149467.4]
  input  [63:0] io_ins_234, // @[:@149467.4]
  input  [63:0] io_ins_235, // @[:@149467.4]
  input  [63:0] io_ins_236, // @[:@149467.4]
  input  [63:0] io_ins_237, // @[:@149467.4]
  input  [63:0] io_ins_238, // @[:@149467.4]
  input  [63:0] io_ins_239, // @[:@149467.4]
  input  [63:0] io_ins_240, // @[:@149467.4]
  input  [63:0] io_ins_241, // @[:@149467.4]
  input  [63:0] io_ins_242, // @[:@149467.4]
  input  [63:0] io_ins_243, // @[:@149467.4]
  input  [63:0] io_ins_244, // @[:@149467.4]
  input  [63:0] io_ins_245, // @[:@149467.4]
  input  [63:0] io_ins_246, // @[:@149467.4]
  input  [63:0] io_ins_247, // @[:@149467.4]
  input  [63:0] io_ins_248, // @[:@149467.4]
  input  [63:0] io_ins_249, // @[:@149467.4]
  input  [63:0] io_ins_250, // @[:@149467.4]
  input  [63:0] io_ins_251, // @[:@149467.4]
  input  [63:0] io_ins_252, // @[:@149467.4]
  input  [63:0] io_ins_253, // @[:@149467.4]
  input  [63:0] io_ins_254, // @[:@149467.4]
  input  [63:0] io_ins_255, // @[:@149467.4]
  input  [63:0] io_ins_256, // @[:@149467.4]
  input  [63:0] io_ins_257, // @[:@149467.4]
  input  [63:0] io_ins_258, // @[:@149467.4]
  input  [63:0] io_ins_259, // @[:@149467.4]
  input  [63:0] io_ins_260, // @[:@149467.4]
  input  [63:0] io_ins_261, // @[:@149467.4]
  input  [63:0] io_ins_262, // @[:@149467.4]
  input  [63:0] io_ins_263, // @[:@149467.4]
  input  [63:0] io_ins_264, // @[:@149467.4]
  input  [63:0] io_ins_265, // @[:@149467.4]
  input  [63:0] io_ins_266, // @[:@149467.4]
  input  [63:0] io_ins_267, // @[:@149467.4]
  input  [63:0] io_ins_268, // @[:@149467.4]
  input  [63:0] io_ins_269, // @[:@149467.4]
  input  [63:0] io_ins_270, // @[:@149467.4]
  input  [63:0] io_ins_271, // @[:@149467.4]
  input  [63:0] io_ins_272, // @[:@149467.4]
  input  [63:0] io_ins_273, // @[:@149467.4]
  input  [63:0] io_ins_274, // @[:@149467.4]
  input  [63:0] io_ins_275, // @[:@149467.4]
  input  [63:0] io_ins_276, // @[:@149467.4]
  input  [63:0] io_ins_277, // @[:@149467.4]
  input  [63:0] io_ins_278, // @[:@149467.4]
  input  [63:0] io_ins_279, // @[:@149467.4]
  input  [63:0] io_ins_280, // @[:@149467.4]
  input  [63:0] io_ins_281, // @[:@149467.4]
  input  [63:0] io_ins_282, // @[:@149467.4]
  input  [63:0] io_ins_283, // @[:@149467.4]
  input  [63:0] io_ins_284, // @[:@149467.4]
  input  [63:0] io_ins_285, // @[:@149467.4]
  input  [63:0] io_ins_286, // @[:@149467.4]
  input  [63:0] io_ins_287, // @[:@149467.4]
  input  [63:0] io_ins_288, // @[:@149467.4]
  input  [63:0] io_ins_289, // @[:@149467.4]
  input  [63:0] io_ins_290, // @[:@149467.4]
  input  [63:0] io_ins_291, // @[:@149467.4]
  input  [63:0] io_ins_292, // @[:@149467.4]
  input  [63:0] io_ins_293, // @[:@149467.4]
  input  [63:0] io_ins_294, // @[:@149467.4]
  input  [63:0] io_ins_295, // @[:@149467.4]
  input  [63:0] io_ins_296, // @[:@149467.4]
  input  [63:0] io_ins_297, // @[:@149467.4]
  input  [63:0] io_ins_298, // @[:@149467.4]
  input  [63:0] io_ins_299, // @[:@149467.4]
  input  [63:0] io_ins_300, // @[:@149467.4]
  input  [63:0] io_ins_301, // @[:@149467.4]
  input  [63:0] io_ins_302, // @[:@149467.4]
  input  [63:0] io_ins_303, // @[:@149467.4]
  input  [63:0] io_ins_304, // @[:@149467.4]
  input  [63:0] io_ins_305, // @[:@149467.4]
  input  [63:0] io_ins_306, // @[:@149467.4]
  input  [63:0] io_ins_307, // @[:@149467.4]
  input  [63:0] io_ins_308, // @[:@149467.4]
  input  [63:0] io_ins_309, // @[:@149467.4]
  input  [63:0] io_ins_310, // @[:@149467.4]
  input  [63:0] io_ins_311, // @[:@149467.4]
  input  [63:0] io_ins_312, // @[:@149467.4]
  input  [63:0] io_ins_313, // @[:@149467.4]
  input  [63:0] io_ins_314, // @[:@149467.4]
  input  [63:0] io_ins_315, // @[:@149467.4]
  input  [63:0] io_ins_316, // @[:@149467.4]
  input  [63:0] io_ins_317, // @[:@149467.4]
  input  [63:0] io_ins_318, // @[:@149467.4]
  input  [63:0] io_ins_319, // @[:@149467.4]
  input  [63:0] io_ins_320, // @[:@149467.4]
  input  [63:0] io_ins_321, // @[:@149467.4]
  input  [63:0] io_ins_322, // @[:@149467.4]
  input  [63:0] io_ins_323, // @[:@149467.4]
  input  [63:0] io_ins_324, // @[:@149467.4]
  input  [63:0] io_ins_325, // @[:@149467.4]
  input  [63:0] io_ins_326, // @[:@149467.4]
  input  [63:0] io_ins_327, // @[:@149467.4]
  input  [63:0] io_ins_328, // @[:@149467.4]
  input  [63:0] io_ins_329, // @[:@149467.4]
  input  [63:0] io_ins_330, // @[:@149467.4]
  input  [63:0] io_ins_331, // @[:@149467.4]
  input  [63:0] io_ins_332, // @[:@149467.4]
  input  [63:0] io_ins_333, // @[:@149467.4]
  input  [63:0] io_ins_334, // @[:@149467.4]
  input  [63:0] io_ins_335, // @[:@149467.4]
  input  [63:0] io_ins_336, // @[:@149467.4]
  input  [63:0] io_ins_337, // @[:@149467.4]
  input  [63:0] io_ins_338, // @[:@149467.4]
  input  [63:0] io_ins_339, // @[:@149467.4]
  input  [63:0] io_ins_340, // @[:@149467.4]
  input  [63:0] io_ins_341, // @[:@149467.4]
  input  [63:0] io_ins_342, // @[:@149467.4]
  input  [63:0] io_ins_343, // @[:@149467.4]
  input  [63:0] io_ins_344, // @[:@149467.4]
  input  [63:0] io_ins_345, // @[:@149467.4]
  input  [63:0] io_ins_346, // @[:@149467.4]
  input  [63:0] io_ins_347, // @[:@149467.4]
  input  [63:0] io_ins_348, // @[:@149467.4]
  input  [63:0] io_ins_349, // @[:@149467.4]
  input  [63:0] io_ins_350, // @[:@149467.4]
  input  [63:0] io_ins_351, // @[:@149467.4]
  input  [63:0] io_ins_352, // @[:@149467.4]
  input  [63:0] io_ins_353, // @[:@149467.4]
  input  [63:0] io_ins_354, // @[:@149467.4]
  input  [63:0] io_ins_355, // @[:@149467.4]
  input  [63:0] io_ins_356, // @[:@149467.4]
  input  [63:0] io_ins_357, // @[:@149467.4]
  input  [63:0] io_ins_358, // @[:@149467.4]
  input  [63:0] io_ins_359, // @[:@149467.4]
  input  [63:0] io_ins_360, // @[:@149467.4]
  input  [63:0] io_ins_361, // @[:@149467.4]
  input  [63:0] io_ins_362, // @[:@149467.4]
  input  [63:0] io_ins_363, // @[:@149467.4]
  input  [63:0] io_ins_364, // @[:@149467.4]
  input  [63:0] io_ins_365, // @[:@149467.4]
  input  [63:0] io_ins_366, // @[:@149467.4]
  input  [63:0] io_ins_367, // @[:@149467.4]
  input  [63:0] io_ins_368, // @[:@149467.4]
  input  [63:0] io_ins_369, // @[:@149467.4]
  input  [63:0] io_ins_370, // @[:@149467.4]
  input  [63:0] io_ins_371, // @[:@149467.4]
  input  [63:0] io_ins_372, // @[:@149467.4]
  input  [63:0] io_ins_373, // @[:@149467.4]
  input  [63:0] io_ins_374, // @[:@149467.4]
  input  [63:0] io_ins_375, // @[:@149467.4]
  input  [63:0] io_ins_376, // @[:@149467.4]
  input  [63:0] io_ins_377, // @[:@149467.4]
  input  [63:0] io_ins_378, // @[:@149467.4]
  input  [63:0] io_ins_379, // @[:@149467.4]
  input  [63:0] io_ins_380, // @[:@149467.4]
  input  [63:0] io_ins_381, // @[:@149467.4]
  input  [63:0] io_ins_382, // @[:@149467.4]
  input  [63:0] io_ins_383, // @[:@149467.4]
  input  [63:0] io_ins_384, // @[:@149467.4]
  input  [63:0] io_ins_385, // @[:@149467.4]
  input  [63:0] io_ins_386, // @[:@149467.4]
  input  [63:0] io_ins_387, // @[:@149467.4]
  input  [63:0] io_ins_388, // @[:@149467.4]
  input  [63:0] io_ins_389, // @[:@149467.4]
  input  [63:0] io_ins_390, // @[:@149467.4]
  input  [63:0] io_ins_391, // @[:@149467.4]
  input  [63:0] io_ins_392, // @[:@149467.4]
  input  [63:0] io_ins_393, // @[:@149467.4]
  input  [63:0] io_ins_394, // @[:@149467.4]
  input  [63:0] io_ins_395, // @[:@149467.4]
  input  [63:0] io_ins_396, // @[:@149467.4]
  input  [63:0] io_ins_397, // @[:@149467.4]
  input  [63:0] io_ins_398, // @[:@149467.4]
  input  [63:0] io_ins_399, // @[:@149467.4]
  input  [63:0] io_ins_400, // @[:@149467.4]
  input  [63:0] io_ins_401, // @[:@149467.4]
  input  [63:0] io_ins_402, // @[:@149467.4]
  input  [63:0] io_ins_403, // @[:@149467.4]
  input  [63:0] io_ins_404, // @[:@149467.4]
  input  [63:0] io_ins_405, // @[:@149467.4]
  input  [63:0] io_ins_406, // @[:@149467.4]
  input  [63:0] io_ins_407, // @[:@149467.4]
  input  [63:0] io_ins_408, // @[:@149467.4]
  input  [63:0] io_ins_409, // @[:@149467.4]
  input  [63:0] io_ins_410, // @[:@149467.4]
  input  [63:0] io_ins_411, // @[:@149467.4]
  input  [63:0] io_ins_412, // @[:@149467.4]
  input  [63:0] io_ins_413, // @[:@149467.4]
  input  [63:0] io_ins_414, // @[:@149467.4]
  input  [63:0] io_ins_415, // @[:@149467.4]
  input  [63:0] io_ins_416, // @[:@149467.4]
  input  [63:0] io_ins_417, // @[:@149467.4]
  input  [63:0] io_ins_418, // @[:@149467.4]
  input  [63:0] io_ins_419, // @[:@149467.4]
  input  [63:0] io_ins_420, // @[:@149467.4]
  input  [63:0] io_ins_421, // @[:@149467.4]
  input  [63:0] io_ins_422, // @[:@149467.4]
  input  [63:0] io_ins_423, // @[:@149467.4]
  input  [63:0] io_ins_424, // @[:@149467.4]
  input  [63:0] io_ins_425, // @[:@149467.4]
  input  [63:0] io_ins_426, // @[:@149467.4]
  input  [63:0] io_ins_427, // @[:@149467.4]
  input  [63:0] io_ins_428, // @[:@149467.4]
  input  [63:0] io_ins_429, // @[:@149467.4]
  input  [63:0] io_ins_430, // @[:@149467.4]
  input  [63:0] io_ins_431, // @[:@149467.4]
  input  [63:0] io_ins_432, // @[:@149467.4]
  input  [63:0] io_ins_433, // @[:@149467.4]
  input  [63:0] io_ins_434, // @[:@149467.4]
  input  [63:0] io_ins_435, // @[:@149467.4]
  input  [63:0] io_ins_436, // @[:@149467.4]
  input  [63:0] io_ins_437, // @[:@149467.4]
  input  [63:0] io_ins_438, // @[:@149467.4]
  input  [63:0] io_ins_439, // @[:@149467.4]
  input  [63:0] io_ins_440, // @[:@149467.4]
  input  [63:0] io_ins_441, // @[:@149467.4]
  input  [63:0] io_ins_442, // @[:@149467.4]
  input  [63:0] io_ins_443, // @[:@149467.4]
  input  [63:0] io_ins_444, // @[:@149467.4]
  input  [63:0] io_ins_445, // @[:@149467.4]
  input  [63:0] io_ins_446, // @[:@149467.4]
  input  [63:0] io_ins_447, // @[:@149467.4]
  input  [63:0] io_ins_448, // @[:@149467.4]
  input  [63:0] io_ins_449, // @[:@149467.4]
  input  [63:0] io_ins_450, // @[:@149467.4]
  input  [63:0] io_ins_451, // @[:@149467.4]
  input  [63:0] io_ins_452, // @[:@149467.4]
  input  [63:0] io_ins_453, // @[:@149467.4]
  input  [63:0] io_ins_454, // @[:@149467.4]
  input  [63:0] io_ins_455, // @[:@149467.4]
  input  [63:0] io_ins_456, // @[:@149467.4]
  input  [63:0] io_ins_457, // @[:@149467.4]
  input  [63:0] io_ins_458, // @[:@149467.4]
  input  [63:0] io_ins_459, // @[:@149467.4]
  input  [63:0] io_ins_460, // @[:@149467.4]
  input  [63:0] io_ins_461, // @[:@149467.4]
  input  [63:0] io_ins_462, // @[:@149467.4]
  input  [63:0] io_ins_463, // @[:@149467.4]
  input  [63:0] io_ins_464, // @[:@149467.4]
  input  [63:0] io_ins_465, // @[:@149467.4]
  input  [63:0] io_ins_466, // @[:@149467.4]
  input  [63:0] io_ins_467, // @[:@149467.4]
  input  [63:0] io_ins_468, // @[:@149467.4]
  input  [63:0] io_ins_469, // @[:@149467.4]
  input  [63:0] io_ins_470, // @[:@149467.4]
  input  [63:0] io_ins_471, // @[:@149467.4]
  input  [63:0] io_ins_472, // @[:@149467.4]
  input  [63:0] io_ins_473, // @[:@149467.4]
  input  [63:0] io_ins_474, // @[:@149467.4]
  input  [63:0] io_ins_475, // @[:@149467.4]
  input  [63:0] io_ins_476, // @[:@149467.4]
  input  [63:0] io_ins_477, // @[:@149467.4]
  input  [63:0] io_ins_478, // @[:@149467.4]
  input  [63:0] io_ins_479, // @[:@149467.4]
  input  [63:0] io_ins_480, // @[:@149467.4]
  input  [63:0] io_ins_481, // @[:@149467.4]
  input  [63:0] io_ins_482, // @[:@149467.4]
  input  [63:0] io_ins_483, // @[:@149467.4]
  input  [63:0] io_ins_484, // @[:@149467.4]
  input  [63:0] io_ins_485, // @[:@149467.4]
  input  [63:0] io_ins_486, // @[:@149467.4]
  input  [63:0] io_ins_487, // @[:@149467.4]
  input  [63:0] io_ins_488, // @[:@149467.4]
  input  [63:0] io_ins_489, // @[:@149467.4]
  input  [63:0] io_ins_490, // @[:@149467.4]
  input  [63:0] io_ins_491, // @[:@149467.4]
  input  [63:0] io_ins_492, // @[:@149467.4]
  input  [63:0] io_ins_493, // @[:@149467.4]
  input  [63:0] io_ins_494, // @[:@149467.4]
  input  [63:0] io_ins_495, // @[:@149467.4]
  input  [63:0] io_ins_496, // @[:@149467.4]
  input  [63:0] io_ins_497, // @[:@149467.4]
  input  [63:0] io_ins_498, // @[:@149467.4]
  input  [63:0] io_ins_499, // @[:@149467.4]
  input  [63:0] io_ins_500, // @[:@149467.4]
  input  [63:0] io_ins_501, // @[:@149467.4]
  input  [63:0] io_ins_502, // @[:@149467.4]
  input  [8:0]  io_sel, // @[:@149467.4]
  output [63:0] io_out // @[:@149467.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@149469.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@149469.4]
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@149469.4]
  assign io_out = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@149469.4]
endmodule
module RegFile( // @[:@149471.2]
  input         clock, // @[:@149472.4]
  input         reset, // @[:@149473.4]
  input  [39:0] io_raddr, // @[:@149474.4]
  input         io_wen, // @[:@149474.4]
  input  [39:0] io_waddr, // @[:@149474.4]
  input  [63:0] io_wdata, // @[:@149474.4]
  output [63:0] io_rdata, // @[:@149474.4]
  input         io_reset, // @[:@149474.4]
  output [63:0] io_argIns_0, // @[:@149474.4]
  output [63:0] io_argIns_1, // @[:@149474.4]
  output [63:0] io_argIns_2, // @[:@149474.4]
  output [63:0] io_argIns_3, // @[:@149474.4]
  input         io_argOuts_0_valid, // @[:@149474.4]
  input  [63:0] io_argOuts_0_bits, // @[:@149474.4]
  input         io_argOuts_1_valid, // @[:@149474.4]
  input  [63:0] io_argOuts_1_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_2_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_3_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_4_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_5_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_6_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_7_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_8_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_9_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_10_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_11_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_12_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_13_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_14_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_15_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_16_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_17_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_18_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_19_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_20_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_21_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_22_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_23_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_24_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_25_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_26_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_27_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_28_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_29_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_30_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_31_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_32_bits, // @[:@149474.4]
  input  [63:0] io_argOuts_43_bits, // @[:@149474.4]
  output [63:0] io_argEchos_1 // @[:@149474.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@151484.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@151484.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@151484.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@151484.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@151484.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@151484.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@151496.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@151496.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@151496.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@151496.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@151496.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@151496.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@151515.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@151515.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@151515.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@151515.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@151515.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@151515.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@151527.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@151527.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@151527.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@151527.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@151527.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@151527.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@151539.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@151539.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@151539.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@151539.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@151539.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@151539.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@151553.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@151553.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@151553.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@151553.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@151553.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@151553.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@151567.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@151567.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@151567.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@151567.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@151567.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@151567.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@151581.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@151581.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@151581.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@151581.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@151581.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@151581.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@151595.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@151595.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@151595.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@151595.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@151595.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@151595.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@151609.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@151609.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@151609.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@151609.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@151609.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@151609.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@151623.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@151623.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@151623.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@151623.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@151623.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@151623.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@151637.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@151637.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@151637.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@151637.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@151637.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@151637.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@151651.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@151651.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@151651.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@151651.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@151651.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@151651.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@151665.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@151665.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@151665.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@151665.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@151665.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@151665.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@151679.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@151679.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@151679.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@151679.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@151679.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@151679.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@151693.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@151693.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@151693.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@151693.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@151693.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@151693.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@151707.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@151707.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@151707.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@151707.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@151707.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@151707.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@151721.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@151721.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@151721.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@151721.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@151721.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@151721.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@151735.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@151735.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@151735.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@151735.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@151735.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@151735.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@151749.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@151749.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@151749.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@151749.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@151749.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@151749.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@151763.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@151763.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@151763.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@151763.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@151763.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@151763.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@151777.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@151777.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@151777.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@151777.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@151777.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@151777.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@151791.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@151791.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@151791.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@151791.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@151791.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@151791.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@151805.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@151805.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@151805.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@151805.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@151805.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@151805.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@151819.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@151819.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@151819.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@151819.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@151819.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@151819.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@151833.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@151833.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@151833.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@151833.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@151833.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@151833.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@151847.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@151847.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@151847.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@151847.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@151847.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@151847.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@151861.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@151861.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@151861.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@151861.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@151861.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@151861.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@151875.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@151875.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@151875.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@151875.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@151875.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@151875.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@151889.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@151889.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@151889.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@151889.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@151889.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@151889.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@151903.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@151903.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@151903.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@151903.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@151903.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@151903.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@151917.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@151917.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@151917.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@151917.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@151917.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@151917.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@151931.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@151931.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@151931.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@151931.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@151931.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@151931.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@151945.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@151945.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@151945.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@151945.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@151945.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@151945.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@151959.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@151959.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@151959.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@151959.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@151959.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@151959.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@151973.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@151973.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@151973.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@151973.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@151973.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@151973.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@151987.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@151987.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@151987.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@151987.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@151987.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@151987.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@152001.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@152001.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@152001.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@152001.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@152001.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@152001.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@152015.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@152015.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@152015.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@152015.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@152015.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@152015.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@152029.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@152029.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@152029.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@152029.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@152029.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@152029.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@152043.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@152043.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@152043.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@152043.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@152043.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@152043.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@152057.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@152057.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@152057.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@152057.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@152057.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@152057.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@152071.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@152071.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@152071.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@152071.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@152071.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@152071.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@152085.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@152085.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@152085.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@152085.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@152085.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@152085.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@152099.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@152099.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@152099.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@152099.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@152099.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@152099.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@152113.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@152113.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@152113.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@152113.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@152113.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@152113.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@152127.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@152127.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@152127.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@152127.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@152127.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@152127.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@152141.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@152141.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@152141.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@152141.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@152141.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@152141.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@152155.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@152155.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@152155.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@152155.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@152155.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@152155.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@152169.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@152169.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@152169.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@152169.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@152169.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@152169.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@152183.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@152183.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@152183.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@152183.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@152183.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@152183.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@152197.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@152197.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@152197.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@152197.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@152197.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@152197.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@152211.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@152211.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@152211.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@152211.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@152211.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@152211.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@152225.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@152225.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@152225.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@152225.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@152225.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@152225.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@152239.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@152239.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@152239.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@152239.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@152239.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@152239.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@152253.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@152253.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@152253.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@152253.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@152253.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@152253.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@152267.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@152267.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@152267.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@152267.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@152267.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@152267.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@152281.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@152281.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@152281.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@152281.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@152281.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@152281.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@152295.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@152295.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@152295.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@152295.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@152295.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@152295.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@152309.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@152309.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@152309.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@152309.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@152309.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@152309.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@152323.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@152323.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@152323.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@152323.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@152323.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@152323.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@152337.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@152337.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@152337.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@152337.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@152337.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@152337.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@152351.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@152351.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@152351.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@152351.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@152351.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@152351.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@152365.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@152365.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@152365.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@152365.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@152365.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@152365.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@152379.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@152379.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@152379.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@152379.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@152379.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@152379.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@152393.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@152393.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@152393.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@152393.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@152393.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@152393.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@152407.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@152407.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@152407.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@152407.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@152407.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@152407.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@152421.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@152421.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@152421.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@152421.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@152421.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@152421.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@152435.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@152435.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@152435.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@152435.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@152435.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@152435.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@152449.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@152449.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@152449.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@152449.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@152449.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@152449.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@152463.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@152463.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@152463.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@152463.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@152463.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@152463.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@152477.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@152477.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@152477.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@152477.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@152477.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@152477.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@152491.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@152491.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@152491.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@152491.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@152491.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@152491.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@152505.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@152505.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@152505.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@152505.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@152505.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@152505.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@152519.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@152519.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@152519.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@152519.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@152519.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@152519.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@152533.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@152533.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@152533.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@152533.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@152533.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@152533.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@152547.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@152547.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@152547.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@152547.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@152547.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@152547.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@152561.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@152561.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@152561.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@152561.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@152561.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@152561.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@152575.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@152575.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@152575.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@152575.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@152575.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@152575.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@152589.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@152589.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@152589.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@152589.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@152589.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@152589.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@152603.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@152603.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@152603.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@152603.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@152603.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@152603.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@152617.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@152617.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@152617.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@152617.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@152617.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@152617.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@152631.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@152631.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@152631.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@152631.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@152631.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@152631.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@152645.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@152645.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@152645.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@152645.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@152645.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@152645.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@152659.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@152659.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@152659.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@152659.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@152659.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@152659.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@152673.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@152673.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@152673.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@152673.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@152673.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@152673.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@152687.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@152687.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@152687.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@152687.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@152687.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@152687.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@152701.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@152701.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@152701.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@152701.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@152701.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@152701.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@152715.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@152715.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@152715.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@152715.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@152715.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@152715.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@152729.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@152729.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@152729.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@152729.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@152729.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@152729.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@152743.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@152743.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@152743.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@152743.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@152743.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@152743.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@152757.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@152757.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@152757.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@152757.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@152757.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@152757.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@152771.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@152771.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@152771.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@152771.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@152771.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@152771.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@152785.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@152785.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@152785.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@152785.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@152785.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@152785.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@152799.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@152799.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@152799.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@152799.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@152799.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@152799.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@152813.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@152813.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@152813.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@152813.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@152813.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@152813.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@152827.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@152827.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@152827.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@152827.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@152827.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@152827.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@152841.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@152841.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@152841.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@152841.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@152841.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@152841.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@152855.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@152855.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@152855.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@152855.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@152855.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@152855.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@152869.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@152869.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@152869.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@152869.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@152869.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@152869.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@152883.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@152883.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@152883.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@152883.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@152883.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@152883.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@152897.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@152897.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@152897.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@152897.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@152897.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@152897.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@152911.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@152911.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@152911.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@152911.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@152911.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@152911.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@152925.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@152925.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@152925.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@152925.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@152925.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@152925.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@152939.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@152939.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@152939.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@152939.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@152939.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@152939.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@152953.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@152953.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@152953.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@152953.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@152953.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@152953.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@152967.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@152967.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@152967.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@152967.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@152967.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@152967.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@152981.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@152981.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@152981.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@152981.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@152981.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@152981.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@152995.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@152995.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@152995.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@152995.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@152995.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@152995.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@153009.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@153009.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@153009.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@153009.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@153009.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@153009.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@153023.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@153023.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@153023.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@153023.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@153023.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@153023.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@153037.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@153037.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@153037.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@153037.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@153037.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@153037.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@153051.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@153051.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@153051.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@153051.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@153051.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@153051.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@153065.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@153065.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@153065.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@153065.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@153065.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@153065.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@153079.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@153079.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@153079.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@153079.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@153079.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@153079.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@153093.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@153093.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@153093.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@153093.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@153093.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@153093.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@153107.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@153107.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@153107.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@153107.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@153107.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@153107.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@153121.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@153121.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@153121.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@153121.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@153121.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@153121.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@153135.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@153135.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@153135.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@153135.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@153135.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@153135.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@153149.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@153149.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@153149.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@153149.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@153149.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@153149.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@153163.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@153163.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@153163.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@153163.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@153163.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@153163.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@153177.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@153177.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@153177.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@153177.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@153177.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@153177.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@153191.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@153191.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@153191.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@153191.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@153191.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@153191.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@153205.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@153205.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@153205.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@153205.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@153205.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@153205.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@153219.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@153219.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@153219.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@153219.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@153219.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@153219.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@153233.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@153233.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@153233.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@153233.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@153233.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@153233.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@153247.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@153247.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@153247.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@153247.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@153247.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@153247.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@153261.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@153261.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@153261.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@153261.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@153261.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@153261.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@153275.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@153275.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@153275.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@153275.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@153275.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@153275.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@153289.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@153289.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@153289.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@153289.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@153289.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@153289.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@153303.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@153303.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@153303.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@153303.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@153303.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@153303.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@153317.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@153317.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@153317.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@153317.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@153317.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@153317.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@153331.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@153331.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@153331.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@153331.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@153331.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@153331.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@153345.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@153345.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@153345.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@153345.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@153345.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@153345.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@153359.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@153359.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@153359.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@153359.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@153359.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@153359.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@153373.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@153373.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@153373.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@153373.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@153373.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@153373.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@153387.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@153387.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@153387.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@153387.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@153387.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@153387.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@153401.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@153401.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@153401.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@153401.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@153401.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@153401.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@153415.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@153415.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@153415.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@153415.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@153415.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@153415.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@153429.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@153429.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@153429.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@153429.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@153429.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@153429.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@153443.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@153443.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@153443.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@153443.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@153443.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@153443.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@153457.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@153457.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@153457.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@153457.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@153457.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@153457.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@153471.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@153471.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@153471.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@153471.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@153471.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@153471.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@153485.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@153485.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@153485.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@153485.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@153485.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@153485.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@153499.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@153499.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@153499.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@153499.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@153499.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@153499.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@153513.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@153513.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@153513.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@153513.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@153513.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@153513.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@153527.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@153527.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@153527.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@153527.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@153527.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@153527.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@153541.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@153541.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@153541.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@153541.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@153541.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@153541.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@153555.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@153555.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@153555.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@153555.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@153555.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@153555.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@153569.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@153569.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@153569.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@153569.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@153569.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@153569.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@153583.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@153583.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@153583.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@153583.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@153583.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@153583.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@153597.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@153597.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@153597.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@153597.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@153597.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@153597.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@153611.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@153611.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@153611.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@153611.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@153611.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@153611.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@153625.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@153625.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@153625.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@153625.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@153625.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@153625.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@153639.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@153639.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@153639.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@153639.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@153639.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@153639.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@153653.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@153653.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@153653.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@153653.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@153653.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@153653.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@153667.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@153667.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@153667.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@153667.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@153667.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@153667.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@153681.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@153681.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@153681.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@153681.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@153681.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@153681.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@153695.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@153695.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@153695.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@153695.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@153695.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@153695.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@153709.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@153709.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@153709.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@153709.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@153709.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@153709.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@153723.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@153723.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@153723.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@153723.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@153723.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@153723.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@153737.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@153737.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@153737.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@153737.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@153737.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@153737.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@153751.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@153751.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@153751.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@153751.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@153751.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@153751.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@153765.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@153765.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@153765.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@153765.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@153765.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@153765.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@153779.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@153779.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@153779.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@153779.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@153779.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@153779.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@153793.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@153793.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@153793.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@153793.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@153793.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@153793.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@153807.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@153807.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@153807.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@153807.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@153807.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@153807.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@153821.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@153821.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@153821.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@153821.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@153821.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@153821.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@153835.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@153835.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@153835.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@153835.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@153835.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@153835.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@153849.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@153849.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@153849.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@153849.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@153849.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@153849.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@153863.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@153863.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@153863.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@153863.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@153863.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@153863.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@153877.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@153877.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@153877.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@153877.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@153877.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@153877.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@153891.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@153891.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@153891.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@153891.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@153891.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@153891.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@153905.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@153905.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@153905.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@153905.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@153905.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@153905.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@153919.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@153919.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@153919.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@153919.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@153919.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@153919.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@153933.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@153933.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@153933.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@153933.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@153933.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@153933.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@153947.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@153947.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@153947.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@153947.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@153947.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@153947.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@153961.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@153961.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@153961.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@153961.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@153961.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@153961.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@153975.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@153975.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@153975.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@153975.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@153975.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@153975.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@153989.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@153989.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@153989.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@153989.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@153989.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@153989.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@154003.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@154003.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@154003.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@154003.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@154003.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@154003.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@154017.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@154017.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@154017.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@154017.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@154017.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@154017.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@154031.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@154031.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@154031.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@154031.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@154031.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@154031.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@154045.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@154045.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@154045.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@154045.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@154045.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@154045.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@154059.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@154059.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@154059.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@154059.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@154059.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@154059.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@154073.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@154073.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@154073.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@154073.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@154073.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@154073.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@154087.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@154087.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@154087.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@154087.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@154087.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@154087.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@154101.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@154101.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@154101.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@154101.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@154101.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@154101.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@154115.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@154115.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@154115.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@154115.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@154115.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@154115.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@154129.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@154129.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@154129.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@154129.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@154129.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@154129.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@154143.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@154143.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@154143.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@154143.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@154143.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@154143.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@154157.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@154157.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@154157.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@154157.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@154157.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@154157.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@154171.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@154171.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@154171.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@154171.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@154171.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@154171.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@154185.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@154185.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@154185.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@154185.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@154185.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@154185.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@154199.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@154199.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@154199.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@154199.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@154199.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@154199.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@154213.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@154213.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@154213.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@154213.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@154213.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@154213.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@154227.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@154227.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@154227.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@154227.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@154227.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@154227.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@154241.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@154241.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@154241.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@154241.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@154241.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@154241.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@154255.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@154255.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@154255.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@154255.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@154255.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@154255.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@154269.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@154269.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@154269.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@154269.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@154269.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@154269.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@154283.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@154283.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@154283.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@154283.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@154283.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@154283.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@154297.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@154297.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@154297.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@154297.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@154297.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@154297.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@154311.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@154311.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@154311.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@154311.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@154311.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@154311.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@154325.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@154325.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@154325.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@154325.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@154325.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@154325.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@154339.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@154339.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@154339.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@154339.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@154339.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@154339.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@154353.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@154353.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@154353.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@154353.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@154353.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@154353.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@154367.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@154367.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@154367.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@154367.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@154367.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@154367.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@154381.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@154381.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@154381.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@154381.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@154381.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@154381.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@154395.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@154395.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@154395.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@154395.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@154395.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@154395.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@154409.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@154409.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@154409.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@154409.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@154409.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@154409.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@154423.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@154423.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@154423.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@154423.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@154423.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@154423.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@154437.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@154437.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@154437.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@154437.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@154437.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@154437.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@154451.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@154451.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@154451.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@154451.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@154451.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@154451.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@154465.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@154465.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@154465.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@154465.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@154465.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@154465.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@154479.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@154479.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@154479.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@154479.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@154479.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@154479.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@154493.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@154493.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@154493.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@154493.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@154493.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@154493.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@154507.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@154507.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@154507.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@154507.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@154507.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@154507.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@154521.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@154521.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@154521.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@154521.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@154521.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@154521.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@154535.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@154535.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@154535.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@154535.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@154535.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@154535.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@154549.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@154549.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@154549.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@154549.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@154549.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@154549.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@154563.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@154563.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@154563.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@154563.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@154563.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@154563.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@154577.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@154577.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@154577.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@154577.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@154577.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@154577.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@154591.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@154591.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@154591.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@154591.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@154591.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@154591.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@154605.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@154605.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@154605.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@154605.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@154605.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@154605.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@154619.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@154619.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@154619.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@154619.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@154619.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@154619.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@154633.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@154633.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@154633.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@154633.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@154633.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@154633.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@154647.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@154647.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@154647.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@154647.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@154647.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@154647.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@154661.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@154661.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@154661.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@154661.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@154661.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@154661.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@154675.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@154675.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@154675.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@154675.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@154675.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@154675.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@154689.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@154689.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@154689.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@154689.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@154689.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@154689.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@154703.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@154703.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@154703.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@154703.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@154703.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@154703.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@154717.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@154717.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@154717.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@154717.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@154717.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@154717.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@154731.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@154731.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@154731.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@154731.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@154731.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@154731.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@154745.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@154745.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@154745.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@154745.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@154745.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@154745.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@154759.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@154759.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@154759.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@154759.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@154759.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@154759.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@154773.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@154773.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@154773.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@154773.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@154773.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@154773.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@154787.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@154787.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@154787.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@154787.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@154787.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@154787.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@154801.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@154801.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@154801.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@154801.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@154801.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@154801.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@154815.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@154815.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@154815.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@154815.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@154815.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@154815.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@154829.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@154829.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@154829.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@154829.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@154829.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@154829.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@154843.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@154843.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@154843.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@154843.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@154843.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@154843.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@154857.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@154857.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@154857.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@154857.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@154857.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@154857.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@154871.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@154871.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@154871.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@154871.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@154871.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@154871.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@154885.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@154885.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@154885.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@154885.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@154885.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@154885.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@154899.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@154899.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@154899.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@154899.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@154899.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@154899.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@154913.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@154913.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@154913.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@154913.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@154913.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@154913.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@154927.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@154927.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@154927.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@154927.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@154927.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@154927.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@154941.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@154941.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@154941.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@154941.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@154941.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@154941.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@154955.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@154955.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@154955.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@154955.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@154955.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@154955.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@154969.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@154969.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@154969.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@154969.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@154969.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@154969.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@154983.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@154983.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@154983.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@154983.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@154983.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@154983.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@154997.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@154997.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@154997.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@154997.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@154997.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@154997.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@155011.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@155011.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@155011.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@155011.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@155011.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@155011.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@155025.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@155025.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@155025.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@155025.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@155025.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@155025.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@155039.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@155039.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@155039.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@155039.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@155039.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@155039.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@155053.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@155053.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@155053.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@155053.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@155053.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@155053.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@155067.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@155067.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@155067.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@155067.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@155067.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@155067.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@155081.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@155081.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@155081.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@155081.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@155081.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@155081.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@155095.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@155095.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@155095.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@155095.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@155095.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@155095.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@155109.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@155109.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@155109.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@155109.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@155109.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@155109.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@155123.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@155123.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@155123.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@155123.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@155123.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@155123.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@155137.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@155137.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@155137.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@155137.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@155137.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@155137.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@155151.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@155151.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@155151.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@155151.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@155151.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@155151.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@155165.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@155165.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@155165.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@155165.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@155165.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@155165.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@155179.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@155179.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@155179.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@155179.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@155179.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@155179.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@155193.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@155193.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@155193.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@155193.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@155193.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@155193.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@155207.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@155207.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@155207.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@155207.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@155207.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@155207.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@155221.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@155221.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@155221.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@155221.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@155221.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@155221.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@155235.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@155235.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@155235.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@155235.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@155235.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@155235.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@155249.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@155249.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@155249.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@155249.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@155249.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@155249.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@155263.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@155263.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@155263.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@155263.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@155263.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@155263.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@155277.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@155277.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@155277.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@155277.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@155277.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@155277.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@155291.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@155291.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@155291.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@155291.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@155291.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@155291.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@155305.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@155305.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@155305.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@155305.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@155305.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@155305.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@155319.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@155319.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@155319.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@155319.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@155319.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@155319.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@155333.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@155333.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@155333.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@155333.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@155333.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@155333.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@155347.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@155347.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@155347.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@155347.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@155347.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@155347.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@155361.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@155361.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@155361.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@155361.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@155361.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@155361.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@155375.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@155375.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@155375.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@155375.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@155375.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@155375.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@155389.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@155389.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@155389.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@155389.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@155389.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@155389.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@155403.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@155403.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@155403.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@155403.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@155403.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@155403.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@155417.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@155417.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@155417.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@155417.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@155417.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@155417.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@155431.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@155431.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@155431.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@155431.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@155431.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@155431.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@155445.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@155445.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@155445.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@155445.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@155445.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@155445.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@155459.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@155459.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@155459.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@155459.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@155459.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@155459.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@155473.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@155473.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@155473.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@155473.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@155473.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@155473.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@155487.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@155487.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@155487.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@155487.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@155487.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@155487.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@155501.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@155501.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@155501.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@155501.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@155501.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@155501.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@155515.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@155515.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@155515.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@155515.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@155515.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@155515.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@155529.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@155529.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@155529.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@155529.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@155529.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@155529.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@155543.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@155543.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@155543.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@155543.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@155543.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@155543.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@155557.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@155557.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@155557.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@155557.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@155557.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@155557.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@155571.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@155571.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@155571.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@155571.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@155571.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@155571.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@155585.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@155585.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@155585.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@155585.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@155585.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@155585.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@155599.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@155599.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@155599.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@155599.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@155599.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@155599.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@155613.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@155613.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@155613.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@155613.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@155613.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@155613.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@155627.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@155627.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@155627.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@155627.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@155627.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@155627.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@155641.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@155641.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@155641.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@155641.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@155641.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@155641.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@155655.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@155655.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@155655.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@155655.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@155655.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@155655.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@155669.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@155669.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@155669.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@155669.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@155669.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@155669.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@155683.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@155683.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@155683.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@155683.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@155683.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@155683.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@155697.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@155697.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@155697.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@155697.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@155697.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@155697.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@155711.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@155711.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@155711.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@155711.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@155711.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@155711.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@155725.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@155725.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@155725.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@155725.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@155725.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@155725.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@155739.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@155739.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@155739.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@155739.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@155739.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@155739.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@155753.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@155753.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@155753.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@155753.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@155753.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@155753.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@155767.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@155767.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@155767.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@155767.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@155767.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@155767.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@155781.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@155781.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@155781.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@155781.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@155781.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@155781.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@155795.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@155795.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@155795.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@155795.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@155795.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@155795.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@155809.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@155809.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@155809.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@155809.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@155809.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@155809.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@155823.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@155823.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@155823.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@155823.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@155823.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@155823.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@155837.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@155837.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@155837.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@155837.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@155837.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@155837.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@155851.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@155851.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@155851.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@155851.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@155851.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@155851.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@155865.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@155865.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@155865.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@155865.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@155865.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@155865.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@155879.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@155879.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@155879.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@155879.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@155879.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@155879.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@155893.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@155893.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@155893.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@155893.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@155893.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@155893.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@155907.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@155907.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@155907.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@155907.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@155907.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@155907.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@155921.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@155921.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@155921.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@155921.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@155921.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@155921.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@155935.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@155935.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@155935.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@155935.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@155935.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@155935.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@155949.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@155949.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@155949.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@155949.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@155949.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@155949.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@155963.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@155963.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@155963.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@155963.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@155963.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@155963.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@155977.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@155977.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@155977.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@155977.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@155977.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@155977.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@155991.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@155991.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@155991.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@155991.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@155991.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@155991.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@156005.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@156005.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@156005.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@156005.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@156005.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@156005.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@156019.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@156019.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@156019.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@156019.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@156019.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@156019.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@156033.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@156033.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@156033.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@156033.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@156033.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@156033.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@156047.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@156047.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@156047.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@156047.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@156047.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@156047.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@156061.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@156061.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@156061.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@156061.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@156061.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@156061.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@156075.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@156075.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@156075.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@156075.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@156075.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@156075.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@156089.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@156089.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@156089.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@156089.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@156089.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@156089.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@156103.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@156103.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@156103.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@156103.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@156103.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@156103.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@156117.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@156117.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@156117.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@156117.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@156117.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@156117.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@156131.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@156131.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@156131.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@156131.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@156131.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@156131.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@156145.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@156145.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@156145.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@156145.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@156145.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@156145.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@156159.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@156159.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@156159.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@156159.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@156159.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@156159.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@156173.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@156173.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@156173.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@156173.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@156173.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@156173.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@156187.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@156187.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@156187.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@156187.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@156187.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@156187.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@156201.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@156201.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@156201.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@156201.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@156201.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@156201.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@156215.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@156215.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@156215.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@156215.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@156215.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@156215.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@156229.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@156229.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@156229.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@156229.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@156229.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@156229.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@156243.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@156243.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@156243.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@156243.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@156243.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@156243.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@156257.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@156257.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@156257.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@156257.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@156257.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@156257.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@156271.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@156271.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@156271.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@156271.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@156271.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@156271.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@156285.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@156285.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@156285.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@156285.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@156285.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@156285.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@156299.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@156299.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@156299.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@156299.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@156299.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@156299.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@156313.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@156313.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@156313.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@156313.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@156313.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@156313.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@156327.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@156327.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@156327.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@156327.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@156327.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@156327.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@156341.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@156341.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@156341.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@156341.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@156341.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@156341.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@156355.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@156355.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@156355.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@156355.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@156355.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@156355.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@156369.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@156369.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@156369.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@156369.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@156369.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@156369.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@156383.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@156383.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@156383.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@156383.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@156383.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@156383.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@156397.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@156397.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@156397.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@156397.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@156397.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@156397.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@156411.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@156411.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@156411.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@156411.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@156411.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@156411.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@156425.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@156425.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@156425.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@156425.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@156425.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@156425.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@156439.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@156439.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@156439.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@156439.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@156439.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@156439.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@156453.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@156453.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@156453.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@156453.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@156453.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@156453.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@156467.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@156467.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@156467.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@156467.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@156467.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@156467.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@156481.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@156481.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@156481.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@156481.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@156481.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@156481.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@156495.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@156495.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@156495.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@156495.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@156495.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@156495.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@156509.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@156509.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@156509.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@156509.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@156509.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@156509.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@156523.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@156523.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@156523.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@156523.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@156523.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@156523.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@156537.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@156537.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@156537.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@156537.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@156537.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@156537.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@156551.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@156551.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@156551.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@156551.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@156551.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@156551.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@156565.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@156565.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@156565.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@156565.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@156565.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@156565.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@156579.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@156579.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@156579.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@156579.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@156579.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@156579.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@156593.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@156593.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@156593.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@156593.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@156593.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@156593.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@156607.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@156607.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@156607.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@156607.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@156607.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@156607.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@156621.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@156621.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@156621.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@156621.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@156621.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@156621.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@156635.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@156635.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@156635.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@156635.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@156635.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@156635.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@156649.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@156649.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@156649.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@156649.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@156649.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@156649.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@156663.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@156663.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@156663.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@156663.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@156663.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@156663.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@156677.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@156677.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@156677.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@156677.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@156677.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@156677.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@156691.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@156691.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@156691.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@156691.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@156691.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@156691.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@156705.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@156705.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@156705.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@156705.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@156705.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@156705.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@156719.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@156719.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@156719.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@156719.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@156719.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@156719.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@156733.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@156733.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@156733.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@156733.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@156733.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@156733.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@156747.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@156747.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@156747.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@156747.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@156747.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@156747.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@156761.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@156761.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@156761.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@156761.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@156761.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@156761.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@156775.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@156775.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@156775.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@156775.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@156775.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@156775.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@156789.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@156789.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@156789.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@156789.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@156789.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@156789.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@156803.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@156803.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@156803.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@156803.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@156803.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@156803.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@156817.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@156817.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@156817.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@156817.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@156817.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@156817.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@156831.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@156831.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@156831.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@156831.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@156831.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@156831.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@156845.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@156845.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@156845.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@156845.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@156845.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@156845.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@156859.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@156859.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@156859.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@156859.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@156859.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@156859.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@156873.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@156873.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@156873.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@156873.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@156873.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@156873.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@156887.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@156887.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@156887.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@156887.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@156887.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@156887.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@156901.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@156901.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@156901.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@156901.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@156901.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@156901.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@156915.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@156915.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@156915.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@156915.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@156915.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@156915.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@156929.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@156929.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@156929.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@156929.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@156929.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@156929.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@156943.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@156943.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@156943.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@156943.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@156943.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@156943.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@156957.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@156957.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@156957.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@156957.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@156957.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@156957.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@156971.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@156971.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@156971.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@156971.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@156971.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@156971.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@156985.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@156985.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@156985.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@156985.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@156985.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@156985.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@156999.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@156999.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@156999.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@156999.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@156999.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@156999.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@157013.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@157013.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@157013.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@157013.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@157013.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@157013.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@157027.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@157027.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@157027.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@157027.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@157027.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@157027.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@157041.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@157041.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@157041.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@157041.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@157041.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@157041.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@157055.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@157055.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@157055.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@157055.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@157055.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@157055.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@157069.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@157069.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@157069.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@157069.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@157069.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@157069.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@157083.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@157083.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@157083.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@157083.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@157083.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@157083.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@157097.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@157097.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@157097.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@157097.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@157097.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@157097.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@157111.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@157111.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@157111.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@157111.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@157111.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@157111.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@157125.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@157125.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@157125.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@157125.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@157125.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@157125.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@157139.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@157139.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@157139.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@157139.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@157139.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@157139.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@157153.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@157153.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@157153.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@157153.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@157153.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@157153.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@157167.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@157167.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@157167.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@157167.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@157167.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@157167.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@157181.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@157181.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@157181.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@157181.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@157181.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@157181.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@157195.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@157195.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@157195.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@157195.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@157195.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@157195.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@157209.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@157209.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@157209.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@157209.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@157209.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@157209.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@157223.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@157223.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@157223.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@157223.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@157223.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@157223.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@157237.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@157237.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@157237.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@157237.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@157237.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@157237.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@157251.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@157251.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@157251.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@157251.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@157251.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@157251.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@157265.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@157265.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@157265.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@157265.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@157265.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@157265.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@157279.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@157279.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@157279.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@157279.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@157279.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@157279.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@157293.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@157293.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@157293.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@157293.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@157293.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@157293.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@157307.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@157307.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@157307.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@157307.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@157307.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@157307.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@157321.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@157321.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@157321.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@157321.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@157321.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@157321.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@157335.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@157335.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@157335.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@157335.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@157335.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@157335.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@157349.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@157349.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@157349.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@157349.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@157349.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@157349.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@157363.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@157363.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@157363.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@157363.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@157363.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@157363.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@157377.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@157377.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@157377.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@157377.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@157377.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@157377.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@157391.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@157391.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@157391.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@157391.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@157391.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@157391.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@157405.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@157405.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@157405.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@157405.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@157405.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@157405.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@157419.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@157419.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@157419.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@157419.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@157419.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@157419.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@157433.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@157433.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@157433.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@157433.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@157433.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@157433.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@157447.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@157447.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@157447.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@157447.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@157447.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@157447.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@157461.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@157461.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@157461.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@157461.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@157461.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@157461.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@157475.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@157475.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@157475.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@157475.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@157475.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@157475.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@157489.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@157489.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@157489.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@157489.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@157489.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@157489.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@157503.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@157503.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@157503.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@157503.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@157503.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@157503.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@157517.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@157517.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@157517.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@157517.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@157517.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@157517.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@157531.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@157531.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@157531.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@157531.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@157531.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@157531.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@157545.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@157545.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@157545.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@157545.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@157545.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@157545.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@157559.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@157559.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@157559.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@157559.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@157559.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@157559.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@157573.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@157573.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@157573.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@157573.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@157573.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@157573.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@157587.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@157587.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@157587.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@157587.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@157587.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@157587.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@157601.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@157601.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@157601.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@157601.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@157601.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@157601.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@157615.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@157615.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@157615.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@157615.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@157615.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@157615.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@157629.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@157629.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@157629.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@157629.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@157629.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@157629.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@157643.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@157643.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@157643.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@157643.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@157643.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@157643.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@157657.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@157657.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@157657.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@157657.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@157657.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@157657.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@157671.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@157671.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@157671.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@157671.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@157671.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@157671.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@157685.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@157685.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@157685.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@157685.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@157685.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@157685.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@157699.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@157699.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@157699.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@157699.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@157699.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@157699.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@157713.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@157713.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@157713.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@157713.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@157713.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@157713.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@157727.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@157727.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@157727.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@157727.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@157727.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@157727.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@157741.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@157741.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@157741.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@157741.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@157741.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@157741.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@157755.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@157755.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@157755.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@157755.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@157755.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@157755.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@157769.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@157769.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@157769.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@157769.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@157769.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@157769.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@157783.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@157783.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@157783.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@157783.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@157783.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@157783.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@157797.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@157797.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@157797.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@157797.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@157797.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@157797.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@157811.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@157811.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@157811.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@157811.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@157811.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@157811.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@157825.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@157825.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@157825.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@157825.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@157825.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@157825.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@157839.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@157839.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@157839.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@157839.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@157839.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@157839.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@157853.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@157853.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@157853.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@157853.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@157853.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@157853.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@157867.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@157867.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@157867.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@157867.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@157867.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@157867.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@157881.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@157881.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@157881.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@157881.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@157881.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@157881.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@157895.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@157895.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@157895.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@157895.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@157895.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@157895.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@157909.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@157909.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@157909.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@157909.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@157909.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@157909.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@157923.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@157923.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@157923.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@157923.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@157923.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@157923.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@157937.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@157937.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@157937.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@157937.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@157937.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@157937.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@157951.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@157951.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@157951.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@157951.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@157951.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@157951.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@157965.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@157965.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@157965.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@157965.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@157965.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@157965.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@157979.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@157979.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@157979.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@157979.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@157979.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@157979.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@157993.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@157993.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@157993.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@157993.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@157993.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@157993.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@158007.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@158007.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@158007.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@158007.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@158007.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@158007.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@158021.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@158021.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@158021.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@158021.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@158021.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@158021.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@158035.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@158035.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@158035.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@158035.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@158035.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@158035.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@158049.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@158049.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@158049.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@158049.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@158049.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@158049.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@158063.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@158063.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@158063.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@158063.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@158063.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@158063.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@158077.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@158077.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@158077.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@158077.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@158077.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@158077.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@158091.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@158091.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@158091.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@158091.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@158091.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@158091.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@158105.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@158105.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@158105.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@158105.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@158105.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@158105.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@158119.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@158119.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@158119.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@158119.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@158119.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@158119.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@158133.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@158133.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@158133.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@158133.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@158133.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@158133.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@158147.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@158147.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@158147.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@158147.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@158147.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@158147.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@158161.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@158161.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@158161.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@158161.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@158161.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@158161.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@158175.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@158175.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@158175.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@158175.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@158175.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@158175.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@158189.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@158189.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@158189.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@158189.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@158189.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@158189.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@158203.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@158203.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@158203.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@158203.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@158203.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@158203.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@158217.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@158217.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@158217.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@158217.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@158217.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@158217.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@158231.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@158231.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@158231.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@158231.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@158231.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@158231.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@158245.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@158245.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@158245.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@158245.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@158245.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@158245.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@158259.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@158259.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@158259.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@158259.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@158259.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@158259.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@158273.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@158273.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@158273.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@158273.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@158273.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@158273.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@158287.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@158287.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@158287.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@158287.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@158287.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@158287.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@158301.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@158301.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@158301.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@158301.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@158301.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@158301.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@158315.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@158315.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@158315.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@158315.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@158315.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@158315.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@158329.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@158329.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@158329.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@158329.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@158329.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@158329.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@158343.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@158343.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@158343.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@158343.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@158343.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@158343.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@158357.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@158357.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@158357.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@158357.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@158357.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@158357.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@158371.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@158371.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@158371.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@158371.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@158371.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@158371.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@158385.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@158385.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@158385.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@158385.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@158385.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@158385.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@158399.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@158399.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@158399.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@158399.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@158399.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@158399.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@158413.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@158413.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@158413.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@158413.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@158413.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@158413.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@158427.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@158427.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@158427.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@158427.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@158427.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@158427.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@158441.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@158441.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@158441.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@158441.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@158441.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@158441.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@158455.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@158455.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@158455.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@158455.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@158455.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@158455.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@158469.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@158469.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@158469.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@158469.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@158469.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@158469.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@158483.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@158483.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@158483.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@158483.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@158483.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@158483.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@158497.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@158497.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@158497.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@158497.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@158497.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@158497.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@158511.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@158511.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@158511.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@158511.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@158511.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@158511.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@158525.4]
  wire [8:0] rport_io_sel; // @[RegFile.scala 95:21:@158525.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@158525.4]
  wire  _T_3078; // @[RegFile.scala 80:42:@151487.4]
  wire  _T_3084; // @[RegFile.scala 68:46:@151499.4]
  wire  _T_3085; // @[RegFile.scala 68:34:@151500.4]
  wire  _T_3098; // @[RegFile.scala 80:42:@151518.4]
  wire  _T_3104; // @[RegFile.scala 80:42:@151530.4]
  wire  _T_3110; // @[RegFile.scala 74:80:@151542.4]
  wire  _T_3111; // @[RegFile.scala 74:68:@151543.4]
  wire [39:0] _T_7111; // @[RegFile.scala 99:30:@159535.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@151484.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@151496.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@151515.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@151527.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@151539.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@151553.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@151567.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@151581.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@151595.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@151609.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@151623.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@151637.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@151651.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@151665.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@151679.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@151693.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@151707.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@151721.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@151735.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@151749.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@151763.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@151777.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@151791.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@151805.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@151819.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@151833.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@151847.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@151861.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@151875.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@151889.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@151903.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@151917.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@151931.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@151945.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@151959.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@151973.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@151987.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@152001.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@152015.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@152029.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@152043.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@152057.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@152071.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@152085.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@152099.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@152113.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@152127.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@152141.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@152155.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@152169.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@152183.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@152197.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@152211.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@152225.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@152239.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@152253.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@152267.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@152281.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@152295.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@152309.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@152323.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@152337.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@152351.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@152365.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@152379.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@152393.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@152407.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@152421.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@152435.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@152449.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@152463.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@152477.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@152491.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@152505.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@152519.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@152533.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@152547.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@152561.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@152575.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@152589.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@152603.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@152617.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@152631.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@152645.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@152659.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@152673.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@152687.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@152701.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@152715.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@152729.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@152743.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@152757.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@152771.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@152785.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@152799.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@152813.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@152827.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@152841.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@152855.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@152869.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@152883.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@152897.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@152911.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@152925.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@152939.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@152953.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@152967.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@152981.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@152995.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@153009.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@153023.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@153037.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@153051.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@153065.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@153079.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@153093.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@153107.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@153121.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@153135.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@153149.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@153163.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@153177.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@153191.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@153205.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@153219.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@153233.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@153247.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@153261.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@153275.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@153289.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@153303.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@153317.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@153331.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@153345.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@153359.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@153373.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@153387.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@153401.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@153415.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@153429.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@153443.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@153457.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@153471.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@153485.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@153499.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@153513.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@153527.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@153541.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@153555.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@153569.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@153583.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@153597.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@153611.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@153625.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@153639.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@153653.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@153667.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@153681.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@153695.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@153709.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@153723.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@153737.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@153751.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@153765.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@153779.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@153793.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@153807.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@153821.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@153835.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@153849.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@153863.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@153877.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@153891.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@153905.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@153919.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@153933.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@153947.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@153961.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@153975.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@153989.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@154003.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@154017.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@154031.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@154045.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@154059.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@154073.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@154087.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@154101.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@154115.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@154129.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@154143.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@154157.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@154171.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@154185.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@154199.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@154213.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@154227.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@154241.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@154255.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@154269.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@154283.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@154297.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@154311.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@154325.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@154339.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@154353.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@154367.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@154381.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@154395.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@154409.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@154423.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@154437.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@154451.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@154465.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@154479.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@154493.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@154507.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@154521.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@154535.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@154549.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@154563.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@154577.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@154591.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@154605.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@154619.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@154633.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@154647.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@154661.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@154675.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@154689.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@154703.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@154717.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@154731.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@154745.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@154759.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@154773.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@154787.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@154801.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@154815.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@154829.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@154843.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@154857.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@154871.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@154885.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@154899.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@154913.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@154927.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@154941.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@154955.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@154969.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@154983.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@154997.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@155011.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@155025.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@155039.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@155053.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@155067.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@155081.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@155095.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@155109.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@155123.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@155137.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@155151.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@155165.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@155179.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@155193.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@155207.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@155221.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@155235.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@155249.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@155263.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@155277.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@155291.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@155305.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@155319.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@155333.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@155347.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@155361.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@155375.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@155389.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@155403.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@155417.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@155431.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@155445.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@155459.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@155473.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@155487.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@155501.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@155515.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@155529.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@155543.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@155557.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@155571.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@155585.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@155599.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@155613.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@155627.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@155641.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@155655.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@155669.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@155683.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@155697.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@155711.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@155725.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@155739.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@155753.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@155767.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@155781.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@155795.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@155809.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@155823.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@155837.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@155851.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@155865.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@155879.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@155893.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@155907.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@155921.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@155935.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@155949.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@155963.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@155977.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@155991.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@156005.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@156019.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@156033.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@156047.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@156061.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@156075.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@156089.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@156103.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@156117.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@156131.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@156145.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@156159.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@156173.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@156187.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@156201.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@156215.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@156229.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@156243.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@156257.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@156271.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@156285.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@156299.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@156313.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@156327.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@156341.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@156355.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@156369.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@156383.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@156397.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@156411.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@156425.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@156439.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@156453.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@156467.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@156481.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@156495.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@156509.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@156523.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@156537.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@156551.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@156565.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@156579.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@156593.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@156607.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@156621.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@156635.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@156649.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@156663.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@156677.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@156691.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@156705.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@156719.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@156733.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@156747.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@156761.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@156775.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@156789.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@156803.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@156817.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@156831.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@156845.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@156859.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@156873.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@156887.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@156901.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@156915.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@156929.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@156943.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@156957.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@156971.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@156985.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@156999.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@157013.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@157027.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@157041.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@157055.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@157069.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@157083.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@157097.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@157111.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@157125.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@157139.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@157153.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@157167.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@157181.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@157195.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@157209.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@157223.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@157237.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@157251.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@157265.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@157279.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@157293.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@157307.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@157321.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@157335.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@157349.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@157363.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@157377.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@157391.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@157405.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@157419.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@157433.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@157447.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@157461.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@157475.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@157489.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@157503.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@157517.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@157531.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@157545.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@157559.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@157573.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@157587.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@157601.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@157615.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@157629.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@157643.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@157657.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@157671.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@157685.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@157699.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@157713.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@157727.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@157741.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@157755.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@157769.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@157783.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@157797.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@157811.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@157825.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@157839.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@157853.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@157867.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@157881.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@157895.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@157909.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@157923.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@157937.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@157951.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@157965.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@157979.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@157993.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@158007.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@158021.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@158035.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@158049.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@158063.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@158077.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@158091.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@158105.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@158119.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@158133.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@158147.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@158161.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@158175.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@158189.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@158203.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@158217.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@158231.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@158245.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@158259.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@158273.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@158287.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@158301.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@158315.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@158329.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@158343.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@158357.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@158371.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@158385.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@158399.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@158413.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@158427.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@158441.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@158455.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@158469.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@158483.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@158497.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@158511.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  MuxN_4 rport ( // @[RegFile.scala 95:21:@158525.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3078 = io_waddr == 40'h0; // @[RegFile.scala 80:42:@151487.4]
  assign _T_3084 = io_waddr == 40'h2; // @[RegFile.scala 68:46:@151499.4]
  assign _T_3085 = io_wen & _T_3084; // @[RegFile.scala 68:34:@151500.4]
  assign _T_3098 = io_waddr == 40'h4; // @[RegFile.scala 80:42:@151518.4]
  assign _T_3104 = io_waddr == 40'h6; // @[RegFile.scala 80:42:@151530.4]
  assign _T_3110 = io_waddr == 40'h8; // @[RegFile.scala 74:80:@151542.4]
  assign _T_3111 = io_wen & _T_3110; // @[RegFile.scala 74:68:@151543.4]
  assign _T_7111 = io_raddr / 40'h2; // @[RegFile.scala 99:30:@159535.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 100:14:@159537.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@159543.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@159544.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@159545.4]
  assign io_argIns_3 = regs_3_io_out; // @[RegFile.scala 111:13:@159546.4]
  assign io_argEchos_1 = regs_4_io_out; // @[RegFile.scala 77:37:@151549.4]
  assign regs_0_clock = clock; // @[:@151485.4]
  assign regs_0_reset = reset; // @[:@151486.4 RegFile.scala 82:16:@151492.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@151490.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@151494.4]
  assign regs_0_io_enable = io_wen & _T_3078; // @[RegFile.scala 80:20:@151489.4]
  assign regs_1_clock = clock; // @[:@151497.4]
  assign regs_1_reset = reset; // @[:@151498.4 RegFile.scala 70:16:@151510.4]
  assign regs_1_io_in = _T_3085 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@151508.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@151513.4]
  assign regs_1_io_enable = _T_3085 ? _T_3085 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@151504.4]
  assign regs_2_clock = clock; // @[:@151516.4]
  assign regs_2_reset = reset; // @[:@151517.4 RegFile.scala 82:16:@151523.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@151521.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@151525.4]
  assign regs_2_io_enable = io_wen & _T_3098; // @[RegFile.scala 80:20:@151520.4]
  assign regs_3_clock = clock; // @[:@151528.4]
  assign regs_3_reset = reset; // @[:@151529.4 RegFile.scala 82:16:@151535.4]
  assign regs_3_io_in = io_wdata; // @[RegFile.scala 81:16:@151533.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 83:19:@151537.4]
  assign regs_3_io_enable = io_wen & _T_3104; // @[RegFile.scala 80:20:@151532.4]
  assign regs_4_clock = clock; // @[:@151540.4]
  assign regs_4_reset = io_reset; // @[:@151541.4 RegFile.scala 76:16:@151548.4]
  assign regs_4_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@151547.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@151551.4]
  assign regs_4_io_enable = io_argOuts_1_valid | _T_3111; // @[RegFile.scala 74:20:@151545.4]
  assign regs_5_clock = clock; // @[:@151554.4]
  assign regs_5_reset = io_reset; // @[:@151555.4 RegFile.scala 76:16:@151562.4]
  assign regs_5_io_in = io_argOuts_2_bits; // @[RegFile.scala 75:16:@151561.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@151565.4]
  assign regs_5_io_enable = 1'h1; // @[RegFile.scala 74:20:@151559.4]
  assign regs_6_clock = clock; // @[:@151568.4]
  assign regs_6_reset = io_reset; // @[:@151569.4 RegFile.scala 76:16:@151576.4]
  assign regs_6_io_in = io_argOuts_3_bits; // @[RegFile.scala 75:16:@151575.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@151579.4]
  assign regs_6_io_enable = 1'h1; // @[RegFile.scala 74:20:@151573.4]
  assign regs_7_clock = clock; // @[:@151582.4]
  assign regs_7_reset = io_reset; // @[:@151583.4 RegFile.scala 76:16:@151590.4]
  assign regs_7_io_in = io_argOuts_4_bits; // @[RegFile.scala 75:16:@151589.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@151593.4]
  assign regs_7_io_enable = 1'h1; // @[RegFile.scala 74:20:@151587.4]
  assign regs_8_clock = clock; // @[:@151596.4]
  assign regs_8_reset = io_reset; // @[:@151597.4 RegFile.scala 76:16:@151604.4]
  assign regs_8_io_in = io_argOuts_5_bits; // @[RegFile.scala 75:16:@151603.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@151607.4]
  assign regs_8_io_enable = 1'h1; // @[RegFile.scala 74:20:@151601.4]
  assign regs_9_clock = clock; // @[:@151610.4]
  assign regs_9_reset = io_reset; // @[:@151611.4 RegFile.scala 76:16:@151618.4]
  assign regs_9_io_in = io_argOuts_6_bits; // @[RegFile.scala 75:16:@151617.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@151621.4]
  assign regs_9_io_enable = 1'h1; // @[RegFile.scala 74:20:@151615.4]
  assign regs_10_clock = clock; // @[:@151624.4]
  assign regs_10_reset = io_reset; // @[:@151625.4 RegFile.scala 76:16:@151632.4]
  assign regs_10_io_in = io_argOuts_7_bits; // @[RegFile.scala 75:16:@151631.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@151635.4]
  assign regs_10_io_enable = 1'h1; // @[RegFile.scala 74:20:@151629.4]
  assign regs_11_clock = clock; // @[:@151638.4]
  assign regs_11_reset = io_reset; // @[:@151639.4 RegFile.scala 76:16:@151646.4]
  assign regs_11_io_in = io_argOuts_8_bits; // @[RegFile.scala 75:16:@151645.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@151649.4]
  assign regs_11_io_enable = 1'h1; // @[RegFile.scala 74:20:@151643.4]
  assign regs_12_clock = clock; // @[:@151652.4]
  assign regs_12_reset = io_reset; // @[:@151653.4 RegFile.scala 76:16:@151660.4]
  assign regs_12_io_in = io_argOuts_9_bits; // @[RegFile.scala 75:16:@151659.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@151663.4]
  assign regs_12_io_enable = 1'h1; // @[RegFile.scala 74:20:@151657.4]
  assign regs_13_clock = clock; // @[:@151666.4]
  assign regs_13_reset = io_reset; // @[:@151667.4 RegFile.scala 76:16:@151674.4]
  assign regs_13_io_in = io_argOuts_10_bits; // @[RegFile.scala 75:16:@151673.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@151677.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 74:20:@151671.4]
  assign regs_14_clock = clock; // @[:@151680.4]
  assign regs_14_reset = io_reset; // @[:@151681.4 RegFile.scala 76:16:@151688.4]
  assign regs_14_io_in = io_argOuts_11_bits; // @[RegFile.scala 75:16:@151687.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@151691.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 74:20:@151685.4]
  assign regs_15_clock = clock; // @[:@151694.4]
  assign regs_15_reset = io_reset; // @[:@151695.4 RegFile.scala 76:16:@151702.4]
  assign regs_15_io_in = io_argOuts_12_bits; // @[RegFile.scala 75:16:@151701.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@151705.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 74:20:@151699.4]
  assign regs_16_clock = clock; // @[:@151708.4]
  assign regs_16_reset = io_reset; // @[:@151709.4 RegFile.scala 76:16:@151716.4]
  assign regs_16_io_in = io_argOuts_13_bits; // @[RegFile.scala 75:16:@151715.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@151719.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 74:20:@151713.4]
  assign regs_17_clock = clock; // @[:@151722.4]
  assign regs_17_reset = io_reset; // @[:@151723.4 RegFile.scala 76:16:@151730.4]
  assign regs_17_io_in = io_argOuts_14_bits; // @[RegFile.scala 75:16:@151729.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@151733.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 74:20:@151727.4]
  assign regs_18_clock = clock; // @[:@151736.4]
  assign regs_18_reset = io_reset; // @[:@151737.4 RegFile.scala 76:16:@151744.4]
  assign regs_18_io_in = io_argOuts_15_bits; // @[RegFile.scala 75:16:@151743.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@151747.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 74:20:@151741.4]
  assign regs_19_clock = clock; // @[:@151750.4]
  assign regs_19_reset = io_reset; // @[:@151751.4 RegFile.scala 76:16:@151758.4]
  assign regs_19_io_in = io_argOuts_16_bits; // @[RegFile.scala 75:16:@151757.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@151761.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@151755.4]
  assign regs_20_clock = clock; // @[:@151764.4]
  assign regs_20_reset = io_reset; // @[:@151765.4 RegFile.scala 76:16:@151772.4]
  assign regs_20_io_in = io_argOuts_17_bits; // @[RegFile.scala 75:16:@151771.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@151775.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@151769.4]
  assign regs_21_clock = clock; // @[:@151778.4]
  assign regs_21_reset = io_reset; // @[:@151779.4 RegFile.scala 76:16:@151786.4]
  assign regs_21_io_in = io_argOuts_18_bits; // @[RegFile.scala 75:16:@151785.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@151789.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@151783.4]
  assign regs_22_clock = clock; // @[:@151792.4]
  assign regs_22_reset = io_reset; // @[:@151793.4 RegFile.scala 76:16:@151800.4]
  assign regs_22_io_in = io_argOuts_19_bits; // @[RegFile.scala 75:16:@151799.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@151803.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@151797.4]
  assign regs_23_clock = clock; // @[:@151806.4]
  assign regs_23_reset = io_reset; // @[:@151807.4 RegFile.scala 76:16:@151814.4]
  assign regs_23_io_in = io_argOuts_20_bits; // @[RegFile.scala 75:16:@151813.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@151817.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@151811.4]
  assign regs_24_clock = clock; // @[:@151820.4]
  assign regs_24_reset = io_reset; // @[:@151821.4 RegFile.scala 76:16:@151828.4]
  assign regs_24_io_in = io_argOuts_21_bits; // @[RegFile.scala 75:16:@151827.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@151831.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@151825.4]
  assign regs_25_clock = clock; // @[:@151834.4]
  assign regs_25_reset = io_reset; // @[:@151835.4 RegFile.scala 76:16:@151842.4]
  assign regs_25_io_in = io_argOuts_22_bits; // @[RegFile.scala 75:16:@151841.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@151845.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@151839.4]
  assign regs_26_clock = clock; // @[:@151848.4]
  assign regs_26_reset = io_reset; // @[:@151849.4 RegFile.scala 76:16:@151856.4]
  assign regs_26_io_in = io_argOuts_23_bits; // @[RegFile.scala 75:16:@151855.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@151859.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@151853.4]
  assign regs_27_clock = clock; // @[:@151862.4]
  assign regs_27_reset = io_reset; // @[:@151863.4 RegFile.scala 76:16:@151870.4]
  assign regs_27_io_in = io_argOuts_24_bits; // @[RegFile.scala 75:16:@151869.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@151873.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@151867.4]
  assign regs_28_clock = clock; // @[:@151876.4]
  assign regs_28_reset = io_reset; // @[:@151877.4 RegFile.scala 76:16:@151884.4]
  assign regs_28_io_in = io_argOuts_25_bits; // @[RegFile.scala 75:16:@151883.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@151887.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@151881.4]
  assign regs_29_clock = clock; // @[:@151890.4]
  assign regs_29_reset = io_reset; // @[:@151891.4 RegFile.scala 76:16:@151898.4]
  assign regs_29_io_in = io_argOuts_26_bits; // @[RegFile.scala 75:16:@151897.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@151901.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@151895.4]
  assign regs_30_clock = clock; // @[:@151904.4]
  assign regs_30_reset = io_reset; // @[:@151905.4 RegFile.scala 76:16:@151912.4]
  assign regs_30_io_in = io_argOuts_27_bits; // @[RegFile.scala 75:16:@151911.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@151915.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@151909.4]
  assign regs_31_clock = clock; // @[:@151918.4]
  assign regs_31_reset = io_reset; // @[:@151919.4 RegFile.scala 76:16:@151926.4]
  assign regs_31_io_in = io_argOuts_28_bits; // @[RegFile.scala 75:16:@151925.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@151929.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@151923.4]
  assign regs_32_clock = clock; // @[:@151932.4]
  assign regs_32_reset = io_reset; // @[:@151933.4 RegFile.scala 76:16:@151940.4]
  assign regs_32_io_in = io_argOuts_29_bits; // @[RegFile.scala 75:16:@151939.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@151943.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@151937.4]
  assign regs_33_clock = clock; // @[:@151946.4]
  assign regs_33_reset = io_reset; // @[:@151947.4 RegFile.scala 76:16:@151954.4]
  assign regs_33_io_in = io_argOuts_30_bits; // @[RegFile.scala 75:16:@151953.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@151957.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@151951.4]
  assign regs_34_clock = clock; // @[:@151960.4]
  assign regs_34_reset = io_reset; // @[:@151961.4 RegFile.scala 76:16:@151968.4]
  assign regs_34_io_in = io_argOuts_31_bits; // @[RegFile.scala 75:16:@151967.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@151971.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@151965.4]
  assign regs_35_clock = clock; // @[:@151974.4]
  assign regs_35_reset = io_reset; // @[:@151975.4 RegFile.scala 76:16:@151982.4]
  assign regs_35_io_in = io_argOuts_32_bits; // @[RegFile.scala 75:16:@151981.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@151985.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@151979.4]
  assign regs_36_clock = clock; // @[:@151988.4]
  assign regs_36_reset = io_reset; // @[:@151989.4 RegFile.scala 76:16:@151996.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@151995.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@151999.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@151993.4]
  assign regs_37_clock = clock; // @[:@152002.4]
  assign regs_37_reset = io_reset; // @[:@152003.4 RegFile.scala 76:16:@152010.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@152009.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@152013.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@152007.4]
  assign regs_38_clock = clock; // @[:@152016.4]
  assign regs_38_reset = io_reset; // @[:@152017.4 RegFile.scala 76:16:@152024.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@152023.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@152027.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@152021.4]
  assign regs_39_clock = clock; // @[:@152030.4]
  assign regs_39_reset = io_reset; // @[:@152031.4 RegFile.scala 76:16:@152038.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@152037.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@152041.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@152035.4]
  assign regs_40_clock = clock; // @[:@152044.4]
  assign regs_40_reset = io_reset; // @[:@152045.4 RegFile.scala 76:16:@152052.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@152051.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@152055.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@152049.4]
  assign regs_41_clock = clock; // @[:@152058.4]
  assign regs_41_reset = io_reset; // @[:@152059.4 RegFile.scala 76:16:@152066.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@152065.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@152069.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@152063.4]
  assign regs_42_clock = clock; // @[:@152072.4]
  assign regs_42_reset = io_reset; // @[:@152073.4 RegFile.scala 76:16:@152080.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@152079.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@152083.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@152077.4]
  assign regs_43_clock = clock; // @[:@152086.4]
  assign regs_43_reset = io_reset; // @[:@152087.4 RegFile.scala 76:16:@152094.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@152093.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@152097.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@152091.4]
  assign regs_44_clock = clock; // @[:@152100.4]
  assign regs_44_reset = io_reset; // @[:@152101.4 RegFile.scala 76:16:@152108.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@152107.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@152111.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@152105.4]
  assign regs_45_clock = clock; // @[:@152114.4]
  assign regs_45_reset = io_reset; // @[:@152115.4 RegFile.scala 76:16:@152122.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@152121.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@152125.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@152119.4]
  assign regs_46_clock = clock; // @[:@152128.4]
  assign regs_46_reset = io_reset; // @[:@152129.4 RegFile.scala 76:16:@152136.4]
  assign regs_46_io_in = io_argOuts_43_bits; // @[RegFile.scala 75:16:@152135.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@152139.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@152133.4]
  assign regs_47_clock = clock; // @[:@152142.4]
  assign regs_47_reset = io_reset; // @[:@152143.4 RegFile.scala 76:16:@152150.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@152149.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@152153.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@152147.4]
  assign regs_48_clock = clock; // @[:@152156.4]
  assign regs_48_reset = io_reset; // @[:@152157.4 RegFile.scala 76:16:@152164.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@152163.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@152167.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@152161.4]
  assign regs_49_clock = clock; // @[:@152170.4]
  assign regs_49_reset = io_reset; // @[:@152171.4 RegFile.scala 76:16:@152178.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@152177.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@152181.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@152175.4]
  assign regs_50_clock = clock; // @[:@152184.4]
  assign regs_50_reset = io_reset; // @[:@152185.4 RegFile.scala 76:16:@152192.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@152191.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@152195.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@152189.4]
  assign regs_51_clock = clock; // @[:@152198.4]
  assign regs_51_reset = io_reset; // @[:@152199.4 RegFile.scala 76:16:@152206.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@152205.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@152209.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@152203.4]
  assign regs_52_clock = clock; // @[:@152212.4]
  assign regs_52_reset = io_reset; // @[:@152213.4 RegFile.scala 76:16:@152220.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@152219.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@152223.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@152217.4]
  assign regs_53_clock = clock; // @[:@152226.4]
  assign regs_53_reset = io_reset; // @[:@152227.4 RegFile.scala 76:16:@152234.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@152233.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@152237.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@152231.4]
  assign regs_54_clock = clock; // @[:@152240.4]
  assign regs_54_reset = io_reset; // @[:@152241.4 RegFile.scala 76:16:@152248.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@152247.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@152251.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@152245.4]
  assign regs_55_clock = clock; // @[:@152254.4]
  assign regs_55_reset = io_reset; // @[:@152255.4 RegFile.scala 76:16:@152262.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@152261.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@152265.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@152259.4]
  assign regs_56_clock = clock; // @[:@152268.4]
  assign regs_56_reset = io_reset; // @[:@152269.4 RegFile.scala 76:16:@152276.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@152275.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@152279.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@152273.4]
  assign regs_57_clock = clock; // @[:@152282.4]
  assign regs_57_reset = io_reset; // @[:@152283.4 RegFile.scala 76:16:@152290.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@152289.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@152293.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@152287.4]
  assign regs_58_clock = clock; // @[:@152296.4]
  assign regs_58_reset = io_reset; // @[:@152297.4 RegFile.scala 76:16:@152304.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@152303.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@152307.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@152301.4]
  assign regs_59_clock = clock; // @[:@152310.4]
  assign regs_59_reset = io_reset; // @[:@152311.4 RegFile.scala 76:16:@152318.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@152317.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@152321.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@152315.4]
  assign regs_60_clock = clock; // @[:@152324.4]
  assign regs_60_reset = io_reset; // @[:@152325.4 RegFile.scala 76:16:@152332.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@152331.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@152335.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@152329.4]
  assign regs_61_clock = clock; // @[:@152338.4]
  assign regs_61_reset = io_reset; // @[:@152339.4 RegFile.scala 76:16:@152346.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@152345.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@152349.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@152343.4]
  assign regs_62_clock = clock; // @[:@152352.4]
  assign regs_62_reset = io_reset; // @[:@152353.4 RegFile.scala 76:16:@152360.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@152359.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@152363.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@152357.4]
  assign regs_63_clock = clock; // @[:@152366.4]
  assign regs_63_reset = io_reset; // @[:@152367.4 RegFile.scala 76:16:@152374.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@152373.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@152377.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@152371.4]
  assign regs_64_clock = clock; // @[:@152380.4]
  assign regs_64_reset = io_reset; // @[:@152381.4 RegFile.scala 76:16:@152388.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@152387.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@152391.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@152385.4]
  assign regs_65_clock = clock; // @[:@152394.4]
  assign regs_65_reset = io_reset; // @[:@152395.4 RegFile.scala 76:16:@152402.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@152401.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@152405.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@152399.4]
  assign regs_66_clock = clock; // @[:@152408.4]
  assign regs_66_reset = io_reset; // @[:@152409.4 RegFile.scala 76:16:@152416.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@152415.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@152419.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@152413.4]
  assign regs_67_clock = clock; // @[:@152422.4]
  assign regs_67_reset = io_reset; // @[:@152423.4 RegFile.scala 76:16:@152430.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@152429.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@152433.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@152427.4]
  assign regs_68_clock = clock; // @[:@152436.4]
  assign regs_68_reset = io_reset; // @[:@152437.4 RegFile.scala 76:16:@152444.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@152443.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@152447.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@152441.4]
  assign regs_69_clock = clock; // @[:@152450.4]
  assign regs_69_reset = io_reset; // @[:@152451.4 RegFile.scala 76:16:@152458.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@152457.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@152461.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@152455.4]
  assign regs_70_clock = clock; // @[:@152464.4]
  assign regs_70_reset = io_reset; // @[:@152465.4 RegFile.scala 76:16:@152472.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@152471.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@152475.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@152469.4]
  assign regs_71_clock = clock; // @[:@152478.4]
  assign regs_71_reset = io_reset; // @[:@152479.4 RegFile.scala 76:16:@152486.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@152485.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@152489.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@152483.4]
  assign regs_72_clock = clock; // @[:@152492.4]
  assign regs_72_reset = io_reset; // @[:@152493.4 RegFile.scala 76:16:@152500.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@152499.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@152503.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@152497.4]
  assign regs_73_clock = clock; // @[:@152506.4]
  assign regs_73_reset = io_reset; // @[:@152507.4 RegFile.scala 76:16:@152514.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@152513.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@152517.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@152511.4]
  assign regs_74_clock = clock; // @[:@152520.4]
  assign regs_74_reset = io_reset; // @[:@152521.4 RegFile.scala 76:16:@152528.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@152527.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@152531.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@152525.4]
  assign regs_75_clock = clock; // @[:@152534.4]
  assign regs_75_reset = io_reset; // @[:@152535.4 RegFile.scala 76:16:@152542.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@152541.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@152545.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@152539.4]
  assign regs_76_clock = clock; // @[:@152548.4]
  assign regs_76_reset = io_reset; // @[:@152549.4 RegFile.scala 76:16:@152556.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@152555.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@152559.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@152553.4]
  assign regs_77_clock = clock; // @[:@152562.4]
  assign regs_77_reset = io_reset; // @[:@152563.4 RegFile.scala 76:16:@152570.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@152569.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@152573.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@152567.4]
  assign regs_78_clock = clock; // @[:@152576.4]
  assign regs_78_reset = io_reset; // @[:@152577.4 RegFile.scala 76:16:@152584.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@152583.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@152587.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@152581.4]
  assign regs_79_clock = clock; // @[:@152590.4]
  assign regs_79_reset = io_reset; // @[:@152591.4 RegFile.scala 76:16:@152598.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@152597.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@152601.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@152595.4]
  assign regs_80_clock = clock; // @[:@152604.4]
  assign regs_80_reset = io_reset; // @[:@152605.4 RegFile.scala 76:16:@152612.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@152611.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@152615.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@152609.4]
  assign regs_81_clock = clock; // @[:@152618.4]
  assign regs_81_reset = io_reset; // @[:@152619.4 RegFile.scala 76:16:@152626.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@152625.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@152629.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@152623.4]
  assign regs_82_clock = clock; // @[:@152632.4]
  assign regs_82_reset = io_reset; // @[:@152633.4 RegFile.scala 76:16:@152640.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@152639.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@152643.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@152637.4]
  assign regs_83_clock = clock; // @[:@152646.4]
  assign regs_83_reset = io_reset; // @[:@152647.4 RegFile.scala 76:16:@152654.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@152653.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@152657.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@152651.4]
  assign regs_84_clock = clock; // @[:@152660.4]
  assign regs_84_reset = io_reset; // @[:@152661.4 RegFile.scala 76:16:@152668.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@152667.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@152671.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@152665.4]
  assign regs_85_clock = clock; // @[:@152674.4]
  assign regs_85_reset = io_reset; // @[:@152675.4 RegFile.scala 76:16:@152682.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@152681.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@152685.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@152679.4]
  assign regs_86_clock = clock; // @[:@152688.4]
  assign regs_86_reset = io_reset; // @[:@152689.4 RegFile.scala 76:16:@152696.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@152695.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@152699.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@152693.4]
  assign regs_87_clock = clock; // @[:@152702.4]
  assign regs_87_reset = io_reset; // @[:@152703.4 RegFile.scala 76:16:@152710.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@152709.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@152713.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@152707.4]
  assign regs_88_clock = clock; // @[:@152716.4]
  assign regs_88_reset = io_reset; // @[:@152717.4 RegFile.scala 76:16:@152724.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@152723.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@152727.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@152721.4]
  assign regs_89_clock = clock; // @[:@152730.4]
  assign regs_89_reset = io_reset; // @[:@152731.4 RegFile.scala 76:16:@152738.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@152737.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@152741.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@152735.4]
  assign regs_90_clock = clock; // @[:@152744.4]
  assign regs_90_reset = io_reset; // @[:@152745.4 RegFile.scala 76:16:@152752.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@152751.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@152755.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@152749.4]
  assign regs_91_clock = clock; // @[:@152758.4]
  assign regs_91_reset = io_reset; // @[:@152759.4 RegFile.scala 76:16:@152766.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@152765.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@152769.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@152763.4]
  assign regs_92_clock = clock; // @[:@152772.4]
  assign regs_92_reset = io_reset; // @[:@152773.4 RegFile.scala 76:16:@152780.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@152779.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@152783.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@152777.4]
  assign regs_93_clock = clock; // @[:@152786.4]
  assign regs_93_reset = io_reset; // @[:@152787.4 RegFile.scala 76:16:@152794.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@152793.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@152797.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@152791.4]
  assign regs_94_clock = clock; // @[:@152800.4]
  assign regs_94_reset = io_reset; // @[:@152801.4 RegFile.scala 76:16:@152808.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@152807.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@152811.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@152805.4]
  assign regs_95_clock = clock; // @[:@152814.4]
  assign regs_95_reset = io_reset; // @[:@152815.4 RegFile.scala 76:16:@152822.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@152821.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@152825.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@152819.4]
  assign regs_96_clock = clock; // @[:@152828.4]
  assign regs_96_reset = io_reset; // @[:@152829.4 RegFile.scala 76:16:@152836.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@152835.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@152839.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@152833.4]
  assign regs_97_clock = clock; // @[:@152842.4]
  assign regs_97_reset = io_reset; // @[:@152843.4 RegFile.scala 76:16:@152850.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@152849.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@152853.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@152847.4]
  assign regs_98_clock = clock; // @[:@152856.4]
  assign regs_98_reset = io_reset; // @[:@152857.4 RegFile.scala 76:16:@152864.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@152863.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@152867.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@152861.4]
  assign regs_99_clock = clock; // @[:@152870.4]
  assign regs_99_reset = io_reset; // @[:@152871.4 RegFile.scala 76:16:@152878.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@152877.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@152881.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@152875.4]
  assign regs_100_clock = clock; // @[:@152884.4]
  assign regs_100_reset = io_reset; // @[:@152885.4 RegFile.scala 76:16:@152892.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@152891.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@152895.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@152889.4]
  assign regs_101_clock = clock; // @[:@152898.4]
  assign regs_101_reset = io_reset; // @[:@152899.4 RegFile.scala 76:16:@152906.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@152905.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@152909.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@152903.4]
  assign regs_102_clock = clock; // @[:@152912.4]
  assign regs_102_reset = io_reset; // @[:@152913.4 RegFile.scala 76:16:@152920.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@152919.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@152923.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@152917.4]
  assign regs_103_clock = clock; // @[:@152926.4]
  assign regs_103_reset = io_reset; // @[:@152927.4 RegFile.scala 76:16:@152934.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@152933.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@152937.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@152931.4]
  assign regs_104_clock = clock; // @[:@152940.4]
  assign regs_104_reset = io_reset; // @[:@152941.4 RegFile.scala 76:16:@152948.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@152947.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@152951.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@152945.4]
  assign regs_105_clock = clock; // @[:@152954.4]
  assign regs_105_reset = io_reset; // @[:@152955.4 RegFile.scala 76:16:@152962.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@152961.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@152965.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@152959.4]
  assign regs_106_clock = clock; // @[:@152968.4]
  assign regs_106_reset = io_reset; // @[:@152969.4 RegFile.scala 76:16:@152976.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@152975.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@152979.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@152973.4]
  assign regs_107_clock = clock; // @[:@152982.4]
  assign regs_107_reset = io_reset; // @[:@152983.4 RegFile.scala 76:16:@152990.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@152989.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@152993.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@152987.4]
  assign regs_108_clock = clock; // @[:@152996.4]
  assign regs_108_reset = io_reset; // @[:@152997.4 RegFile.scala 76:16:@153004.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@153003.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@153007.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@153001.4]
  assign regs_109_clock = clock; // @[:@153010.4]
  assign regs_109_reset = io_reset; // @[:@153011.4 RegFile.scala 76:16:@153018.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@153017.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@153021.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@153015.4]
  assign regs_110_clock = clock; // @[:@153024.4]
  assign regs_110_reset = io_reset; // @[:@153025.4 RegFile.scala 76:16:@153032.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@153031.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@153035.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@153029.4]
  assign regs_111_clock = clock; // @[:@153038.4]
  assign regs_111_reset = io_reset; // @[:@153039.4 RegFile.scala 76:16:@153046.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@153045.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@153049.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@153043.4]
  assign regs_112_clock = clock; // @[:@153052.4]
  assign regs_112_reset = io_reset; // @[:@153053.4 RegFile.scala 76:16:@153060.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@153059.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@153063.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@153057.4]
  assign regs_113_clock = clock; // @[:@153066.4]
  assign regs_113_reset = io_reset; // @[:@153067.4 RegFile.scala 76:16:@153074.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@153073.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@153077.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@153071.4]
  assign regs_114_clock = clock; // @[:@153080.4]
  assign regs_114_reset = io_reset; // @[:@153081.4 RegFile.scala 76:16:@153088.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@153087.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@153091.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@153085.4]
  assign regs_115_clock = clock; // @[:@153094.4]
  assign regs_115_reset = io_reset; // @[:@153095.4 RegFile.scala 76:16:@153102.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@153101.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@153105.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@153099.4]
  assign regs_116_clock = clock; // @[:@153108.4]
  assign regs_116_reset = io_reset; // @[:@153109.4 RegFile.scala 76:16:@153116.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@153115.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@153119.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@153113.4]
  assign regs_117_clock = clock; // @[:@153122.4]
  assign regs_117_reset = io_reset; // @[:@153123.4 RegFile.scala 76:16:@153130.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@153129.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@153133.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@153127.4]
  assign regs_118_clock = clock; // @[:@153136.4]
  assign regs_118_reset = io_reset; // @[:@153137.4 RegFile.scala 76:16:@153144.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@153143.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@153147.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@153141.4]
  assign regs_119_clock = clock; // @[:@153150.4]
  assign regs_119_reset = io_reset; // @[:@153151.4 RegFile.scala 76:16:@153158.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@153157.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@153161.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@153155.4]
  assign regs_120_clock = clock; // @[:@153164.4]
  assign regs_120_reset = io_reset; // @[:@153165.4 RegFile.scala 76:16:@153172.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@153171.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@153175.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@153169.4]
  assign regs_121_clock = clock; // @[:@153178.4]
  assign regs_121_reset = io_reset; // @[:@153179.4 RegFile.scala 76:16:@153186.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@153185.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@153189.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@153183.4]
  assign regs_122_clock = clock; // @[:@153192.4]
  assign regs_122_reset = io_reset; // @[:@153193.4 RegFile.scala 76:16:@153200.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@153199.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@153203.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@153197.4]
  assign regs_123_clock = clock; // @[:@153206.4]
  assign regs_123_reset = io_reset; // @[:@153207.4 RegFile.scala 76:16:@153214.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@153213.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@153217.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@153211.4]
  assign regs_124_clock = clock; // @[:@153220.4]
  assign regs_124_reset = io_reset; // @[:@153221.4 RegFile.scala 76:16:@153228.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@153227.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@153231.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@153225.4]
  assign regs_125_clock = clock; // @[:@153234.4]
  assign regs_125_reset = io_reset; // @[:@153235.4 RegFile.scala 76:16:@153242.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@153241.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@153245.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@153239.4]
  assign regs_126_clock = clock; // @[:@153248.4]
  assign regs_126_reset = io_reset; // @[:@153249.4 RegFile.scala 76:16:@153256.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@153255.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@153259.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@153253.4]
  assign regs_127_clock = clock; // @[:@153262.4]
  assign regs_127_reset = io_reset; // @[:@153263.4 RegFile.scala 76:16:@153270.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@153269.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@153273.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@153267.4]
  assign regs_128_clock = clock; // @[:@153276.4]
  assign regs_128_reset = io_reset; // @[:@153277.4 RegFile.scala 76:16:@153284.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@153283.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@153287.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@153281.4]
  assign regs_129_clock = clock; // @[:@153290.4]
  assign regs_129_reset = io_reset; // @[:@153291.4 RegFile.scala 76:16:@153298.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@153297.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@153301.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@153295.4]
  assign regs_130_clock = clock; // @[:@153304.4]
  assign regs_130_reset = io_reset; // @[:@153305.4 RegFile.scala 76:16:@153312.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@153311.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@153315.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@153309.4]
  assign regs_131_clock = clock; // @[:@153318.4]
  assign regs_131_reset = io_reset; // @[:@153319.4 RegFile.scala 76:16:@153326.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@153325.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@153329.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@153323.4]
  assign regs_132_clock = clock; // @[:@153332.4]
  assign regs_132_reset = io_reset; // @[:@153333.4 RegFile.scala 76:16:@153340.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@153339.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@153343.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@153337.4]
  assign regs_133_clock = clock; // @[:@153346.4]
  assign regs_133_reset = io_reset; // @[:@153347.4 RegFile.scala 76:16:@153354.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@153353.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@153357.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@153351.4]
  assign regs_134_clock = clock; // @[:@153360.4]
  assign regs_134_reset = io_reset; // @[:@153361.4 RegFile.scala 76:16:@153368.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@153367.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@153371.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@153365.4]
  assign regs_135_clock = clock; // @[:@153374.4]
  assign regs_135_reset = io_reset; // @[:@153375.4 RegFile.scala 76:16:@153382.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@153381.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@153385.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@153379.4]
  assign regs_136_clock = clock; // @[:@153388.4]
  assign regs_136_reset = io_reset; // @[:@153389.4 RegFile.scala 76:16:@153396.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@153395.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@153399.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@153393.4]
  assign regs_137_clock = clock; // @[:@153402.4]
  assign regs_137_reset = io_reset; // @[:@153403.4 RegFile.scala 76:16:@153410.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@153409.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@153413.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@153407.4]
  assign regs_138_clock = clock; // @[:@153416.4]
  assign regs_138_reset = io_reset; // @[:@153417.4 RegFile.scala 76:16:@153424.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@153423.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@153427.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@153421.4]
  assign regs_139_clock = clock; // @[:@153430.4]
  assign regs_139_reset = io_reset; // @[:@153431.4 RegFile.scala 76:16:@153438.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@153437.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@153441.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@153435.4]
  assign regs_140_clock = clock; // @[:@153444.4]
  assign regs_140_reset = io_reset; // @[:@153445.4 RegFile.scala 76:16:@153452.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@153451.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@153455.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@153449.4]
  assign regs_141_clock = clock; // @[:@153458.4]
  assign regs_141_reset = io_reset; // @[:@153459.4 RegFile.scala 76:16:@153466.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@153465.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@153469.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@153463.4]
  assign regs_142_clock = clock; // @[:@153472.4]
  assign regs_142_reset = io_reset; // @[:@153473.4 RegFile.scala 76:16:@153480.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@153479.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@153483.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@153477.4]
  assign regs_143_clock = clock; // @[:@153486.4]
  assign regs_143_reset = io_reset; // @[:@153487.4 RegFile.scala 76:16:@153494.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@153493.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@153497.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@153491.4]
  assign regs_144_clock = clock; // @[:@153500.4]
  assign regs_144_reset = io_reset; // @[:@153501.4 RegFile.scala 76:16:@153508.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@153507.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@153511.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@153505.4]
  assign regs_145_clock = clock; // @[:@153514.4]
  assign regs_145_reset = io_reset; // @[:@153515.4 RegFile.scala 76:16:@153522.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@153521.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@153525.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@153519.4]
  assign regs_146_clock = clock; // @[:@153528.4]
  assign regs_146_reset = io_reset; // @[:@153529.4 RegFile.scala 76:16:@153536.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@153535.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@153539.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@153533.4]
  assign regs_147_clock = clock; // @[:@153542.4]
  assign regs_147_reset = io_reset; // @[:@153543.4 RegFile.scala 76:16:@153550.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@153549.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@153553.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@153547.4]
  assign regs_148_clock = clock; // @[:@153556.4]
  assign regs_148_reset = io_reset; // @[:@153557.4 RegFile.scala 76:16:@153564.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@153563.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@153567.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@153561.4]
  assign regs_149_clock = clock; // @[:@153570.4]
  assign regs_149_reset = io_reset; // @[:@153571.4 RegFile.scala 76:16:@153578.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@153577.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@153581.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@153575.4]
  assign regs_150_clock = clock; // @[:@153584.4]
  assign regs_150_reset = io_reset; // @[:@153585.4 RegFile.scala 76:16:@153592.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@153591.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@153595.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@153589.4]
  assign regs_151_clock = clock; // @[:@153598.4]
  assign regs_151_reset = io_reset; // @[:@153599.4 RegFile.scala 76:16:@153606.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@153605.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@153609.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@153603.4]
  assign regs_152_clock = clock; // @[:@153612.4]
  assign regs_152_reset = io_reset; // @[:@153613.4 RegFile.scala 76:16:@153620.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@153619.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@153623.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@153617.4]
  assign regs_153_clock = clock; // @[:@153626.4]
  assign regs_153_reset = io_reset; // @[:@153627.4 RegFile.scala 76:16:@153634.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@153633.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@153637.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@153631.4]
  assign regs_154_clock = clock; // @[:@153640.4]
  assign regs_154_reset = io_reset; // @[:@153641.4 RegFile.scala 76:16:@153648.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@153647.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@153651.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@153645.4]
  assign regs_155_clock = clock; // @[:@153654.4]
  assign regs_155_reset = io_reset; // @[:@153655.4 RegFile.scala 76:16:@153662.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@153661.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@153665.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@153659.4]
  assign regs_156_clock = clock; // @[:@153668.4]
  assign regs_156_reset = io_reset; // @[:@153669.4 RegFile.scala 76:16:@153676.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@153675.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@153679.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@153673.4]
  assign regs_157_clock = clock; // @[:@153682.4]
  assign regs_157_reset = io_reset; // @[:@153683.4 RegFile.scala 76:16:@153690.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@153689.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@153693.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@153687.4]
  assign regs_158_clock = clock; // @[:@153696.4]
  assign regs_158_reset = io_reset; // @[:@153697.4 RegFile.scala 76:16:@153704.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@153703.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@153707.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@153701.4]
  assign regs_159_clock = clock; // @[:@153710.4]
  assign regs_159_reset = io_reset; // @[:@153711.4 RegFile.scala 76:16:@153718.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@153717.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@153721.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@153715.4]
  assign regs_160_clock = clock; // @[:@153724.4]
  assign regs_160_reset = io_reset; // @[:@153725.4 RegFile.scala 76:16:@153732.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@153731.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@153735.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@153729.4]
  assign regs_161_clock = clock; // @[:@153738.4]
  assign regs_161_reset = io_reset; // @[:@153739.4 RegFile.scala 76:16:@153746.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@153745.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@153749.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@153743.4]
  assign regs_162_clock = clock; // @[:@153752.4]
  assign regs_162_reset = io_reset; // @[:@153753.4 RegFile.scala 76:16:@153760.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@153759.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@153763.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@153757.4]
  assign regs_163_clock = clock; // @[:@153766.4]
  assign regs_163_reset = io_reset; // @[:@153767.4 RegFile.scala 76:16:@153774.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@153773.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@153777.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@153771.4]
  assign regs_164_clock = clock; // @[:@153780.4]
  assign regs_164_reset = io_reset; // @[:@153781.4 RegFile.scala 76:16:@153788.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@153787.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@153791.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@153785.4]
  assign regs_165_clock = clock; // @[:@153794.4]
  assign regs_165_reset = io_reset; // @[:@153795.4 RegFile.scala 76:16:@153802.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@153801.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@153805.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@153799.4]
  assign regs_166_clock = clock; // @[:@153808.4]
  assign regs_166_reset = io_reset; // @[:@153809.4 RegFile.scala 76:16:@153816.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@153815.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@153819.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@153813.4]
  assign regs_167_clock = clock; // @[:@153822.4]
  assign regs_167_reset = io_reset; // @[:@153823.4 RegFile.scala 76:16:@153830.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@153829.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@153833.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@153827.4]
  assign regs_168_clock = clock; // @[:@153836.4]
  assign regs_168_reset = io_reset; // @[:@153837.4 RegFile.scala 76:16:@153844.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@153843.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@153847.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@153841.4]
  assign regs_169_clock = clock; // @[:@153850.4]
  assign regs_169_reset = io_reset; // @[:@153851.4 RegFile.scala 76:16:@153858.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@153857.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@153861.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@153855.4]
  assign regs_170_clock = clock; // @[:@153864.4]
  assign regs_170_reset = io_reset; // @[:@153865.4 RegFile.scala 76:16:@153872.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@153871.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@153875.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@153869.4]
  assign regs_171_clock = clock; // @[:@153878.4]
  assign regs_171_reset = io_reset; // @[:@153879.4 RegFile.scala 76:16:@153886.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@153885.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@153889.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@153883.4]
  assign regs_172_clock = clock; // @[:@153892.4]
  assign regs_172_reset = io_reset; // @[:@153893.4 RegFile.scala 76:16:@153900.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@153899.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@153903.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@153897.4]
  assign regs_173_clock = clock; // @[:@153906.4]
  assign regs_173_reset = io_reset; // @[:@153907.4 RegFile.scala 76:16:@153914.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@153913.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@153917.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@153911.4]
  assign regs_174_clock = clock; // @[:@153920.4]
  assign regs_174_reset = io_reset; // @[:@153921.4 RegFile.scala 76:16:@153928.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@153927.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@153931.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@153925.4]
  assign regs_175_clock = clock; // @[:@153934.4]
  assign regs_175_reset = io_reset; // @[:@153935.4 RegFile.scala 76:16:@153942.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@153941.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@153945.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@153939.4]
  assign regs_176_clock = clock; // @[:@153948.4]
  assign regs_176_reset = io_reset; // @[:@153949.4 RegFile.scala 76:16:@153956.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@153955.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@153959.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@153953.4]
  assign regs_177_clock = clock; // @[:@153962.4]
  assign regs_177_reset = io_reset; // @[:@153963.4 RegFile.scala 76:16:@153970.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@153969.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@153973.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@153967.4]
  assign regs_178_clock = clock; // @[:@153976.4]
  assign regs_178_reset = io_reset; // @[:@153977.4 RegFile.scala 76:16:@153984.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@153983.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@153987.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@153981.4]
  assign regs_179_clock = clock; // @[:@153990.4]
  assign regs_179_reset = io_reset; // @[:@153991.4 RegFile.scala 76:16:@153998.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@153997.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@154001.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@153995.4]
  assign regs_180_clock = clock; // @[:@154004.4]
  assign regs_180_reset = io_reset; // @[:@154005.4 RegFile.scala 76:16:@154012.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@154011.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@154015.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@154009.4]
  assign regs_181_clock = clock; // @[:@154018.4]
  assign regs_181_reset = io_reset; // @[:@154019.4 RegFile.scala 76:16:@154026.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@154025.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@154029.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@154023.4]
  assign regs_182_clock = clock; // @[:@154032.4]
  assign regs_182_reset = io_reset; // @[:@154033.4 RegFile.scala 76:16:@154040.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@154039.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@154043.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@154037.4]
  assign regs_183_clock = clock; // @[:@154046.4]
  assign regs_183_reset = io_reset; // @[:@154047.4 RegFile.scala 76:16:@154054.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@154053.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@154057.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@154051.4]
  assign regs_184_clock = clock; // @[:@154060.4]
  assign regs_184_reset = io_reset; // @[:@154061.4 RegFile.scala 76:16:@154068.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@154067.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@154071.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@154065.4]
  assign regs_185_clock = clock; // @[:@154074.4]
  assign regs_185_reset = io_reset; // @[:@154075.4 RegFile.scala 76:16:@154082.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@154081.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@154085.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@154079.4]
  assign regs_186_clock = clock; // @[:@154088.4]
  assign regs_186_reset = io_reset; // @[:@154089.4 RegFile.scala 76:16:@154096.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@154095.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@154099.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@154093.4]
  assign regs_187_clock = clock; // @[:@154102.4]
  assign regs_187_reset = io_reset; // @[:@154103.4 RegFile.scala 76:16:@154110.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@154109.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@154113.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@154107.4]
  assign regs_188_clock = clock; // @[:@154116.4]
  assign regs_188_reset = io_reset; // @[:@154117.4 RegFile.scala 76:16:@154124.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@154123.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@154127.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@154121.4]
  assign regs_189_clock = clock; // @[:@154130.4]
  assign regs_189_reset = io_reset; // @[:@154131.4 RegFile.scala 76:16:@154138.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@154137.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@154141.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@154135.4]
  assign regs_190_clock = clock; // @[:@154144.4]
  assign regs_190_reset = io_reset; // @[:@154145.4 RegFile.scala 76:16:@154152.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@154151.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@154155.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@154149.4]
  assign regs_191_clock = clock; // @[:@154158.4]
  assign regs_191_reset = io_reset; // @[:@154159.4 RegFile.scala 76:16:@154166.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@154165.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@154169.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@154163.4]
  assign regs_192_clock = clock; // @[:@154172.4]
  assign regs_192_reset = io_reset; // @[:@154173.4 RegFile.scala 76:16:@154180.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@154179.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@154183.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@154177.4]
  assign regs_193_clock = clock; // @[:@154186.4]
  assign regs_193_reset = io_reset; // @[:@154187.4 RegFile.scala 76:16:@154194.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@154193.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@154197.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@154191.4]
  assign regs_194_clock = clock; // @[:@154200.4]
  assign regs_194_reset = io_reset; // @[:@154201.4 RegFile.scala 76:16:@154208.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@154207.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@154211.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@154205.4]
  assign regs_195_clock = clock; // @[:@154214.4]
  assign regs_195_reset = io_reset; // @[:@154215.4 RegFile.scala 76:16:@154222.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@154221.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@154225.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@154219.4]
  assign regs_196_clock = clock; // @[:@154228.4]
  assign regs_196_reset = io_reset; // @[:@154229.4 RegFile.scala 76:16:@154236.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@154235.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@154239.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@154233.4]
  assign regs_197_clock = clock; // @[:@154242.4]
  assign regs_197_reset = io_reset; // @[:@154243.4 RegFile.scala 76:16:@154250.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@154249.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@154253.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@154247.4]
  assign regs_198_clock = clock; // @[:@154256.4]
  assign regs_198_reset = io_reset; // @[:@154257.4 RegFile.scala 76:16:@154264.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@154263.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@154267.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@154261.4]
  assign regs_199_clock = clock; // @[:@154270.4]
  assign regs_199_reset = io_reset; // @[:@154271.4 RegFile.scala 76:16:@154278.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@154277.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@154281.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@154275.4]
  assign regs_200_clock = clock; // @[:@154284.4]
  assign regs_200_reset = io_reset; // @[:@154285.4 RegFile.scala 76:16:@154292.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@154291.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@154295.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@154289.4]
  assign regs_201_clock = clock; // @[:@154298.4]
  assign regs_201_reset = io_reset; // @[:@154299.4 RegFile.scala 76:16:@154306.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@154305.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@154309.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@154303.4]
  assign regs_202_clock = clock; // @[:@154312.4]
  assign regs_202_reset = io_reset; // @[:@154313.4 RegFile.scala 76:16:@154320.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@154319.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@154323.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@154317.4]
  assign regs_203_clock = clock; // @[:@154326.4]
  assign regs_203_reset = io_reset; // @[:@154327.4 RegFile.scala 76:16:@154334.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@154333.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@154337.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@154331.4]
  assign regs_204_clock = clock; // @[:@154340.4]
  assign regs_204_reset = io_reset; // @[:@154341.4 RegFile.scala 76:16:@154348.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@154347.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@154351.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@154345.4]
  assign regs_205_clock = clock; // @[:@154354.4]
  assign regs_205_reset = io_reset; // @[:@154355.4 RegFile.scala 76:16:@154362.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@154361.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@154365.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@154359.4]
  assign regs_206_clock = clock; // @[:@154368.4]
  assign regs_206_reset = io_reset; // @[:@154369.4 RegFile.scala 76:16:@154376.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@154375.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@154379.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@154373.4]
  assign regs_207_clock = clock; // @[:@154382.4]
  assign regs_207_reset = io_reset; // @[:@154383.4 RegFile.scala 76:16:@154390.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@154389.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@154393.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@154387.4]
  assign regs_208_clock = clock; // @[:@154396.4]
  assign regs_208_reset = io_reset; // @[:@154397.4 RegFile.scala 76:16:@154404.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@154403.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@154407.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@154401.4]
  assign regs_209_clock = clock; // @[:@154410.4]
  assign regs_209_reset = io_reset; // @[:@154411.4 RegFile.scala 76:16:@154418.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@154417.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@154421.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@154415.4]
  assign regs_210_clock = clock; // @[:@154424.4]
  assign regs_210_reset = io_reset; // @[:@154425.4 RegFile.scala 76:16:@154432.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@154431.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@154435.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@154429.4]
  assign regs_211_clock = clock; // @[:@154438.4]
  assign regs_211_reset = io_reset; // @[:@154439.4 RegFile.scala 76:16:@154446.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@154445.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@154449.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@154443.4]
  assign regs_212_clock = clock; // @[:@154452.4]
  assign regs_212_reset = io_reset; // @[:@154453.4 RegFile.scala 76:16:@154460.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@154459.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@154463.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@154457.4]
  assign regs_213_clock = clock; // @[:@154466.4]
  assign regs_213_reset = io_reset; // @[:@154467.4 RegFile.scala 76:16:@154474.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@154473.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@154477.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@154471.4]
  assign regs_214_clock = clock; // @[:@154480.4]
  assign regs_214_reset = io_reset; // @[:@154481.4 RegFile.scala 76:16:@154488.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@154487.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@154491.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@154485.4]
  assign regs_215_clock = clock; // @[:@154494.4]
  assign regs_215_reset = io_reset; // @[:@154495.4 RegFile.scala 76:16:@154502.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@154501.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@154505.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@154499.4]
  assign regs_216_clock = clock; // @[:@154508.4]
  assign regs_216_reset = io_reset; // @[:@154509.4 RegFile.scala 76:16:@154516.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@154515.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@154519.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@154513.4]
  assign regs_217_clock = clock; // @[:@154522.4]
  assign regs_217_reset = io_reset; // @[:@154523.4 RegFile.scala 76:16:@154530.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@154529.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@154533.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@154527.4]
  assign regs_218_clock = clock; // @[:@154536.4]
  assign regs_218_reset = io_reset; // @[:@154537.4 RegFile.scala 76:16:@154544.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@154543.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@154547.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@154541.4]
  assign regs_219_clock = clock; // @[:@154550.4]
  assign regs_219_reset = io_reset; // @[:@154551.4 RegFile.scala 76:16:@154558.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@154557.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@154561.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@154555.4]
  assign regs_220_clock = clock; // @[:@154564.4]
  assign regs_220_reset = io_reset; // @[:@154565.4 RegFile.scala 76:16:@154572.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@154571.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@154575.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@154569.4]
  assign regs_221_clock = clock; // @[:@154578.4]
  assign regs_221_reset = io_reset; // @[:@154579.4 RegFile.scala 76:16:@154586.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@154585.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@154589.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@154583.4]
  assign regs_222_clock = clock; // @[:@154592.4]
  assign regs_222_reset = io_reset; // @[:@154593.4 RegFile.scala 76:16:@154600.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@154599.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@154603.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@154597.4]
  assign regs_223_clock = clock; // @[:@154606.4]
  assign regs_223_reset = io_reset; // @[:@154607.4 RegFile.scala 76:16:@154614.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@154613.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@154617.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@154611.4]
  assign regs_224_clock = clock; // @[:@154620.4]
  assign regs_224_reset = io_reset; // @[:@154621.4 RegFile.scala 76:16:@154628.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@154627.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@154631.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@154625.4]
  assign regs_225_clock = clock; // @[:@154634.4]
  assign regs_225_reset = io_reset; // @[:@154635.4 RegFile.scala 76:16:@154642.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@154641.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@154645.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@154639.4]
  assign regs_226_clock = clock; // @[:@154648.4]
  assign regs_226_reset = io_reset; // @[:@154649.4 RegFile.scala 76:16:@154656.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@154655.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@154659.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@154653.4]
  assign regs_227_clock = clock; // @[:@154662.4]
  assign regs_227_reset = io_reset; // @[:@154663.4 RegFile.scala 76:16:@154670.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@154669.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@154673.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@154667.4]
  assign regs_228_clock = clock; // @[:@154676.4]
  assign regs_228_reset = io_reset; // @[:@154677.4 RegFile.scala 76:16:@154684.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@154683.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@154687.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@154681.4]
  assign regs_229_clock = clock; // @[:@154690.4]
  assign regs_229_reset = io_reset; // @[:@154691.4 RegFile.scala 76:16:@154698.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@154697.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@154701.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@154695.4]
  assign regs_230_clock = clock; // @[:@154704.4]
  assign regs_230_reset = io_reset; // @[:@154705.4 RegFile.scala 76:16:@154712.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@154711.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@154715.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@154709.4]
  assign regs_231_clock = clock; // @[:@154718.4]
  assign regs_231_reset = io_reset; // @[:@154719.4 RegFile.scala 76:16:@154726.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@154725.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@154729.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@154723.4]
  assign regs_232_clock = clock; // @[:@154732.4]
  assign regs_232_reset = io_reset; // @[:@154733.4 RegFile.scala 76:16:@154740.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@154739.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@154743.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@154737.4]
  assign regs_233_clock = clock; // @[:@154746.4]
  assign regs_233_reset = io_reset; // @[:@154747.4 RegFile.scala 76:16:@154754.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@154753.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@154757.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@154751.4]
  assign regs_234_clock = clock; // @[:@154760.4]
  assign regs_234_reset = io_reset; // @[:@154761.4 RegFile.scala 76:16:@154768.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@154767.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@154771.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@154765.4]
  assign regs_235_clock = clock; // @[:@154774.4]
  assign regs_235_reset = io_reset; // @[:@154775.4 RegFile.scala 76:16:@154782.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@154781.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@154785.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@154779.4]
  assign regs_236_clock = clock; // @[:@154788.4]
  assign regs_236_reset = io_reset; // @[:@154789.4 RegFile.scala 76:16:@154796.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@154795.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@154799.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@154793.4]
  assign regs_237_clock = clock; // @[:@154802.4]
  assign regs_237_reset = io_reset; // @[:@154803.4 RegFile.scala 76:16:@154810.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@154809.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@154813.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@154807.4]
  assign regs_238_clock = clock; // @[:@154816.4]
  assign regs_238_reset = io_reset; // @[:@154817.4 RegFile.scala 76:16:@154824.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@154823.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@154827.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@154821.4]
  assign regs_239_clock = clock; // @[:@154830.4]
  assign regs_239_reset = io_reset; // @[:@154831.4 RegFile.scala 76:16:@154838.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@154837.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@154841.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@154835.4]
  assign regs_240_clock = clock; // @[:@154844.4]
  assign regs_240_reset = io_reset; // @[:@154845.4 RegFile.scala 76:16:@154852.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@154851.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@154855.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@154849.4]
  assign regs_241_clock = clock; // @[:@154858.4]
  assign regs_241_reset = io_reset; // @[:@154859.4 RegFile.scala 76:16:@154866.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@154865.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@154869.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@154863.4]
  assign regs_242_clock = clock; // @[:@154872.4]
  assign regs_242_reset = io_reset; // @[:@154873.4 RegFile.scala 76:16:@154880.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@154879.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@154883.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@154877.4]
  assign regs_243_clock = clock; // @[:@154886.4]
  assign regs_243_reset = io_reset; // @[:@154887.4 RegFile.scala 76:16:@154894.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@154893.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@154897.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@154891.4]
  assign regs_244_clock = clock; // @[:@154900.4]
  assign regs_244_reset = io_reset; // @[:@154901.4 RegFile.scala 76:16:@154908.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@154907.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@154911.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@154905.4]
  assign regs_245_clock = clock; // @[:@154914.4]
  assign regs_245_reset = io_reset; // @[:@154915.4 RegFile.scala 76:16:@154922.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@154921.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@154925.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@154919.4]
  assign regs_246_clock = clock; // @[:@154928.4]
  assign regs_246_reset = io_reset; // @[:@154929.4 RegFile.scala 76:16:@154936.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@154935.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@154939.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@154933.4]
  assign regs_247_clock = clock; // @[:@154942.4]
  assign regs_247_reset = io_reset; // @[:@154943.4 RegFile.scala 76:16:@154950.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@154949.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@154953.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@154947.4]
  assign regs_248_clock = clock; // @[:@154956.4]
  assign regs_248_reset = io_reset; // @[:@154957.4 RegFile.scala 76:16:@154964.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@154963.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@154967.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@154961.4]
  assign regs_249_clock = clock; // @[:@154970.4]
  assign regs_249_reset = io_reset; // @[:@154971.4 RegFile.scala 76:16:@154978.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@154977.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@154981.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@154975.4]
  assign regs_250_clock = clock; // @[:@154984.4]
  assign regs_250_reset = io_reset; // @[:@154985.4 RegFile.scala 76:16:@154992.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@154991.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@154995.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@154989.4]
  assign regs_251_clock = clock; // @[:@154998.4]
  assign regs_251_reset = io_reset; // @[:@154999.4 RegFile.scala 76:16:@155006.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@155005.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@155009.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@155003.4]
  assign regs_252_clock = clock; // @[:@155012.4]
  assign regs_252_reset = io_reset; // @[:@155013.4 RegFile.scala 76:16:@155020.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@155019.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@155023.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@155017.4]
  assign regs_253_clock = clock; // @[:@155026.4]
  assign regs_253_reset = io_reset; // @[:@155027.4 RegFile.scala 76:16:@155034.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@155033.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@155037.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@155031.4]
  assign regs_254_clock = clock; // @[:@155040.4]
  assign regs_254_reset = io_reset; // @[:@155041.4 RegFile.scala 76:16:@155048.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@155047.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@155051.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@155045.4]
  assign regs_255_clock = clock; // @[:@155054.4]
  assign regs_255_reset = io_reset; // @[:@155055.4 RegFile.scala 76:16:@155062.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@155061.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@155065.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@155059.4]
  assign regs_256_clock = clock; // @[:@155068.4]
  assign regs_256_reset = io_reset; // @[:@155069.4 RegFile.scala 76:16:@155076.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@155075.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@155079.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@155073.4]
  assign regs_257_clock = clock; // @[:@155082.4]
  assign regs_257_reset = io_reset; // @[:@155083.4 RegFile.scala 76:16:@155090.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@155089.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@155093.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@155087.4]
  assign regs_258_clock = clock; // @[:@155096.4]
  assign regs_258_reset = io_reset; // @[:@155097.4 RegFile.scala 76:16:@155104.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@155103.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@155107.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@155101.4]
  assign regs_259_clock = clock; // @[:@155110.4]
  assign regs_259_reset = io_reset; // @[:@155111.4 RegFile.scala 76:16:@155118.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@155117.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@155121.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@155115.4]
  assign regs_260_clock = clock; // @[:@155124.4]
  assign regs_260_reset = io_reset; // @[:@155125.4 RegFile.scala 76:16:@155132.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@155131.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@155135.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@155129.4]
  assign regs_261_clock = clock; // @[:@155138.4]
  assign regs_261_reset = io_reset; // @[:@155139.4 RegFile.scala 76:16:@155146.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@155145.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@155149.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@155143.4]
  assign regs_262_clock = clock; // @[:@155152.4]
  assign regs_262_reset = io_reset; // @[:@155153.4 RegFile.scala 76:16:@155160.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@155159.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@155163.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@155157.4]
  assign regs_263_clock = clock; // @[:@155166.4]
  assign regs_263_reset = io_reset; // @[:@155167.4 RegFile.scala 76:16:@155174.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@155173.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@155177.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@155171.4]
  assign regs_264_clock = clock; // @[:@155180.4]
  assign regs_264_reset = io_reset; // @[:@155181.4 RegFile.scala 76:16:@155188.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@155187.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@155191.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@155185.4]
  assign regs_265_clock = clock; // @[:@155194.4]
  assign regs_265_reset = io_reset; // @[:@155195.4 RegFile.scala 76:16:@155202.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@155201.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@155205.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@155199.4]
  assign regs_266_clock = clock; // @[:@155208.4]
  assign regs_266_reset = io_reset; // @[:@155209.4 RegFile.scala 76:16:@155216.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@155215.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@155219.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@155213.4]
  assign regs_267_clock = clock; // @[:@155222.4]
  assign regs_267_reset = io_reset; // @[:@155223.4 RegFile.scala 76:16:@155230.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@155229.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@155233.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@155227.4]
  assign regs_268_clock = clock; // @[:@155236.4]
  assign regs_268_reset = io_reset; // @[:@155237.4 RegFile.scala 76:16:@155244.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@155243.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@155247.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@155241.4]
  assign regs_269_clock = clock; // @[:@155250.4]
  assign regs_269_reset = io_reset; // @[:@155251.4 RegFile.scala 76:16:@155258.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@155257.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@155261.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@155255.4]
  assign regs_270_clock = clock; // @[:@155264.4]
  assign regs_270_reset = io_reset; // @[:@155265.4 RegFile.scala 76:16:@155272.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@155271.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@155275.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@155269.4]
  assign regs_271_clock = clock; // @[:@155278.4]
  assign regs_271_reset = io_reset; // @[:@155279.4 RegFile.scala 76:16:@155286.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@155285.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@155289.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@155283.4]
  assign regs_272_clock = clock; // @[:@155292.4]
  assign regs_272_reset = io_reset; // @[:@155293.4 RegFile.scala 76:16:@155300.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@155299.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@155303.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@155297.4]
  assign regs_273_clock = clock; // @[:@155306.4]
  assign regs_273_reset = io_reset; // @[:@155307.4 RegFile.scala 76:16:@155314.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@155313.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@155317.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@155311.4]
  assign regs_274_clock = clock; // @[:@155320.4]
  assign regs_274_reset = io_reset; // @[:@155321.4 RegFile.scala 76:16:@155328.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@155327.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@155331.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@155325.4]
  assign regs_275_clock = clock; // @[:@155334.4]
  assign regs_275_reset = io_reset; // @[:@155335.4 RegFile.scala 76:16:@155342.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@155341.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@155345.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@155339.4]
  assign regs_276_clock = clock; // @[:@155348.4]
  assign regs_276_reset = io_reset; // @[:@155349.4 RegFile.scala 76:16:@155356.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@155355.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@155359.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@155353.4]
  assign regs_277_clock = clock; // @[:@155362.4]
  assign regs_277_reset = io_reset; // @[:@155363.4 RegFile.scala 76:16:@155370.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@155369.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@155373.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@155367.4]
  assign regs_278_clock = clock; // @[:@155376.4]
  assign regs_278_reset = io_reset; // @[:@155377.4 RegFile.scala 76:16:@155384.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@155383.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@155387.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@155381.4]
  assign regs_279_clock = clock; // @[:@155390.4]
  assign regs_279_reset = io_reset; // @[:@155391.4 RegFile.scala 76:16:@155398.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@155397.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@155401.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@155395.4]
  assign regs_280_clock = clock; // @[:@155404.4]
  assign regs_280_reset = io_reset; // @[:@155405.4 RegFile.scala 76:16:@155412.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@155411.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@155415.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@155409.4]
  assign regs_281_clock = clock; // @[:@155418.4]
  assign regs_281_reset = io_reset; // @[:@155419.4 RegFile.scala 76:16:@155426.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@155425.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@155429.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@155423.4]
  assign regs_282_clock = clock; // @[:@155432.4]
  assign regs_282_reset = io_reset; // @[:@155433.4 RegFile.scala 76:16:@155440.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@155439.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@155443.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@155437.4]
  assign regs_283_clock = clock; // @[:@155446.4]
  assign regs_283_reset = io_reset; // @[:@155447.4 RegFile.scala 76:16:@155454.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@155453.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@155457.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@155451.4]
  assign regs_284_clock = clock; // @[:@155460.4]
  assign regs_284_reset = io_reset; // @[:@155461.4 RegFile.scala 76:16:@155468.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@155467.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@155471.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@155465.4]
  assign regs_285_clock = clock; // @[:@155474.4]
  assign regs_285_reset = io_reset; // @[:@155475.4 RegFile.scala 76:16:@155482.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@155481.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@155485.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@155479.4]
  assign regs_286_clock = clock; // @[:@155488.4]
  assign regs_286_reset = io_reset; // @[:@155489.4 RegFile.scala 76:16:@155496.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@155495.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@155499.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@155493.4]
  assign regs_287_clock = clock; // @[:@155502.4]
  assign regs_287_reset = io_reset; // @[:@155503.4 RegFile.scala 76:16:@155510.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@155509.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@155513.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@155507.4]
  assign regs_288_clock = clock; // @[:@155516.4]
  assign regs_288_reset = io_reset; // @[:@155517.4 RegFile.scala 76:16:@155524.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@155523.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@155527.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@155521.4]
  assign regs_289_clock = clock; // @[:@155530.4]
  assign regs_289_reset = io_reset; // @[:@155531.4 RegFile.scala 76:16:@155538.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@155537.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@155541.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@155535.4]
  assign regs_290_clock = clock; // @[:@155544.4]
  assign regs_290_reset = io_reset; // @[:@155545.4 RegFile.scala 76:16:@155552.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@155551.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@155555.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@155549.4]
  assign regs_291_clock = clock; // @[:@155558.4]
  assign regs_291_reset = io_reset; // @[:@155559.4 RegFile.scala 76:16:@155566.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@155565.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@155569.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@155563.4]
  assign regs_292_clock = clock; // @[:@155572.4]
  assign regs_292_reset = io_reset; // @[:@155573.4 RegFile.scala 76:16:@155580.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@155579.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@155583.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@155577.4]
  assign regs_293_clock = clock; // @[:@155586.4]
  assign regs_293_reset = io_reset; // @[:@155587.4 RegFile.scala 76:16:@155594.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@155593.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@155597.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@155591.4]
  assign regs_294_clock = clock; // @[:@155600.4]
  assign regs_294_reset = io_reset; // @[:@155601.4 RegFile.scala 76:16:@155608.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@155607.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@155611.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@155605.4]
  assign regs_295_clock = clock; // @[:@155614.4]
  assign regs_295_reset = io_reset; // @[:@155615.4 RegFile.scala 76:16:@155622.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@155621.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@155625.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@155619.4]
  assign regs_296_clock = clock; // @[:@155628.4]
  assign regs_296_reset = io_reset; // @[:@155629.4 RegFile.scala 76:16:@155636.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@155635.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@155639.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@155633.4]
  assign regs_297_clock = clock; // @[:@155642.4]
  assign regs_297_reset = io_reset; // @[:@155643.4 RegFile.scala 76:16:@155650.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@155649.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@155653.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@155647.4]
  assign regs_298_clock = clock; // @[:@155656.4]
  assign regs_298_reset = io_reset; // @[:@155657.4 RegFile.scala 76:16:@155664.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@155663.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@155667.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@155661.4]
  assign regs_299_clock = clock; // @[:@155670.4]
  assign regs_299_reset = io_reset; // @[:@155671.4 RegFile.scala 76:16:@155678.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@155677.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@155681.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@155675.4]
  assign regs_300_clock = clock; // @[:@155684.4]
  assign regs_300_reset = io_reset; // @[:@155685.4 RegFile.scala 76:16:@155692.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@155691.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@155695.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@155689.4]
  assign regs_301_clock = clock; // @[:@155698.4]
  assign regs_301_reset = io_reset; // @[:@155699.4 RegFile.scala 76:16:@155706.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@155705.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@155709.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@155703.4]
  assign regs_302_clock = clock; // @[:@155712.4]
  assign regs_302_reset = io_reset; // @[:@155713.4 RegFile.scala 76:16:@155720.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@155719.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@155723.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@155717.4]
  assign regs_303_clock = clock; // @[:@155726.4]
  assign regs_303_reset = io_reset; // @[:@155727.4 RegFile.scala 76:16:@155734.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@155733.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@155737.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@155731.4]
  assign regs_304_clock = clock; // @[:@155740.4]
  assign regs_304_reset = io_reset; // @[:@155741.4 RegFile.scala 76:16:@155748.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@155747.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@155751.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@155745.4]
  assign regs_305_clock = clock; // @[:@155754.4]
  assign regs_305_reset = io_reset; // @[:@155755.4 RegFile.scala 76:16:@155762.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@155761.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@155765.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@155759.4]
  assign regs_306_clock = clock; // @[:@155768.4]
  assign regs_306_reset = io_reset; // @[:@155769.4 RegFile.scala 76:16:@155776.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@155775.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@155779.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@155773.4]
  assign regs_307_clock = clock; // @[:@155782.4]
  assign regs_307_reset = io_reset; // @[:@155783.4 RegFile.scala 76:16:@155790.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@155789.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@155793.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@155787.4]
  assign regs_308_clock = clock; // @[:@155796.4]
  assign regs_308_reset = io_reset; // @[:@155797.4 RegFile.scala 76:16:@155804.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@155803.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@155807.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@155801.4]
  assign regs_309_clock = clock; // @[:@155810.4]
  assign regs_309_reset = io_reset; // @[:@155811.4 RegFile.scala 76:16:@155818.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@155817.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@155821.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@155815.4]
  assign regs_310_clock = clock; // @[:@155824.4]
  assign regs_310_reset = io_reset; // @[:@155825.4 RegFile.scala 76:16:@155832.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@155831.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@155835.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@155829.4]
  assign regs_311_clock = clock; // @[:@155838.4]
  assign regs_311_reset = io_reset; // @[:@155839.4 RegFile.scala 76:16:@155846.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@155845.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@155849.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@155843.4]
  assign regs_312_clock = clock; // @[:@155852.4]
  assign regs_312_reset = io_reset; // @[:@155853.4 RegFile.scala 76:16:@155860.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@155859.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@155863.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@155857.4]
  assign regs_313_clock = clock; // @[:@155866.4]
  assign regs_313_reset = io_reset; // @[:@155867.4 RegFile.scala 76:16:@155874.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@155873.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@155877.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@155871.4]
  assign regs_314_clock = clock; // @[:@155880.4]
  assign regs_314_reset = io_reset; // @[:@155881.4 RegFile.scala 76:16:@155888.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@155887.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@155891.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@155885.4]
  assign regs_315_clock = clock; // @[:@155894.4]
  assign regs_315_reset = io_reset; // @[:@155895.4 RegFile.scala 76:16:@155902.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@155901.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@155905.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@155899.4]
  assign regs_316_clock = clock; // @[:@155908.4]
  assign regs_316_reset = io_reset; // @[:@155909.4 RegFile.scala 76:16:@155916.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@155915.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@155919.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@155913.4]
  assign regs_317_clock = clock; // @[:@155922.4]
  assign regs_317_reset = io_reset; // @[:@155923.4 RegFile.scala 76:16:@155930.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@155929.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@155933.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@155927.4]
  assign regs_318_clock = clock; // @[:@155936.4]
  assign regs_318_reset = io_reset; // @[:@155937.4 RegFile.scala 76:16:@155944.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@155943.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@155947.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@155941.4]
  assign regs_319_clock = clock; // @[:@155950.4]
  assign regs_319_reset = io_reset; // @[:@155951.4 RegFile.scala 76:16:@155958.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@155957.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@155961.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@155955.4]
  assign regs_320_clock = clock; // @[:@155964.4]
  assign regs_320_reset = io_reset; // @[:@155965.4 RegFile.scala 76:16:@155972.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@155971.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@155975.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@155969.4]
  assign regs_321_clock = clock; // @[:@155978.4]
  assign regs_321_reset = io_reset; // @[:@155979.4 RegFile.scala 76:16:@155986.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@155985.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@155989.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@155983.4]
  assign regs_322_clock = clock; // @[:@155992.4]
  assign regs_322_reset = io_reset; // @[:@155993.4 RegFile.scala 76:16:@156000.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@155999.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@156003.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@155997.4]
  assign regs_323_clock = clock; // @[:@156006.4]
  assign regs_323_reset = io_reset; // @[:@156007.4 RegFile.scala 76:16:@156014.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@156013.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@156017.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@156011.4]
  assign regs_324_clock = clock; // @[:@156020.4]
  assign regs_324_reset = io_reset; // @[:@156021.4 RegFile.scala 76:16:@156028.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@156027.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@156031.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@156025.4]
  assign regs_325_clock = clock; // @[:@156034.4]
  assign regs_325_reset = io_reset; // @[:@156035.4 RegFile.scala 76:16:@156042.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@156041.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@156045.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@156039.4]
  assign regs_326_clock = clock; // @[:@156048.4]
  assign regs_326_reset = io_reset; // @[:@156049.4 RegFile.scala 76:16:@156056.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@156055.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@156059.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@156053.4]
  assign regs_327_clock = clock; // @[:@156062.4]
  assign regs_327_reset = io_reset; // @[:@156063.4 RegFile.scala 76:16:@156070.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@156069.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@156073.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@156067.4]
  assign regs_328_clock = clock; // @[:@156076.4]
  assign regs_328_reset = io_reset; // @[:@156077.4 RegFile.scala 76:16:@156084.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@156083.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@156087.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@156081.4]
  assign regs_329_clock = clock; // @[:@156090.4]
  assign regs_329_reset = io_reset; // @[:@156091.4 RegFile.scala 76:16:@156098.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@156097.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@156101.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@156095.4]
  assign regs_330_clock = clock; // @[:@156104.4]
  assign regs_330_reset = io_reset; // @[:@156105.4 RegFile.scala 76:16:@156112.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@156111.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@156115.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@156109.4]
  assign regs_331_clock = clock; // @[:@156118.4]
  assign regs_331_reset = io_reset; // @[:@156119.4 RegFile.scala 76:16:@156126.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@156125.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@156129.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@156123.4]
  assign regs_332_clock = clock; // @[:@156132.4]
  assign regs_332_reset = io_reset; // @[:@156133.4 RegFile.scala 76:16:@156140.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@156139.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@156143.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@156137.4]
  assign regs_333_clock = clock; // @[:@156146.4]
  assign regs_333_reset = io_reset; // @[:@156147.4 RegFile.scala 76:16:@156154.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@156153.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@156157.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@156151.4]
  assign regs_334_clock = clock; // @[:@156160.4]
  assign regs_334_reset = io_reset; // @[:@156161.4 RegFile.scala 76:16:@156168.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@156167.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@156171.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@156165.4]
  assign regs_335_clock = clock; // @[:@156174.4]
  assign regs_335_reset = io_reset; // @[:@156175.4 RegFile.scala 76:16:@156182.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@156181.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@156185.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@156179.4]
  assign regs_336_clock = clock; // @[:@156188.4]
  assign regs_336_reset = io_reset; // @[:@156189.4 RegFile.scala 76:16:@156196.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@156195.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@156199.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@156193.4]
  assign regs_337_clock = clock; // @[:@156202.4]
  assign regs_337_reset = io_reset; // @[:@156203.4 RegFile.scala 76:16:@156210.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@156209.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@156213.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@156207.4]
  assign regs_338_clock = clock; // @[:@156216.4]
  assign regs_338_reset = io_reset; // @[:@156217.4 RegFile.scala 76:16:@156224.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@156223.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@156227.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@156221.4]
  assign regs_339_clock = clock; // @[:@156230.4]
  assign regs_339_reset = io_reset; // @[:@156231.4 RegFile.scala 76:16:@156238.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@156237.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@156241.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@156235.4]
  assign regs_340_clock = clock; // @[:@156244.4]
  assign regs_340_reset = io_reset; // @[:@156245.4 RegFile.scala 76:16:@156252.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@156251.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@156255.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@156249.4]
  assign regs_341_clock = clock; // @[:@156258.4]
  assign regs_341_reset = io_reset; // @[:@156259.4 RegFile.scala 76:16:@156266.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@156265.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@156269.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@156263.4]
  assign regs_342_clock = clock; // @[:@156272.4]
  assign regs_342_reset = io_reset; // @[:@156273.4 RegFile.scala 76:16:@156280.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@156279.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@156283.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@156277.4]
  assign regs_343_clock = clock; // @[:@156286.4]
  assign regs_343_reset = io_reset; // @[:@156287.4 RegFile.scala 76:16:@156294.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@156293.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@156297.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@156291.4]
  assign regs_344_clock = clock; // @[:@156300.4]
  assign regs_344_reset = io_reset; // @[:@156301.4 RegFile.scala 76:16:@156308.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@156307.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@156311.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@156305.4]
  assign regs_345_clock = clock; // @[:@156314.4]
  assign regs_345_reset = io_reset; // @[:@156315.4 RegFile.scala 76:16:@156322.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@156321.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@156325.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@156319.4]
  assign regs_346_clock = clock; // @[:@156328.4]
  assign regs_346_reset = io_reset; // @[:@156329.4 RegFile.scala 76:16:@156336.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@156335.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@156339.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@156333.4]
  assign regs_347_clock = clock; // @[:@156342.4]
  assign regs_347_reset = io_reset; // @[:@156343.4 RegFile.scala 76:16:@156350.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@156349.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@156353.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@156347.4]
  assign regs_348_clock = clock; // @[:@156356.4]
  assign regs_348_reset = io_reset; // @[:@156357.4 RegFile.scala 76:16:@156364.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@156363.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@156367.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@156361.4]
  assign regs_349_clock = clock; // @[:@156370.4]
  assign regs_349_reset = io_reset; // @[:@156371.4 RegFile.scala 76:16:@156378.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@156377.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@156381.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@156375.4]
  assign regs_350_clock = clock; // @[:@156384.4]
  assign regs_350_reset = io_reset; // @[:@156385.4 RegFile.scala 76:16:@156392.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@156391.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@156395.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@156389.4]
  assign regs_351_clock = clock; // @[:@156398.4]
  assign regs_351_reset = io_reset; // @[:@156399.4 RegFile.scala 76:16:@156406.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@156405.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@156409.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@156403.4]
  assign regs_352_clock = clock; // @[:@156412.4]
  assign regs_352_reset = io_reset; // @[:@156413.4 RegFile.scala 76:16:@156420.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@156419.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@156423.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@156417.4]
  assign regs_353_clock = clock; // @[:@156426.4]
  assign regs_353_reset = io_reset; // @[:@156427.4 RegFile.scala 76:16:@156434.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@156433.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@156437.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@156431.4]
  assign regs_354_clock = clock; // @[:@156440.4]
  assign regs_354_reset = io_reset; // @[:@156441.4 RegFile.scala 76:16:@156448.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@156447.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@156451.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@156445.4]
  assign regs_355_clock = clock; // @[:@156454.4]
  assign regs_355_reset = io_reset; // @[:@156455.4 RegFile.scala 76:16:@156462.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@156461.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@156465.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@156459.4]
  assign regs_356_clock = clock; // @[:@156468.4]
  assign regs_356_reset = io_reset; // @[:@156469.4 RegFile.scala 76:16:@156476.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@156475.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@156479.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@156473.4]
  assign regs_357_clock = clock; // @[:@156482.4]
  assign regs_357_reset = io_reset; // @[:@156483.4 RegFile.scala 76:16:@156490.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@156489.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@156493.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@156487.4]
  assign regs_358_clock = clock; // @[:@156496.4]
  assign regs_358_reset = io_reset; // @[:@156497.4 RegFile.scala 76:16:@156504.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@156503.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@156507.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@156501.4]
  assign regs_359_clock = clock; // @[:@156510.4]
  assign regs_359_reset = io_reset; // @[:@156511.4 RegFile.scala 76:16:@156518.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@156517.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@156521.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@156515.4]
  assign regs_360_clock = clock; // @[:@156524.4]
  assign regs_360_reset = io_reset; // @[:@156525.4 RegFile.scala 76:16:@156532.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@156531.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@156535.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@156529.4]
  assign regs_361_clock = clock; // @[:@156538.4]
  assign regs_361_reset = io_reset; // @[:@156539.4 RegFile.scala 76:16:@156546.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@156545.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@156549.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@156543.4]
  assign regs_362_clock = clock; // @[:@156552.4]
  assign regs_362_reset = io_reset; // @[:@156553.4 RegFile.scala 76:16:@156560.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@156559.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@156563.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@156557.4]
  assign regs_363_clock = clock; // @[:@156566.4]
  assign regs_363_reset = io_reset; // @[:@156567.4 RegFile.scala 76:16:@156574.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@156573.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@156577.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@156571.4]
  assign regs_364_clock = clock; // @[:@156580.4]
  assign regs_364_reset = io_reset; // @[:@156581.4 RegFile.scala 76:16:@156588.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@156587.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@156591.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@156585.4]
  assign regs_365_clock = clock; // @[:@156594.4]
  assign regs_365_reset = io_reset; // @[:@156595.4 RegFile.scala 76:16:@156602.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@156601.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@156605.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@156599.4]
  assign regs_366_clock = clock; // @[:@156608.4]
  assign regs_366_reset = io_reset; // @[:@156609.4 RegFile.scala 76:16:@156616.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@156615.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@156619.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@156613.4]
  assign regs_367_clock = clock; // @[:@156622.4]
  assign regs_367_reset = io_reset; // @[:@156623.4 RegFile.scala 76:16:@156630.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@156629.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@156633.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@156627.4]
  assign regs_368_clock = clock; // @[:@156636.4]
  assign regs_368_reset = io_reset; // @[:@156637.4 RegFile.scala 76:16:@156644.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@156643.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@156647.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@156641.4]
  assign regs_369_clock = clock; // @[:@156650.4]
  assign regs_369_reset = io_reset; // @[:@156651.4 RegFile.scala 76:16:@156658.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@156657.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@156661.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@156655.4]
  assign regs_370_clock = clock; // @[:@156664.4]
  assign regs_370_reset = io_reset; // @[:@156665.4 RegFile.scala 76:16:@156672.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@156671.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@156675.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@156669.4]
  assign regs_371_clock = clock; // @[:@156678.4]
  assign regs_371_reset = io_reset; // @[:@156679.4 RegFile.scala 76:16:@156686.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@156685.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@156689.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@156683.4]
  assign regs_372_clock = clock; // @[:@156692.4]
  assign regs_372_reset = io_reset; // @[:@156693.4 RegFile.scala 76:16:@156700.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@156699.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@156703.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@156697.4]
  assign regs_373_clock = clock; // @[:@156706.4]
  assign regs_373_reset = io_reset; // @[:@156707.4 RegFile.scala 76:16:@156714.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@156713.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@156717.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@156711.4]
  assign regs_374_clock = clock; // @[:@156720.4]
  assign regs_374_reset = io_reset; // @[:@156721.4 RegFile.scala 76:16:@156728.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@156727.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@156731.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@156725.4]
  assign regs_375_clock = clock; // @[:@156734.4]
  assign regs_375_reset = io_reset; // @[:@156735.4 RegFile.scala 76:16:@156742.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@156741.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@156745.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@156739.4]
  assign regs_376_clock = clock; // @[:@156748.4]
  assign regs_376_reset = io_reset; // @[:@156749.4 RegFile.scala 76:16:@156756.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@156755.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@156759.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@156753.4]
  assign regs_377_clock = clock; // @[:@156762.4]
  assign regs_377_reset = io_reset; // @[:@156763.4 RegFile.scala 76:16:@156770.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@156769.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@156773.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@156767.4]
  assign regs_378_clock = clock; // @[:@156776.4]
  assign regs_378_reset = io_reset; // @[:@156777.4 RegFile.scala 76:16:@156784.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@156783.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@156787.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@156781.4]
  assign regs_379_clock = clock; // @[:@156790.4]
  assign regs_379_reset = io_reset; // @[:@156791.4 RegFile.scala 76:16:@156798.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@156797.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@156801.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@156795.4]
  assign regs_380_clock = clock; // @[:@156804.4]
  assign regs_380_reset = io_reset; // @[:@156805.4 RegFile.scala 76:16:@156812.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@156811.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@156815.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@156809.4]
  assign regs_381_clock = clock; // @[:@156818.4]
  assign regs_381_reset = io_reset; // @[:@156819.4 RegFile.scala 76:16:@156826.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@156825.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@156829.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@156823.4]
  assign regs_382_clock = clock; // @[:@156832.4]
  assign regs_382_reset = io_reset; // @[:@156833.4 RegFile.scala 76:16:@156840.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@156839.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@156843.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@156837.4]
  assign regs_383_clock = clock; // @[:@156846.4]
  assign regs_383_reset = io_reset; // @[:@156847.4 RegFile.scala 76:16:@156854.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@156853.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@156857.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@156851.4]
  assign regs_384_clock = clock; // @[:@156860.4]
  assign regs_384_reset = io_reset; // @[:@156861.4 RegFile.scala 76:16:@156868.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@156867.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@156871.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@156865.4]
  assign regs_385_clock = clock; // @[:@156874.4]
  assign regs_385_reset = io_reset; // @[:@156875.4 RegFile.scala 76:16:@156882.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@156881.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@156885.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@156879.4]
  assign regs_386_clock = clock; // @[:@156888.4]
  assign regs_386_reset = io_reset; // @[:@156889.4 RegFile.scala 76:16:@156896.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@156895.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@156899.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@156893.4]
  assign regs_387_clock = clock; // @[:@156902.4]
  assign regs_387_reset = io_reset; // @[:@156903.4 RegFile.scala 76:16:@156910.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@156909.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@156913.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@156907.4]
  assign regs_388_clock = clock; // @[:@156916.4]
  assign regs_388_reset = io_reset; // @[:@156917.4 RegFile.scala 76:16:@156924.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@156923.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@156927.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@156921.4]
  assign regs_389_clock = clock; // @[:@156930.4]
  assign regs_389_reset = io_reset; // @[:@156931.4 RegFile.scala 76:16:@156938.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@156937.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@156941.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@156935.4]
  assign regs_390_clock = clock; // @[:@156944.4]
  assign regs_390_reset = io_reset; // @[:@156945.4 RegFile.scala 76:16:@156952.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@156951.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@156955.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@156949.4]
  assign regs_391_clock = clock; // @[:@156958.4]
  assign regs_391_reset = io_reset; // @[:@156959.4 RegFile.scala 76:16:@156966.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@156965.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@156969.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@156963.4]
  assign regs_392_clock = clock; // @[:@156972.4]
  assign regs_392_reset = io_reset; // @[:@156973.4 RegFile.scala 76:16:@156980.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@156979.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@156983.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@156977.4]
  assign regs_393_clock = clock; // @[:@156986.4]
  assign regs_393_reset = io_reset; // @[:@156987.4 RegFile.scala 76:16:@156994.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@156993.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@156997.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@156991.4]
  assign regs_394_clock = clock; // @[:@157000.4]
  assign regs_394_reset = io_reset; // @[:@157001.4 RegFile.scala 76:16:@157008.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@157007.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@157011.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@157005.4]
  assign regs_395_clock = clock; // @[:@157014.4]
  assign regs_395_reset = io_reset; // @[:@157015.4 RegFile.scala 76:16:@157022.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@157021.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@157025.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@157019.4]
  assign regs_396_clock = clock; // @[:@157028.4]
  assign regs_396_reset = io_reset; // @[:@157029.4 RegFile.scala 76:16:@157036.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@157035.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@157039.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@157033.4]
  assign regs_397_clock = clock; // @[:@157042.4]
  assign regs_397_reset = io_reset; // @[:@157043.4 RegFile.scala 76:16:@157050.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@157049.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@157053.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@157047.4]
  assign regs_398_clock = clock; // @[:@157056.4]
  assign regs_398_reset = io_reset; // @[:@157057.4 RegFile.scala 76:16:@157064.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@157063.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@157067.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@157061.4]
  assign regs_399_clock = clock; // @[:@157070.4]
  assign regs_399_reset = io_reset; // @[:@157071.4 RegFile.scala 76:16:@157078.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@157077.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@157081.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@157075.4]
  assign regs_400_clock = clock; // @[:@157084.4]
  assign regs_400_reset = io_reset; // @[:@157085.4 RegFile.scala 76:16:@157092.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@157091.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@157095.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@157089.4]
  assign regs_401_clock = clock; // @[:@157098.4]
  assign regs_401_reset = io_reset; // @[:@157099.4 RegFile.scala 76:16:@157106.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@157105.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@157109.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@157103.4]
  assign regs_402_clock = clock; // @[:@157112.4]
  assign regs_402_reset = io_reset; // @[:@157113.4 RegFile.scala 76:16:@157120.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@157119.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@157123.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@157117.4]
  assign regs_403_clock = clock; // @[:@157126.4]
  assign regs_403_reset = io_reset; // @[:@157127.4 RegFile.scala 76:16:@157134.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@157133.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@157137.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@157131.4]
  assign regs_404_clock = clock; // @[:@157140.4]
  assign regs_404_reset = io_reset; // @[:@157141.4 RegFile.scala 76:16:@157148.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@157147.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@157151.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@157145.4]
  assign regs_405_clock = clock; // @[:@157154.4]
  assign regs_405_reset = io_reset; // @[:@157155.4 RegFile.scala 76:16:@157162.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@157161.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@157165.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@157159.4]
  assign regs_406_clock = clock; // @[:@157168.4]
  assign regs_406_reset = io_reset; // @[:@157169.4 RegFile.scala 76:16:@157176.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@157175.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@157179.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@157173.4]
  assign regs_407_clock = clock; // @[:@157182.4]
  assign regs_407_reset = io_reset; // @[:@157183.4 RegFile.scala 76:16:@157190.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@157189.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@157193.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@157187.4]
  assign regs_408_clock = clock; // @[:@157196.4]
  assign regs_408_reset = io_reset; // @[:@157197.4 RegFile.scala 76:16:@157204.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@157203.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@157207.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@157201.4]
  assign regs_409_clock = clock; // @[:@157210.4]
  assign regs_409_reset = io_reset; // @[:@157211.4 RegFile.scala 76:16:@157218.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@157217.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@157221.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@157215.4]
  assign regs_410_clock = clock; // @[:@157224.4]
  assign regs_410_reset = io_reset; // @[:@157225.4 RegFile.scala 76:16:@157232.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@157231.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@157235.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@157229.4]
  assign regs_411_clock = clock; // @[:@157238.4]
  assign regs_411_reset = io_reset; // @[:@157239.4 RegFile.scala 76:16:@157246.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@157245.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@157249.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@157243.4]
  assign regs_412_clock = clock; // @[:@157252.4]
  assign regs_412_reset = io_reset; // @[:@157253.4 RegFile.scala 76:16:@157260.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@157259.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@157263.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@157257.4]
  assign regs_413_clock = clock; // @[:@157266.4]
  assign regs_413_reset = io_reset; // @[:@157267.4 RegFile.scala 76:16:@157274.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@157273.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@157277.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@157271.4]
  assign regs_414_clock = clock; // @[:@157280.4]
  assign regs_414_reset = io_reset; // @[:@157281.4 RegFile.scala 76:16:@157288.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@157287.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@157291.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@157285.4]
  assign regs_415_clock = clock; // @[:@157294.4]
  assign regs_415_reset = io_reset; // @[:@157295.4 RegFile.scala 76:16:@157302.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@157301.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@157305.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@157299.4]
  assign regs_416_clock = clock; // @[:@157308.4]
  assign regs_416_reset = io_reset; // @[:@157309.4 RegFile.scala 76:16:@157316.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@157315.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@157319.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@157313.4]
  assign regs_417_clock = clock; // @[:@157322.4]
  assign regs_417_reset = io_reset; // @[:@157323.4 RegFile.scala 76:16:@157330.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@157329.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@157333.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@157327.4]
  assign regs_418_clock = clock; // @[:@157336.4]
  assign regs_418_reset = io_reset; // @[:@157337.4 RegFile.scala 76:16:@157344.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@157343.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@157347.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@157341.4]
  assign regs_419_clock = clock; // @[:@157350.4]
  assign regs_419_reset = io_reset; // @[:@157351.4 RegFile.scala 76:16:@157358.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@157357.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@157361.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@157355.4]
  assign regs_420_clock = clock; // @[:@157364.4]
  assign regs_420_reset = io_reset; // @[:@157365.4 RegFile.scala 76:16:@157372.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@157371.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@157375.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@157369.4]
  assign regs_421_clock = clock; // @[:@157378.4]
  assign regs_421_reset = io_reset; // @[:@157379.4 RegFile.scala 76:16:@157386.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@157385.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@157389.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@157383.4]
  assign regs_422_clock = clock; // @[:@157392.4]
  assign regs_422_reset = io_reset; // @[:@157393.4 RegFile.scala 76:16:@157400.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@157399.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@157403.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@157397.4]
  assign regs_423_clock = clock; // @[:@157406.4]
  assign regs_423_reset = io_reset; // @[:@157407.4 RegFile.scala 76:16:@157414.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@157413.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@157417.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@157411.4]
  assign regs_424_clock = clock; // @[:@157420.4]
  assign regs_424_reset = io_reset; // @[:@157421.4 RegFile.scala 76:16:@157428.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@157427.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@157431.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@157425.4]
  assign regs_425_clock = clock; // @[:@157434.4]
  assign regs_425_reset = io_reset; // @[:@157435.4 RegFile.scala 76:16:@157442.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@157441.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@157445.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@157439.4]
  assign regs_426_clock = clock; // @[:@157448.4]
  assign regs_426_reset = io_reset; // @[:@157449.4 RegFile.scala 76:16:@157456.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@157455.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@157459.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@157453.4]
  assign regs_427_clock = clock; // @[:@157462.4]
  assign regs_427_reset = io_reset; // @[:@157463.4 RegFile.scala 76:16:@157470.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@157469.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@157473.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@157467.4]
  assign regs_428_clock = clock; // @[:@157476.4]
  assign regs_428_reset = io_reset; // @[:@157477.4 RegFile.scala 76:16:@157484.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@157483.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@157487.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@157481.4]
  assign regs_429_clock = clock; // @[:@157490.4]
  assign regs_429_reset = io_reset; // @[:@157491.4 RegFile.scala 76:16:@157498.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@157497.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@157501.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@157495.4]
  assign regs_430_clock = clock; // @[:@157504.4]
  assign regs_430_reset = io_reset; // @[:@157505.4 RegFile.scala 76:16:@157512.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@157511.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@157515.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@157509.4]
  assign regs_431_clock = clock; // @[:@157518.4]
  assign regs_431_reset = io_reset; // @[:@157519.4 RegFile.scala 76:16:@157526.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@157525.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@157529.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@157523.4]
  assign regs_432_clock = clock; // @[:@157532.4]
  assign regs_432_reset = io_reset; // @[:@157533.4 RegFile.scala 76:16:@157540.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@157539.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@157543.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@157537.4]
  assign regs_433_clock = clock; // @[:@157546.4]
  assign regs_433_reset = io_reset; // @[:@157547.4 RegFile.scala 76:16:@157554.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@157553.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@157557.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@157551.4]
  assign regs_434_clock = clock; // @[:@157560.4]
  assign regs_434_reset = io_reset; // @[:@157561.4 RegFile.scala 76:16:@157568.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@157567.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@157571.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@157565.4]
  assign regs_435_clock = clock; // @[:@157574.4]
  assign regs_435_reset = io_reset; // @[:@157575.4 RegFile.scala 76:16:@157582.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@157581.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@157585.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@157579.4]
  assign regs_436_clock = clock; // @[:@157588.4]
  assign regs_436_reset = io_reset; // @[:@157589.4 RegFile.scala 76:16:@157596.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@157595.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@157599.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@157593.4]
  assign regs_437_clock = clock; // @[:@157602.4]
  assign regs_437_reset = io_reset; // @[:@157603.4 RegFile.scala 76:16:@157610.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@157609.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@157613.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@157607.4]
  assign regs_438_clock = clock; // @[:@157616.4]
  assign regs_438_reset = io_reset; // @[:@157617.4 RegFile.scala 76:16:@157624.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@157623.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@157627.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@157621.4]
  assign regs_439_clock = clock; // @[:@157630.4]
  assign regs_439_reset = io_reset; // @[:@157631.4 RegFile.scala 76:16:@157638.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@157637.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@157641.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@157635.4]
  assign regs_440_clock = clock; // @[:@157644.4]
  assign regs_440_reset = io_reset; // @[:@157645.4 RegFile.scala 76:16:@157652.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@157651.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@157655.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@157649.4]
  assign regs_441_clock = clock; // @[:@157658.4]
  assign regs_441_reset = io_reset; // @[:@157659.4 RegFile.scala 76:16:@157666.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@157665.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@157669.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@157663.4]
  assign regs_442_clock = clock; // @[:@157672.4]
  assign regs_442_reset = io_reset; // @[:@157673.4 RegFile.scala 76:16:@157680.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@157679.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@157683.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@157677.4]
  assign regs_443_clock = clock; // @[:@157686.4]
  assign regs_443_reset = io_reset; // @[:@157687.4 RegFile.scala 76:16:@157694.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@157693.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@157697.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@157691.4]
  assign regs_444_clock = clock; // @[:@157700.4]
  assign regs_444_reset = io_reset; // @[:@157701.4 RegFile.scala 76:16:@157708.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@157707.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@157711.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@157705.4]
  assign regs_445_clock = clock; // @[:@157714.4]
  assign regs_445_reset = io_reset; // @[:@157715.4 RegFile.scala 76:16:@157722.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@157721.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@157725.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@157719.4]
  assign regs_446_clock = clock; // @[:@157728.4]
  assign regs_446_reset = io_reset; // @[:@157729.4 RegFile.scala 76:16:@157736.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@157735.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@157739.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@157733.4]
  assign regs_447_clock = clock; // @[:@157742.4]
  assign regs_447_reset = io_reset; // @[:@157743.4 RegFile.scala 76:16:@157750.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@157749.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@157753.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@157747.4]
  assign regs_448_clock = clock; // @[:@157756.4]
  assign regs_448_reset = io_reset; // @[:@157757.4 RegFile.scala 76:16:@157764.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@157763.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@157767.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@157761.4]
  assign regs_449_clock = clock; // @[:@157770.4]
  assign regs_449_reset = io_reset; // @[:@157771.4 RegFile.scala 76:16:@157778.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@157777.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@157781.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@157775.4]
  assign regs_450_clock = clock; // @[:@157784.4]
  assign regs_450_reset = io_reset; // @[:@157785.4 RegFile.scala 76:16:@157792.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@157791.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@157795.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@157789.4]
  assign regs_451_clock = clock; // @[:@157798.4]
  assign regs_451_reset = io_reset; // @[:@157799.4 RegFile.scala 76:16:@157806.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@157805.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@157809.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@157803.4]
  assign regs_452_clock = clock; // @[:@157812.4]
  assign regs_452_reset = io_reset; // @[:@157813.4 RegFile.scala 76:16:@157820.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@157819.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@157823.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@157817.4]
  assign regs_453_clock = clock; // @[:@157826.4]
  assign regs_453_reset = io_reset; // @[:@157827.4 RegFile.scala 76:16:@157834.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@157833.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@157837.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@157831.4]
  assign regs_454_clock = clock; // @[:@157840.4]
  assign regs_454_reset = io_reset; // @[:@157841.4 RegFile.scala 76:16:@157848.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@157847.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@157851.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@157845.4]
  assign regs_455_clock = clock; // @[:@157854.4]
  assign regs_455_reset = io_reset; // @[:@157855.4 RegFile.scala 76:16:@157862.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@157861.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@157865.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@157859.4]
  assign regs_456_clock = clock; // @[:@157868.4]
  assign regs_456_reset = io_reset; // @[:@157869.4 RegFile.scala 76:16:@157876.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@157875.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@157879.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@157873.4]
  assign regs_457_clock = clock; // @[:@157882.4]
  assign regs_457_reset = io_reset; // @[:@157883.4 RegFile.scala 76:16:@157890.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@157889.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@157893.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@157887.4]
  assign regs_458_clock = clock; // @[:@157896.4]
  assign regs_458_reset = io_reset; // @[:@157897.4 RegFile.scala 76:16:@157904.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@157903.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@157907.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@157901.4]
  assign regs_459_clock = clock; // @[:@157910.4]
  assign regs_459_reset = io_reset; // @[:@157911.4 RegFile.scala 76:16:@157918.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@157917.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@157921.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@157915.4]
  assign regs_460_clock = clock; // @[:@157924.4]
  assign regs_460_reset = io_reset; // @[:@157925.4 RegFile.scala 76:16:@157932.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@157931.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@157935.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@157929.4]
  assign regs_461_clock = clock; // @[:@157938.4]
  assign regs_461_reset = io_reset; // @[:@157939.4 RegFile.scala 76:16:@157946.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@157945.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@157949.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@157943.4]
  assign regs_462_clock = clock; // @[:@157952.4]
  assign regs_462_reset = io_reset; // @[:@157953.4 RegFile.scala 76:16:@157960.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@157959.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@157963.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@157957.4]
  assign regs_463_clock = clock; // @[:@157966.4]
  assign regs_463_reset = io_reset; // @[:@157967.4 RegFile.scala 76:16:@157974.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@157973.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@157977.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@157971.4]
  assign regs_464_clock = clock; // @[:@157980.4]
  assign regs_464_reset = io_reset; // @[:@157981.4 RegFile.scala 76:16:@157988.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@157987.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@157991.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@157985.4]
  assign regs_465_clock = clock; // @[:@157994.4]
  assign regs_465_reset = io_reset; // @[:@157995.4 RegFile.scala 76:16:@158002.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@158001.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@158005.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@157999.4]
  assign regs_466_clock = clock; // @[:@158008.4]
  assign regs_466_reset = io_reset; // @[:@158009.4 RegFile.scala 76:16:@158016.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@158015.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@158019.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@158013.4]
  assign regs_467_clock = clock; // @[:@158022.4]
  assign regs_467_reset = io_reset; // @[:@158023.4 RegFile.scala 76:16:@158030.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@158029.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@158033.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@158027.4]
  assign regs_468_clock = clock; // @[:@158036.4]
  assign regs_468_reset = io_reset; // @[:@158037.4 RegFile.scala 76:16:@158044.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@158043.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@158047.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@158041.4]
  assign regs_469_clock = clock; // @[:@158050.4]
  assign regs_469_reset = io_reset; // @[:@158051.4 RegFile.scala 76:16:@158058.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@158057.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@158061.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@158055.4]
  assign regs_470_clock = clock; // @[:@158064.4]
  assign regs_470_reset = io_reset; // @[:@158065.4 RegFile.scala 76:16:@158072.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@158071.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@158075.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@158069.4]
  assign regs_471_clock = clock; // @[:@158078.4]
  assign regs_471_reset = io_reset; // @[:@158079.4 RegFile.scala 76:16:@158086.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@158085.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@158089.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@158083.4]
  assign regs_472_clock = clock; // @[:@158092.4]
  assign regs_472_reset = io_reset; // @[:@158093.4 RegFile.scala 76:16:@158100.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@158099.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@158103.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@158097.4]
  assign regs_473_clock = clock; // @[:@158106.4]
  assign regs_473_reset = io_reset; // @[:@158107.4 RegFile.scala 76:16:@158114.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@158113.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@158117.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@158111.4]
  assign regs_474_clock = clock; // @[:@158120.4]
  assign regs_474_reset = io_reset; // @[:@158121.4 RegFile.scala 76:16:@158128.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@158127.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@158131.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@158125.4]
  assign regs_475_clock = clock; // @[:@158134.4]
  assign regs_475_reset = io_reset; // @[:@158135.4 RegFile.scala 76:16:@158142.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@158141.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@158145.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@158139.4]
  assign regs_476_clock = clock; // @[:@158148.4]
  assign regs_476_reset = io_reset; // @[:@158149.4 RegFile.scala 76:16:@158156.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@158155.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@158159.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@158153.4]
  assign regs_477_clock = clock; // @[:@158162.4]
  assign regs_477_reset = io_reset; // @[:@158163.4 RegFile.scala 76:16:@158170.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@158169.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@158173.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@158167.4]
  assign regs_478_clock = clock; // @[:@158176.4]
  assign regs_478_reset = io_reset; // @[:@158177.4 RegFile.scala 76:16:@158184.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@158183.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@158187.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@158181.4]
  assign regs_479_clock = clock; // @[:@158190.4]
  assign regs_479_reset = io_reset; // @[:@158191.4 RegFile.scala 76:16:@158198.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@158197.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@158201.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@158195.4]
  assign regs_480_clock = clock; // @[:@158204.4]
  assign regs_480_reset = io_reset; // @[:@158205.4 RegFile.scala 76:16:@158212.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@158211.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@158215.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@158209.4]
  assign regs_481_clock = clock; // @[:@158218.4]
  assign regs_481_reset = io_reset; // @[:@158219.4 RegFile.scala 76:16:@158226.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@158225.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@158229.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@158223.4]
  assign regs_482_clock = clock; // @[:@158232.4]
  assign regs_482_reset = io_reset; // @[:@158233.4 RegFile.scala 76:16:@158240.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@158239.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@158243.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@158237.4]
  assign regs_483_clock = clock; // @[:@158246.4]
  assign regs_483_reset = io_reset; // @[:@158247.4 RegFile.scala 76:16:@158254.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@158253.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@158257.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@158251.4]
  assign regs_484_clock = clock; // @[:@158260.4]
  assign regs_484_reset = io_reset; // @[:@158261.4 RegFile.scala 76:16:@158268.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@158267.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@158271.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@158265.4]
  assign regs_485_clock = clock; // @[:@158274.4]
  assign regs_485_reset = io_reset; // @[:@158275.4 RegFile.scala 76:16:@158282.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@158281.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@158285.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@158279.4]
  assign regs_486_clock = clock; // @[:@158288.4]
  assign regs_486_reset = io_reset; // @[:@158289.4 RegFile.scala 76:16:@158296.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@158295.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@158299.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@158293.4]
  assign regs_487_clock = clock; // @[:@158302.4]
  assign regs_487_reset = io_reset; // @[:@158303.4 RegFile.scala 76:16:@158310.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@158309.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@158313.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@158307.4]
  assign regs_488_clock = clock; // @[:@158316.4]
  assign regs_488_reset = io_reset; // @[:@158317.4 RegFile.scala 76:16:@158324.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@158323.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@158327.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@158321.4]
  assign regs_489_clock = clock; // @[:@158330.4]
  assign regs_489_reset = io_reset; // @[:@158331.4 RegFile.scala 76:16:@158338.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@158337.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@158341.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@158335.4]
  assign regs_490_clock = clock; // @[:@158344.4]
  assign regs_490_reset = io_reset; // @[:@158345.4 RegFile.scala 76:16:@158352.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@158351.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@158355.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@158349.4]
  assign regs_491_clock = clock; // @[:@158358.4]
  assign regs_491_reset = io_reset; // @[:@158359.4 RegFile.scala 76:16:@158366.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@158365.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@158369.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@158363.4]
  assign regs_492_clock = clock; // @[:@158372.4]
  assign regs_492_reset = io_reset; // @[:@158373.4 RegFile.scala 76:16:@158380.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@158379.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@158383.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@158377.4]
  assign regs_493_clock = clock; // @[:@158386.4]
  assign regs_493_reset = io_reset; // @[:@158387.4 RegFile.scala 76:16:@158394.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@158393.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@158397.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@158391.4]
  assign regs_494_clock = clock; // @[:@158400.4]
  assign regs_494_reset = io_reset; // @[:@158401.4 RegFile.scala 76:16:@158408.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@158407.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@158411.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@158405.4]
  assign regs_495_clock = clock; // @[:@158414.4]
  assign regs_495_reset = io_reset; // @[:@158415.4 RegFile.scala 76:16:@158422.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@158421.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@158425.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@158419.4]
  assign regs_496_clock = clock; // @[:@158428.4]
  assign regs_496_reset = io_reset; // @[:@158429.4 RegFile.scala 76:16:@158436.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@158435.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@158439.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@158433.4]
  assign regs_497_clock = clock; // @[:@158442.4]
  assign regs_497_reset = io_reset; // @[:@158443.4 RegFile.scala 76:16:@158450.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@158449.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@158453.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@158447.4]
  assign regs_498_clock = clock; // @[:@158456.4]
  assign regs_498_reset = io_reset; // @[:@158457.4 RegFile.scala 76:16:@158464.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@158463.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@158467.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@158461.4]
  assign regs_499_clock = clock; // @[:@158470.4]
  assign regs_499_reset = io_reset; // @[:@158471.4 RegFile.scala 76:16:@158478.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@158477.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@158481.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@158475.4]
  assign regs_500_clock = clock; // @[:@158484.4]
  assign regs_500_reset = io_reset; // @[:@158485.4 RegFile.scala 76:16:@158492.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@158491.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@158495.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@158489.4]
  assign regs_501_clock = clock; // @[:@158498.4]
  assign regs_501_reset = io_reset; // @[:@158499.4 RegFile.scala 76:16:@158506.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@158505.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@158509.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@158503.4]
  assign regs_502_clock = clock; // @[:@158512.4]
  assign regs_502_reset = io_reset; // @[:@158513.4 RegFile.scala 76:16:@158520.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@158519.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@158523.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@158517.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@159032.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@159033.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@159034.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@159035.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@159036.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@159037.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@159038.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@159039.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@159040.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@159041.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@159042.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@159043.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@159044.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@159045.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@159046.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@159047.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@159048.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@159049.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@159050.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@159051.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@159052.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@159053.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@159054.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@159055.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@159056.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@159057.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@159058.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@159059.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@159060.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@159061.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@159062.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@159063.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@159064.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@159065.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@159066.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@159067.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@159068.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@159069.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@159070.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@159071.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@159072.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@159073.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@159074.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@159075.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@159076.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@159077.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@159078.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@159079.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@159080.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@159081.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@159082.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@159083.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@159084.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@159085.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@159086.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@159087.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@159088.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@159089.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@159090.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@159091.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@159092.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@159093.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@159094.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@159095.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@159096.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@159097.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@159098.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@159099.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@159100.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@159101.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@159102.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@159103.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@159104.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@159105.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@159106.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@159107.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@159108.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@159109.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@159110.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@159111.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@159112.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@159113.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@159114.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@159115.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@159116.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@159117.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@159118.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@159119.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@159120.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@159121.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@159122.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@159123.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@159124.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@159125.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@159126.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@159127.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@159128.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@159129.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@159130.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@159131.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@159132.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@159133.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@159134.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@159135.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@159136.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@159137.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@159138.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@159139.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@159140.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@159141.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@159142.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@159143.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@159144.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@159145.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@159146.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@159147.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@159148.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@159149.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@159150.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@159151.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@159152.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@159153.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@159154.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@159155.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@159156.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@159157.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@159158.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@159159.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@159160.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@159161.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@159162.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@159163.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@159164.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@159165.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@159166.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@159167.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@159168.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@159169.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@159170.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@159171.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@159172.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@159173.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@159174.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@159175.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@159176.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@159177.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@159178.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@159179.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@159180.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@159181.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@159182.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@159183.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@159184.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@159185.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@159186.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@159187.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@159188.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@159189.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@159190.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@159191.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@159192.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@159193.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@159194.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@159195.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@159196.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@159197.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@159198.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@159199.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@159200.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@159201.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@159202.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@159203.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@159204.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@159205.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@159206.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@159207.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@159208.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@159209.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@159210.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@159211.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@159212.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@159213.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@159214.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@159215.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@159216.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@159217.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@159218.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@159219.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@159220.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@159221.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@159222.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@159223.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@159224.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@159225.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@159226.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@159227.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@159228.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@159229.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@159230.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@159231.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@159232.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@159233.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@159234.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@159235.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@159236.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@159237.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@159238.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@159239.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@159240.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@159241.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@159242.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@159243.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@159244.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@159245.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@159246.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@159247.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@159248.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@159249.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@159250.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@159251.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@159252.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@159253.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@159254.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@159255.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@159256.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@159257.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@159258.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@159259.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@159260.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@159261.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@159262.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@159263.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@159264.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@159265.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@159266.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@159267.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@159268.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@159269.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@159270.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@159271.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@159272.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@159273.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@159274.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@159275.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@159276.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@159277.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@159278.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@159279.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@159280.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@159281.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@159282.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@159283.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@159284.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@159285.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@159286.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@159287.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@159288.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@159289.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@159290.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@159291.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@159292.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@159293.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@159294.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@159295.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@159296.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@159297.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@159298.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@159299.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@159300.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@159301.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@159302.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@159303.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@159304.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@159305.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@159306.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@159307.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@159308.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@159309.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@159310.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@159311.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@159312.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@159313.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@159314.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@159315.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@159316.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@159317.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@159318.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@159319.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@159320.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@159321.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@159322.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@159323.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@159324.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@159325.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@159326.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@159327.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@159328.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@159329.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@159330.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@159331.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@159332.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@159333.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@159334.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@159335.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@159336.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@159337.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@159338.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@159339.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@159340.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@159341.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@159342.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@159343.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@159344.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@159345.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@159346.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@159347.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@159348.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@159349.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@159350.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@159351.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@159352.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@159353.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@159354.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@159355.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@159356.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@159357.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@159358.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@159359.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@159360.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@159361.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@159362.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@159363.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@159364.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@159365.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@159366.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@159367.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@159368.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@159369.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@159370.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@159371.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@159372.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@159373.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@159374.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@159375.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@159376.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@159377.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@159378.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@159379.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@159380.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@159381.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@159382.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@159383.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@159384.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@159385.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@159386.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@159387.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@159388.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@159389.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@159390.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@159391.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@159392.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@159393.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@159394.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@159395.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@159396.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@159397.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@159398.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@159399.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@159400.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@159401.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@159402.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@159403.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@159404.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@159405.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@159406.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@159407.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@159408.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@159409.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@159410.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@159411.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@159412.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@159413.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@159414.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@159415.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@159416.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@159417.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@159418.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@159419.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@159420.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@159421.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@159422.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@159423.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@159424.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@159425.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@159426.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@159427.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@159428.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@159429.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@159430.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@159431.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@159432.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@159433.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@159434.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@159435.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@159436.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@159437.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@159438.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@159439.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@159440.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@159441.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@159442.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@159443.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@159444.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@159445.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@159446.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@159447.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@159448.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@159449.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@159450.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@159451.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@159452.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@159453.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@159454.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@159455.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@159456.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@159457.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@159458.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@159459.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@159460.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@159461.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@159462.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@159463.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@159464.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@159465.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@159466.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@159467.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@159468.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@159469.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@159470.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@159471.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@159472.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@159473.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@159474.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@159475.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@159476.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@159477.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@159478.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@159479.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@159480.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@159481.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@159482.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@159483.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@159484.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@159485.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@159486.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@159487.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@159488.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@159489.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@159490.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@159491.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@159492.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@159493.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@159494.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@159495.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@159496.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@159497.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@159498.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@159499.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@159500.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@159501.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@159502.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@159503.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@159504.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@159505.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@159506.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@159507.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@159508.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@159509.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@159510.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@159511.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@159512.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@159513.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@159514.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@159515.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@159516.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@159517.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@159518.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@159519.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@159520.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@159521.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@159522.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@159523.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@159524.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@159525.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@159526.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@159527.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@159528.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@159529.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@159530.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@159531.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@159532.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@159533.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@159534.4]
  assign rport_io_sel = _T_7111[8:0]; // @[RegFile.scala 99:18:@159536.4]
endmodule
module RetimeWrapper_1304( // @[:@159560.2]
  input         clock, // @[:@159561.4]
  input         reset, // @[:@159562.4]
  input  [39:0] io_in, // @[:@159563.4]
  output [39:0] io_out // @[:@159563.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@159565.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@159565.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@159565.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@159565.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@159565.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@159565.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@159565.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@159578.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@159577.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@159576.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@159575.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@159574.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@159572.4]
endmodule
module FringeFF_503( // @[:@159580.2]
  input         clock, // @[:@159581.4]
  input         reset, // @[:@159582.4]
  input  [39:0] io_in, // @[:@159583.4]
  output [39:0] io_out, // @[:@159583.4]
  input         io_enable // @[:@159583.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@159586.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@159586.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@159586.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@159586.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@159591.4 package.scala 96:25:@159592.4]
  RetimeWrapper_1304 RetimeWrapper ( // @[package.scala 93:22:@159586.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@159591.4 package.scala 96:25:@159592.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@159603.4]
  assign RetimeWrapper_clock = clock; // @[:@159587.4]
  assign RetimeWrapper_reset = reset; // @[:@159588.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@159589.4]
endmodule
module FringeCounter( // @[:@159605.2]
  input   clock, // @[:@159606.4]
  input   reset, // @[:@159607.4]
  input   io_enable, // @[:@159608.4]
  output  io_done // @[:@159608.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@159610.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@159610.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@159610.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@159610.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@159610.4]
  wire [40:0] count; // @[Cat.scala 30:58:@159617.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@159618.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@159619.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@159620.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@159622.4]
  FringeFF_503 reg$ ( // @[FringeCounter.scala 24:19:@159610.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@159617.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@159618.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@159619.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@159620.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@159622.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@159633.4]
  assign reg$_clock = clock; // @[:@159611.4]
  assign reg$_reset = reset; // @[:@159612.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@159624.6 FringeCounter.scala 37:15:@159627.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@159615.4]
endmodule
module FringeFF_504( // @[:@159667.2]
  input   clock, // @[:@159668.4]
  input   reset, // @[:@159669.4]
  input   io_in, // @[:@159670.4]
  input   io_reset, // @[:@159670.4]
  output  io_out, // @[:@159670.4]
  input   io_enable // @[:@159670.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@159673.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@159673.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@159673.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@159673.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@159673.4]
  wire  _T_18; // @[package.scala 96:25:@159678.4 package.scala 96:25:@159679.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@159684.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@159673.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@159678.4 package.scala 96:25:@159679.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@159684.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@159690.4]
  assign RetimeWrapper_clock = clock; // @[:@159674.4]
  assign RetimeWrapper_reset = reset; // @[:@159675.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@159677.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@159676.4]
endmodule
module Depulser( // @[:@159692.2]
  input   clock, // @[:@159693.4]
  input   reset, // @[:@159694.4]
  input   io_in, // @[:@159695.4]
  input   io_rst, // @[:@159695.4]
  output  io_out // @[:@159695.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@159697.4]
  wire  r_reset; // @[Depulser.scala 14:17:@159697.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@159697.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@159697.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@159697.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@159697.4]
  FringeFF_504 r ( // @[Depulser.scala 14:17:@159697.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@159706.4]
  assign r_clock = clock; // @[:@159698.4]
  assign r_reset = reset; // @[:@159699.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@159701.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@159705.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@159704.4]
endmodule
module Fringe( // @[:@159708.2]
  input         clock, // @[:@159709.4]
  input         reset, // @[:@159710.4]
  input  [39:0] io_raddr, // @[:@159711.4]
  input         io_wen, // @[:@159711.4]
  input  [39:0] io_waddr, // @[:@159711.4]
  input  [63:0] io_wdata, // @[:@159711.4]
  output [63:0] io_rdata, // @[:@159711.4]
  output        io_enable, // @[:@159711.4]
  input         io_done, // @[:@159711.4]
  output        io_reset, // @[:@159711.4]
  output [63:0] io_argIns_0, // @[:@159711.4]
  output [63:0] io_argIns_1, // @[:@159711.4]
  input         io_argOuts_0_valid, // @[:@159711.4]
  input  [63:0] io_argOuts_0_bits, // @[:@159711.4]
  output [63:0] io_argEchos_0, // @[:@159711.4]
  output        io_memStreams_loads_0_cmd_ready, // @[:@159711.4]
  input         io_memStreams_loads_0_cmd_valid, // @[:@159711.4]
  input  [63:0] io_memStreams_loads_0_cmd_bits_addr, // @[:@159711.4]
  input  [31:0] io_memStreams_loads_0_cmd_bits_size, // @[:@159711.4]
  input         io_memStreams_loads_0_data_ready, // @[:@159711.4]
  output        io_memStreams_loads_0_data_valid, // @[:@159711.4]
  output [31:0] io_memStreams_loads_0_data_bits_rdata_0, // @[:@159711.4]
  output        io_memStreams_stores_0_cmd_ready, // @[:@159711.4]
  input         io_memStreams_stores_0_cmd_valid, // @[:@159711.4]
  input  [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@159711.4]
  input  [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@159711.4]
  output        io_memStreams_stores_0_data_ready, // @[:@159711.4]
  input         io_memStreams_stores_0_data_valid, // @[:@159711.4]
  input  [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@159711.4]
  input         io_memStreams_stores_0_data_bits_wstrb, // @[:@159711.4]
  input         io_memStreams_stores_0_wresp_ready, // @[:@159711.4]
  output        io_memStreams_stores_0_wresp_valid, // @[:@159711.4]
  output        io_memStreams_stores_0_wresp_bits, // @[:@159711.4]
  input         io_dram_0_cmd_ready, // @[:@159711.4]
  output        io_dram_0_cmd_valid, // @[:@159711.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@159711.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@159711.4]
  output        io_dram_0_cmd_bits_isWr, // @[:@159711.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@159711.4]
  input         io_dram_0_wdata_ready, // @[:@159711.4]
  output        io_dram_0_wdata_valid, // @[:@159711.4]
  output [63:0] io_dram_0_wdata_bits_wdata_0, // @[:@159711.4]
  output [63:0] io_dram_0_wdata_bits_wdata_1, // @[:@159711.4]
  output [63:0] io_dram_0_wdata_bits_wdata_2, // @[:@159711.4]
  output [63:0] io_dram_0_wdata_bits_wdata_3, // @[:@159711.4]
  output [63:0] io_dram_0_wdata_bits_wdata_4, // @[:@159711.4]
  output [63:0] io_dram_0_wdata_bits_wdata_5, // @[:@159711.4]
  output [63:0] io_dram_0_wdata_bits_wdata_6, // @[:@159711.4]
  output [63:0] io_dram_0_wdata_bits_wdata_7, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_0, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_1, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_2, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_3, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_4, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_5, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_6, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_7, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_8, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_9, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_10, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_11, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_12, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_13, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_14, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_15, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_16, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_17, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_18, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_19, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_20, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_21, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_22, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_23, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_24, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_25, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_26, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_27, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_28, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_29, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_30, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_31, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_32, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_33, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_34, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_35, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_36, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_37, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_38, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_39, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_40, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_41, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_42, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_43, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_44, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_45, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_46, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_47, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_48, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_49, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_50, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_51, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_52, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_53, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_54, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_55, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_56, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_57, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_58, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_59, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_60, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_61, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_62, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wstrb_63, // @[:@159711.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@159711.4]
  output        io_dram_0_rresp_ready, // @[:@159711.4]
  input         io_dram_0_rresp_valid, // @[:@159711.4]
  input  [63:0] io_dram_0_rresp_bits_rdata_0, // @[:@159711.4]
  input  [63:0] io_dram_0_rresp_bits_rdata_1, // @[:@159711.4]
  input  [63:0] io_dram_0_rresp_bits_rdata_2, // @[:@159711.4]
  input  [63:0] io_dram_0_rresp_bits_rdata_3, // @[:@159711.4]
  input  [63:0] io_dram_0_rresp_bits_rdata_4, // @[:@159711.4]
  input  [63:0] io_dram_0_rresp_bits_rdata_5, // @[:@159711.4]
  input  [63:0] io_dram_0_rresp_bits_rdata_6, // @[:@159711.4]
  input  [63:0] io_dram_0_rresp_bits_rdata_7, // @[:@159711.4]
  input  [31:0] io_dram_0_rresp_bits_tag, // @[:@159711.4]
  output        io_dram_0_wresp_ready, // @[:@159711.4]
  input         io_dram_0_wresp_valid, // @[:@159711.4]
  input  [31:0] io_dram_0_wresp_bits_tag, // @[:@159711.4]
  input         io_dram_1_cmd_ready, // @[:@159711.4]
  output        io_dram_1_cmd_valid, // @[:@159711.4]
  output [63:0] io_dram_1_cmd_bits_addr, // @[:@159711.4]
  output [31:0] io_dram_1_cmd_bits_size, // @[:@159711.4]
  output        io_dram_1_cmd_bits_isWr, // @[:@159711.4]
  output [31:0] io_dram_1_cmd_bits_tag, // @[:@159711.4]
  input         io_dram_1_wdata_ready, // @[:@159711.4]
  output        io_dram_1_wdata_valid, // @[:@159711.4]
  output [63:0] io_dram_1_wdata_bits_wdata_0, // @[:@159711.4]
  output [63:0] io_dram_1_wdata_bits_wdata_1, // @[:@159711.4]
  output [63:0] io_dram_1_wdata_bits_wdata_2, // @[:@159711.4]
  output [63:0] io_dram_1_wdata_bits_wdata_3, // @[:@159711.4]
  output [63:0] io_dram_1_wdata_bits_wdata_4, // @[:@159711.4]
  output [63:0] io_dram_1_wdata_bits_wdata_5, // @[:@159711.4]
  output [63:0] io_dram_1_wdata_bits_wdata_6, // @[:@159711.4]
  output [63:0] io_dram_1_wdata_bits_wdata_7, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_0, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_1, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_2, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_3, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_4, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_5, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_6, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_7, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_8, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_9, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_10, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_11, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_12, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_13, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_14, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_15, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_16, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_17, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_18, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_19, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_20, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_21, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_22, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_23, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_24, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_25, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_26, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_27, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_28, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_29, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_30, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_31, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_32, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_33, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_34, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_35, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_36, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_37, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_38, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_39, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_40, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_41, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_42, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_43, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_44, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_45, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_46, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_47, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_48, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_49, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_50, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_51, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_52, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_53, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_54, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_55, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_56, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_57, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_58, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_59, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_60, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_61, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_62, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wstrb_63, // @[:@159711.4]
  output        io_dram_1_wdata_bits_wlast, // @[:@159711.4]
  output        io_dram_1_rresp_ready, // @[:@159711.4]
  input         io_dram_1_rresp_valid, // @[:@159711.4]
  input  [63:0] io_dram_1_rresp_bits_rdata_0, // @[:@159711.4]
  input  [63:0] io_dram_1_rresp_bits_rdata_1, // @[:@159711.4]
  input  [63:0] io_dram_1_rresp_bits_rdata_2, // @[:@159711.4]
  input  [63:0] io_dram_1_rresp_bits_rdata_3, // @[:@159711.4]
  input  [63:0] io_dram_1_rresp_bits_rdata_4, // @[:@159711.4]
  input  [63:0] io_dram_1_rresp_bits_rdata_5, // @[:@159711.4]
  input  [63:0] io_dram_1_rresp_bits_rdata_6, // @[:@159711.4]
  input  [63:0] io_dram_1_rresp_bits_rdata_7, // @[:@159711.4]
  input  [31:0] io_dram_1_rresp_bits_tag, // @[:@159711.4]
  output        io_dram_1_wresp_ready, // @[:@159711.4]
  input         io_dram_1_wresp_valid, // @[:@159711.4]
  input  [31:0] io_dram_1_wresp_bits_tag, // @[:@159711.4]
  input         io_heap_0_req_valid, // @[:@159711.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@159711.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@159711.4]
  output        io_heap_0_resp_valid, // @[:@159711.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@159711.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@159711.4]
);
  wire  dramArbs_0_clock; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_reset; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_enable; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_app_loads_0_cmd_ready; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_app_loads_0_cmd_valid; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_app_loads_0_cmd_bits_addr; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_app_loads_0_cmd_bits_size; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_app_loads_0_data_ready; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_app_loads_0_data_valid; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_app_loads_0_data_bits_rdata_0; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_app_stores_0_cmd_valid; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_app_stores_0_cmd_bits_addr; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_app_stores_0_cmd_bits_size; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_app_stores_0_data_valid; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_app_stores_0_data_bits_wdata_0; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_app_stores_0_data_bits_wstrb; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_app_stores_0_wresp_ready; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_cmd_ready; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_ready; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_rresp_valid; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_rresp_bits_rdata_0; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_rresp_bits_rdata_1; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_rresp_bits_rdata_2; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_rresp_bits_rdata_3; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_rresp_bits_rdata_4; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_rresp_bits_rdata_5; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_rresp_bits_rdata_6; // @[Fringe.scala 91:25:@159717.4]
  wire [63:0] dramArbs_0_io_dram_rresp_bits_rdata_7; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_dram_rresp_bits_tag; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_0_io_dram_wresp_valid; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_0; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_1; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_2; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_3; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_4; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_5; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_6; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_7; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_8; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_9; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_10; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_11; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_12; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_13; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_14; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_15; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_16; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_17; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_18; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_19; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_20; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_21; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_22; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_23; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_24; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_25; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_26; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_27; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_28; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_29; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_30; // @[Fringe.scala 91:25:@159717.4]
  wire [31:0] dramArbs_0_io_debugSignals_41; // @[Fringe.scala 91:25:@159717.4]
  wire  dramArbs_1_clock; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_reset; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_enable; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_app_loads_0_cmd_ready; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_app_loads_0_cmd_valid; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_app_loads_0_cmd_bits_addr; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_app_loads_0_cmd_bits_size; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_app_loads_0_data_ready; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_app_loads_0_data_valid; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_app_loads_0_data_bits_rdata_0; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_app_stores_0_cmd_ready; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_app_stores_0_cmd_valid; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_app_stores_0_cmd_bits_addr; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_app_stores_0_cmd_bits_size; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_app_stores_0_data_ready; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_app_stores_0_data_valid; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_app_stores_0_data_bits_wdata_0; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_app_stores_0_data_bits_wstrb; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_app_stores_0_wresp_ready; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_app_stores_0_wresp_valid; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_app_stores_0_wresp_bits; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_cmd_ready; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_ready; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_rresp_valid; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_rresp_bits_rdata_0; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_rresp_bits_rdata_1; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_rresp_bits_rdata_2; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_rresp_bits_rdata_3; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_rresp_bits_rdata_4; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_rresp_bits_rdata_5; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_rresp_bits_rdata_6; // @[Fringe.scala 91:25:@160600.4]
  wire [63:0] dramArbs_1_io_dram_rresp_bits_rdata_7; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_dram_rresp_bits_tag; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 91:25:@160600.4]
  wire  dramArbs_1_io_dram_wresp_valid; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_0; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_1; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_2; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_3; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_4; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_5; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_6; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_7; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_8; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_9; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_10; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_11; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_12; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_13; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_14; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_15; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_16; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_17; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_18; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_19; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_20; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_21; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_22; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_23; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_24; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_25; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_26; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_27; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_28; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_29; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_30; // @[Fringe.scala 91:25:@160600.4]
  wire [31:0] dramArbs_1_io_debugSignals_41; // @[Fringe.scala 91:25:@160600.4]
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@161465.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@161465.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@161465.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@161465.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@161465.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@161465.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@161465.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@161465.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@161465.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@161465.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@161465.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@161465.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@161474.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@161474.4]
  wire [39:0] regs_io_raddr; // @[Fringe.scala 116:20:@161474.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@161474.4]
  wire [39:0] regs_io_waddr; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@161474.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argIns_3; // @[Fringe.scala 116:20:@161474.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@161474.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_2_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_3_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_4_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_5_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_6_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_7_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_8_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_9_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_10_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_11_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_12_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_13_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_14_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_15_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_16_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_17_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_18_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_19_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_20_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_21_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_22_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_23_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_24_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_25_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_26_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_27_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_28_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_29_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_30_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_31_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_32_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argOuts_43_bits; // @[Fringe.scala 116:20:@161474.4]
  wire [63:0] regs_io_argEchos_1; // @[Fringe.scala 116:20:@161474.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@163524.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@163524.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@163524.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@163524.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@163543.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@163543.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@163543.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@163543.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@163543.4]
  wire [63:0] _T_548; // @[:@163501.4 :@163502.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@163503.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@163505.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@163507.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@163509.4]
  wire  _T_553; // @[Fringe.scala 134:60:@163511.4]
  wire  _T_557; // @[Fringe.scala 134:74:@163513.4]
  wire  _T_558; // @[Fringe.scala 135:27:@163515.4]
  wire [63:0] _T_568; // @[Fringe.scala 156:22:@163551.4]
  reg  _T_575; // @[package.scala 152:20:@163554.4]
  reg [31:0] _RAND_0;
  wire  _T_576; // @[package.scala 153:13:@163556.4]
  wire  _T_577; // @[package.scala 153:8:@163557.4]
  wire  _T_580; // @[Fringe.scala 160:55:@163561.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@163562.4]
  wire  _T_583; // @[Fringe.scala 161:58:@163565.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@163566.4]
  wire [1:0] _T_587; // @[Fringe.scala 162:57:@163568.4]
  wire [1:0] _T_589; // @[Fringe.scala 162:34:@163569.4]
  wire [63:0] _T_591; // @[Fringe.scala 163:30:@163571.4]
  wire [1:0] _T_592; // @[Fringe.scala 171:37:@163574.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@163553.4 Fringe.scala 163:24:@163572.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@163553.4 Fringe.scala 162:28:@163570.4]
  wire [61:0] _T_593; // @[Fringe.scala 171:37:@163575.4]
  wire  alloc; // @[Fringe.scala 202:38:@164779.4]
  wire  dealloc; // @[Fringe.scala 203:40:@164780.4]
  wire  _T_1097; // @[Fringe.scala 204:37:@164781.4]
  reg  _T_1100; // @[package.scala 152:20:@164782.4]
  reg [31:0] _RAND_1;
  wire  _T_1101; // @[package.scala 153:13:@164784.4]
  DRAMArbiter dramArbs_0 ( // @[Fringe.scala 91:25:@159717.4]
    .clock(dramArbs_0_clock),
    .reset(dramArbs_0_reset),
    .io_enable(dramArbs_0_io_enable),
    .io_app_loads_0_cmd_ready(dramArbs_0_io_app_loads_0_cmd_ready),
    .io_app_loads_0_cmd_valid(dramArbs_0_io_app_loads_0_cmd_valid),
    .io_app_loads_0_cmd_bits_addr(dramArbs_0_io_app_loads_0_cmd_bits_addr),
    .io_app_loads_0_cmd_bits_size(dramArbs_0_io_app_loads_0_cmd_bits_size),
    .io_app_loads_0_data_ready(dramArbs_0_io_app_loads_0_data_ready),
    .io_app_loads_0_data_valid(dramArbs_0_io_app_loads_0_data_valid),
    .io_app_loads_0_data_bits_rdata_0(dramArbs_0_io_app_loads_0_data_bits_rdata_0),
    .io_app_stores_0_cmd_ready(dramArbs_0_io_app_stores_0_cmd_ready),
    .io_app_stores_0_cmd_valid(dramArbs_0_io_app_stores_0_cmd_valid),
    .io_app_stores_0_cmd_bits_addr(dramArbs_0_io_app_stores_0_cmd_bits_addr),
    .io_app_stores_0_cmd_bits_size(dramArbs_0_io_app_stores_0_cmd_bits_size),
    .io_app_stores_0_data_ready(dramArbs_0_io_app_stores_0_data_ready),
    .io_app_stores_0_data_valid(dramArbs_0_io_app_stores_0_data_valid),
    .io_app_stores_0_data_bits_wdata_0(dramArbs_0_io_app_stores_0_data_bits_wdata_0),
    .io_app_stores_0_data_bits_wstrb(dramArbs_0_io_app_stores_0_data_bits_wstrb),
    .io_app_stores_0_wresp_ready(dramArbs_0_io_app_stores_0_wresp_ready),
    .io_app_stores_0_wresp_valid(dramArbs_0_io_app_stores_0_wresp_valid),
    .io_app_stores_0_wresp_bits(dramArbs_0_io_app_stores_0_wresp_bits),
    .io_dram_cmd_ready(dramArbs_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_0_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_0_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_0_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_0_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_0_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_0_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_0_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_0_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wstrb_0(dramArbs_0_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_0_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_0_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_0_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_0_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_0_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_0_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_0_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_0_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_0_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_0_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_0_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_0_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_0_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_0_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_0_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_0_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_0_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_0_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_0_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_0_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_0_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_0_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_0_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_0_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_0_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_0_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_0_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_0_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_0_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_0_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_0_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_0_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_0_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_0_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_0_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_0_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_0_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_0_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_0_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_0_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_0_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_0_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_0_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_0_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_0_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_0_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_0_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_0_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_0_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_0_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_0_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_0_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_0_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_0_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_0_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_0_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_0_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_0_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_0_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_0_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_0_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_0_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_0_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_0_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_0_io_dram_rresp_ready),
    .io_dram_rresp_valid(dramArbs_0_io_dram_rresp_valid),
    .io_dram_rresp_bits_rdata_0(dramArbs_0_io_dram_rresp_bits_rdata_0),
    .io_dram_rresp_bits_rdata_1(dramArbs_0_io_dram_rresp_bits_rdata_1),
    .io_dram_rresp_bits_rdata_2(dramArbs_0_io_dram_rresp_bits_rdata_2),
    .io_dram_rresp_bits_rdata_3(dramArbs_0_io_dram_rresp_bits_rdata_3),
    .io_dram_rresp_bits_rdata_4(dramArbs_0_io_dram_rresp_bits_rdata_4),
    .io_dram_rresp_bits_rdata_5(dramArbs_0_io_dram_rresp_bits_rdata_5),
    .io_dram_rresp_bits_rdata_6(dramArbs_0_io_dram_rresp_bits_rdata_6),
    .io_dram_rresp_bits_rdata_7(dramArbs_0_io_dram_rresp_bits_rdata_7),
    .io_dram_rresp_bits_tag(dramArbs_0_io_dram_rresp_bits_tag),
    .io_dram_wresp_ready(dramArbs_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_0_io_dram_wresp_bits_tag),
    .io_debugSignals_0(dramArbs_0_io_debugSignals_0),
    .io_debugSignals_1(dramArbs_0_io_debugSignals_1),
    .io_debugSignals_2(dramArbs_0_io_debugSignals_2),
    .io_debugSignals_3(dramArbs_0_io_debugSignals_3),
    .io_debugSignals_4(dramArbs_0_io_debugSignals_4),
    .io_debugSignals_5(dramArbs_0_io_debugSignals_5),
    .io_debugSignals_6(dramArbs_0_io_debugSignals_6),
    .io_debugSignals_7(dramArbs_0_io_debugSignals_7),
    .io_debugSignals_8(dramArbs_0_io_debugSignals_8),
    .io_debugSignals_9(dramArbs_0_io_debugSignals_9),
    .io_debugSignals_10(dramArbs_0_io_debugSignals_10),
    .io_debugSignals_11(dramArbs_0_io_debugSignals_11),
    .io_debugSignals_12(dramArbs_0_io_debugSignals_12),
    .io_debugSignals_13(dramArbs_0_io_debugSignals_13),
    .io_debugSignals_14(dramArbs_0_io_debugSignals_14),
    .io_debugSignals_15(dramArbs_0_io_debugSignals_15),
    .io_debugSignals_16(dramArbs_0_io_debugSignals_16),
    .io_debugSignals_17(dramArbs_0_io_debugSignals_17),
    .io_debugSignals_18(dramArbs_0_io_debugSignals_18),
    .io_debugSignals_19(dramArbs_0_io_debugSignals_19),
    .io_debugSignals_20(dramArbs_0_io_debugSignals_20),
    .io_debugSignals_21(dramArbs_0_io_debugSignals_21),
    .io_debugSignals_22(dramArbs_0_io_debugSignals_22),
    .io_debugSignals_23(dramArbs_0_io_debugSignals_23),
    .io_debugSignals_24(dramArbs_0_io_debugSignals_24),
    .io_debugSignals_25(dramArbs_0_io_debugSignals_25),
    .io_debugSignals_26(dramArbs_0_io_debugSignals_26),
    .io_debugSignals_27(dramArbs_0_io_debugSignals_27),
    .io_debugSignals_28(dramArbs_0_io_debugSignals_28),
    .io_debugSignals_29(dramArbs_0_io_debugSignals_29),
    .io_debugSignals_30(dramArbs_0_io_debugSignals_30),
    .io_debugSignals_41(dramArbs_0_io_debugSignals_41)
  );
  DRAMArbiter dramArbs_1 ( // @[Fringe.scala 91:25:@160600.4]
    .clock(dramArbs_1_clock),
    .reset(dramArbs_1_reset),
    .io_enable(dramArbs_1_io_enable),
    .io_app_loads_0_cmd_ready(dramArbs_1_io_app_loads_0_cmd_ready),
    .io_app_loads_0_cmd_valid(dramArbs_1_io_app_loads_0_cmd_valid),
    .io_app_loads_0_cmd_bits_addr(dramArbs_1_io_app_loads_0_cmd_bits_addr),
    .io_app_loads_0_cmd_bits_size(dramArbs_1_io_app_loads_0_cmd_bits_size),
    .io_app_loads_0_data_ready(dramArbs_1_io_app_loads_0_data_ready),
    .io_app_loads_0_data_valid(dramArbs_1_io_app_loads_0_data_valid),
    .io_app_loads_0_data_bits_rdata_0(dramArbs_1_io_app_loads_0_data_bits_rdata_0),
    .io_app_stores_0_cmd_ready(dramArbs_1_io_app_stores_0_cmd_ready),
    .io_app_stores_0_cmd_valid(dramArbs_1_io_app_stores_0_cmd_valid),
    .io_app_stores_0_cmd_bits_addr(dramArbs_1_io_app_stores_0_cmd_bits_addr),
    .io_app_stores_0_cmd_bits_size(dramArbs_1_io_app_stores_0_cmd_bits_size),
    .io_app_stores_0_data_ready(dramArbs_1_io_app_stores_0_data_ready),
    .io_app_stores_0_data_valid(dramArbs_1_io_app_stores_0_data_valid),
    .io_app_stores_0_data_bits_wdata_0(dramArbs_1_io_app_stores_0_data_bits_wdata_0),
    .io_app_stores_0_data_bits_wstrb(dramArbs_1_io_app_stores_0_data_bits_wstrb),
    .io_app_stores_0_wresp_ready(dramArbs_1_io_app_stores_0_wresp_ready),
    .io_app_stores_0_wresp_valid(dramArbs_1_io_app_stores_0_wresp_valid),
    .io_app_stores_0_wresp_bits(dramArbs_1_io_app_stores_0_wresp_bits),
    .io_dram_cmd_ready(dramArbs_1_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_1_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_1_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_1_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_1_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_1_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_1_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_1_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_1_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_1_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_1_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_1_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_1_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_1_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_1_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_1_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wstrb_0(dramArbs_1_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_1_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_1_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_1_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_1_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_1_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_1_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_1_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_1_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_1_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_1_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_1_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_1_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_1_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_1_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_1_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_1_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_1_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_1_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_1_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_1_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_1_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_1_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_1_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_1_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_1_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_1_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_1_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_1_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_1_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_1_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_1_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_1_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_1_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_1_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_1_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_1_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_1_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_1_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_1_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_1_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_1_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_1_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_1_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_1_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_1_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_1_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_1_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_1_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_1_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_1_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_1_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_1_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_1_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_1_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_1_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_1_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_1_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_1_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_1_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_1_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_1_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_1_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_1_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_1_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_1_io_dram_rresp_ready),
    .io_dram_rresp_valid(dramArbs_1_io_dram_rresp_valid),
    .io_dram_rresp_bits_rdata_0(dramArbs_1_io_dram_rresp_bits_rdata_0),
    .io_dram_rresp_bits_rdata_1(dramArbs_1_io_dram_rresp_bits_rdata_1),
    .io_dram_rresp_bits_rdata_2(dramArbs_1_io_dram_rresp_bits_rdata_2),
    .io_dram_rresp_bits_rdata_3(dramArbs_1_io_dram_rresp_bits_rdata_3),
    .io_dram_rresp_bits_rdata_4(dramArbs_1_io_dram_rresp_bits_rdata_4),
    .io_dram_rresp_bits_rdata_5(dramArbs_1_io_dram_rresp_bits_rdata_5),
    .io_dram_rresp_bits_rdata_6(dramArbs_1_io_dram_rresp_bits_rdata_6),
    .io_dram_rresp_bits_rdata_7(dramArbs_1_io_dram_rresp_bits_rdata_7),
    .io_dram_rresp_bits_tag(dramArbs_1_io_dram_rresp_bits_tag),
    .io_dram_wresp_ready(dramArbs_1_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_1_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_1_io_dram_wresp_bits_tag),
    .io_debugSignals_0(dramArbs_1_io_debugSignals_0),
    .io_debugSignals_1(dramArbs_1_io_debugSignals_1),
    .io_debugSignals_2(dramArbs_1_io_debugSignals_2),
    .io_debugSignals_3(dramArbs_1_io_debugSignals_3),
    .io_debugSignals_4(dramArbs_1_io_debugSignals_4),
    .io_debugSignals_5(dramArbs_1_io_debugSignals_5),
    .io_debugSignals_6(dramArbs_1_io_debugSignals_6),
    .io_debugSignals_7(dramArbs_1_io_debugSignals_7),
    .io_debugSignals_8(dramArbs_1_io_debugSignals_8),
    .io_debugSignals_9(dramArbs_1_io_debugSignals_9),
    .io_debugSignals_10(dramArbs_1_io_debugSignals_10),
    .io_debugSignals_11(dramArbs_1_io_debugSignals_11),
    .io_debugSignals_12(dramArbs_1_io_debugSignals_12),
    .io_debugSignals_13(dramArbs_1_io_debugSignals_13),
    .io_debugSignals_14(dramArbs_1_io_debugSignals_14),
    .io_debugSignals_15(dramArbs_1_io_debugSignals_15),
    .io_debugSignals_16(dramArbs_1_io_debugSignals_16),
    .io_debugSignals_17(dramArbs_1_io_debugSignals_17),
    .io_debugSignals_18(dramArbs_1_io_debugSignals_18),
    .io_debugSignals_19(dramArbs_1_io_debugSignals_19),
    .io_debugSignals_20(dramArbs_1_io_debugSignals_20),
    .io_debugSignals_21(dramArbs_1_io_debugSignals_21),
    .io_debugSignals_22(dramArbs_1_io_debugSignals_22),
    .io_debugSignals_23(dramArbs_1_io_debugSignals_23),
    .io_debugSignals_24(dramArbs_1_io_debugSignals_24),
    .io_debugSignals_25(dramArbs_1_io_debugSignals_25),
    .io_debugSignals_26(dramArbs_1_io_debugSignals_26),
    .io_debugSignals_27(dramArbs_1_io_debugSignals_27),
    .io_debugSignals_28(dramArbs_1_io_debugSignals_28),
    .io_debugSignals_29(dramArbs_1_io_debugSignals_29),
    .io_debugSignals_30(dramArbs_1_io_debugSignals_30),
    .io_debugSignals_41(dramArbs_1_io_debugSignals_41)
  );
  DRAMHeap heap ( // @[Fringe.scala 107:20:@161465.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@161474.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argIns_3(regs_io_argIns_3),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits),
    .io_argOuts_2_bits(regs_io_argOuts_2_bits),
    .io_argOuts_3_bits(regs_io_argOuts_3_bits),
    .io_argOuts_4_bits(regs_io_argOuts_4_bits),
    .io_argOuts_5_bits(regs_io_argOuts_5_bits),
    .io_argOuts_6_bits(regs_io_argOuts_6_bits),
    .io_argOuts_7_bits(regs_io_argOuts_7_bits),
    .io_argOuts_8_bits(regs_io_argOuts_8_bits),
    .io_argOuts_9_bits(regs_io_argOuts_9_bits),
    .io_argOuts_10_bits(regs_io_argOuts_10_bits),
    .io_argOuts_11_bits(regs_io_argOuts_11_bits),
    .io_argOuts_12_bits(regs_io_argOuts_12_bits),
    .io_argOuts_13_bits(regs_io_argOuts_13_bits),
    .io_argOuts_14_bits(regs_io_argOuts_14_bits),
    .io_argOuts_15_bits(regs_io_argOuts_15_bits),
    .io_argOuts_16_bits(regs_io_argOuts_16_bits),
    .io_argOuts_17_bits(regs_io_argOuts_17_bits),
    .io_argOuts_18_bits(regs_io_argOuts_18_bits),
    .io_argOuts_19_bits(regs_io_argOuts_19_bits),
    .io_argOuts_20_bits(regs_io_argOuts_20_bits),
    .io_argOuts_21_bits(regs_io_argOuts_21_bits),
    .io_argOuts_22_bits(regs_io_argOuts_22_bits),
    .io_argOuts_23_bits(regs_io_argOuts_23_bits),
    .io_argOuts_24_bits(regs_io_argOuts_24_bits),
    .io_argOuts_25_bits(regs_io_argOuts_25_bits),
    .io_argOuts_26_bits(regs_io_argOuts_26_bits),
    .io_argOuts_27_bits(regs_io_argOuts_27_bits),
    .io_argOuts_28_bits(regs_io_argOuts_28_bits),
    .io_argOuts_29_bits(regs_io_argOuts_29_bits),
    .io_argOuts_30_bits(regs_io_argOuts_30_bits),
    .io_argOuts_31_bits(regs_io_argOuts_31_bits),
    .io_argOuts_32_bits(regs_io_argOuts_32_bits),
    .io_argOuts_43_bits(regs_io_argOuts_43_bits),
    .io_argEchos_1(regs_io_argEchos_1)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@163524.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@163543.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_548 = regs_io_argIns_1; // @[:@163501.4 :@163502.4]
  assign curStatus_done = _T_548[0]; // @[Fringe.scala 133:45:@163503.4]
  assign curStatus_timeout = _T_548[1]; // @[Fringe.scala 133:45:@163505.4]
  assign curStatus_allocDealloc = _T_548[4:2]; // @[Fringe.scala 133:45:@163507.4]
  assign curStatus_sizeAddr = _T_548[63:5]; // @[Fringe.scala 133:45:@163509.4]
  assign _T_553 = regs_io_argIns_0[0]; // @[Fringe.scala 134:60:@163511.4]
  assign _T_557 = curStatus_done == 1'h0; // @[Fringe.scala 134:74:@163513.4]
  assign _T_558 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@163515.4]
  assign _T_568 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@163551.4]
  assign _T_576 = _T_575 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@163556.4]
  assign _T_577 = heap_io_host_0_req_valid & _T_576; // @[package.scala 153:8:@163557.4]
  assign _T_580 = _T_553 & depulser_io_out; // @[Fringe.scala 160:55:@163561.4]
  assign status_bits_done = depulser_io_out ? _T_580 : curStatus_done; // @[Fringe.scala 160:26:@163562.4]
  assign _T_583 = _T_553 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@163565.4]
  assign status_bits_timeout = depulser_io_out ? _T_583 : curStatus_timeout; // @[Fringe.scala 161:29:@163566.4]
  assign _T_587 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@163568.4]
  assign _T_589 = heap_io_host_0_req_valid ? _T_587 : 2'h0; // @[Fringe.scala 162:34:@163569.4]
  assign _T_591 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@163571.4]
  assign _T_592 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@163574.4]
  assign status_bits_sizeAddr = _T_591[58:0]; // @[Fringe.scala 158:20:@163553.4 Fringe.scala 163:24:@163572.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_589}; // @[Fringe.scala 158:20:@163553.4 Fringe.scala 162:28:@163570.4]
  assign _T_593 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@163575.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@164779.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@164780.4]
  assign _T_1097 = alloc | dealloc; // @[Fringe.scala 204:37:@164781.4]
  assign _T_1101 = _T_1100 ^ _T_1097; // @[package.scala 153:13:@164784.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@163499.4]
  assign io_enable = _T_553 & _T_557; // @[Fringe.scala 136:13:@163519.4]
  assign io_reset = _T_558 | reset; // @[Fringe.scala 137:12:@163520.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@163541.4]
  assign io_argIns_1 = regs_io_argIns_3; // @[Fringe.scala 151:51:@163542.4]
  assign io_argEchos_0 = regs_io_argEchos_1; // @[Fringe.scala 174:24:@163578.4]
  assign io_memStreams_loads_0_cmd_ready = dramArbs_0_io_app_loads_0_cmd_ready; // @[Fringe.scala 100:70:@160547.4]
  assign io_memStreams_loads_0_data_valid = dramArbs_0_io_app_loads_0_data_valid; // @[Fringe.scala 100:70:@160542.4]
  assign io_memStreams_loads_0_data_bits_rdata_0 = dramArbs_0_io_app_loads_0_data_bits_rdata_0; // @[Fringe.scala 100:70:@160541.4]
  assign io_memStreams_stores_0_cmd_ready = dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 101:72:@160558.4]
  assign io_memStreams_stores_0_data_ready = dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 101:72:@160554.4]
  assign io_memStreams_stores_0_wresp_valid = dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 101:72:@160549.4]
  assign io_memStreams_stores_0_wresp_bits = dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 101:72:@160548.4]
  assign io_dram_0_cmd_valid = dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 195:72:@164681.4]
  assign io_dram_0_cmd_bits_addr = dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@164680.4]
  assign io_dram_0_cmd_bits_size = dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@164679.4]
  assign io_dram_0_cmd_bits_isWr = dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@164677.4]
  assign io_dram_0_cmd_bits_tag = dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@164676.4]
  assign io_dram_0_wdata_valid = dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 195:72:@164674.4]
  assign io_dram_0_wdata_bits_wdata_0 = dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@164666.4]
  assign io_dram_0_wdata_bits_wdata_1 = dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@164667.4]
  assign io_dram_0_wdata_bits_wdata_2 = dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@164668.4]
  assign io_dram_0_wdata_bits_wdata_3 = dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@164669.4]
  assign io_dram_0_wdata_bits_wdata_4 = dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@164670.4]
  assign io_dram_0_wdata_bits_wdata_5 = dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@164671.4]
  assign io_dram_0_wdata_bits_wdata_6 = dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@164672.4]
  assign io_dram_0_wdata_bits_wdata_7 = dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@164673.4]
  assign io_dram_0_wdata_bits_wstrb_0 = dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@164602.4]
  assign io_dram_0_wdata_bits_wstrb_1 = dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@164603.4]
  assign io_dram_0_wdata_bits_wstrb_2 = dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@164604.4]
  assign io_dram_0_wdata_bits_wstrb_3 = dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@164605.4]
  assign io_dram_0_wdata_bits_wstrb_4 = dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@164606.4]
  assign io_dram_0_wdata_bits_wstrb_5 = dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@164607.4]
  assign io_dram_0_wdata_bits_wstrb_6 = dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@164608.4]
  assign io_dram_0_wdata_bits_wstrb_7 = dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@164609.4]
  assign io_dram_0_wdata_bits_wstrb_8 = dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@164610.4]
  assign io_dram_0_wdata_bits_wstrb_9 = dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@164611.4]
  assign io_dram_0_wdata_bits_wstrb_10 = dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@164612.4]
  assign io_dram_0_wdata_bits_wstrb_11 = dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@164613.4]
  assign io_dram_0_wdata_bits_wstrb_12 = dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@164614.4]
  assign io_dram_0_wdata_bits_wstrb_13 = dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@164615.4]
  assign io_dram_0_wdata_bits_wstrb_14 = dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@164616.4]
  assign io_dram_0_wdata_bits_wstrb_15 = dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@164617.4]
  assign io_dram_0_wdata_bits_wstrb_16 = dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@164618.4]
  assign io_dram_0_wdata_bits_wstrb_17 = dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@164619.4]
  assign io_dram_0_wdata_bits_wstrb_18 = dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@164620.4]
  assign io_dram_0_wdata_bits_wstrb_19 = dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@164621.4]
  assign io_dram_0_wdata_bits_wstrb_20 = dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@164622.4]
  assign io_dram_0_wdata_bits_wstrb_21 = dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@164623.4]
  assign io_dram_0_wdata_bits_wstrb_22 = dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@164624.4]
  assign io_dram_0_wdata_bits_wstrb_23 = dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@164625.4]
  assign io_dram_0_wdata_bits_wstrb_24 = dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@164626.4]
  assign io_dram_0_wdata_bits_wstrb_25 = dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@164627.4]
  assign io_dram_0_wdata_bits_wstrb_26 = dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@164628.4]
  assign io_dram_0_wdata_bits_wstrb_27 = dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@164629.4]
  assign io_dram_0_wdata_bits_wstrb_28 = dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@164630.4]
  assign io_dram_0_wdata_bits_wstrb_29 = dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@164631.4]
  assign io_dram_0_wdata_bits_wstrb_30 = dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@164632.4]
  assign io_dram_0_wdata_bits_wstrb_31 = dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@164633.4]
  assign io_dram_0_wdata_bits_wstrb_32 = dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@164634.4]
  assign io_dram_0_wdata_bits_wstrb_33 = dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@164635.4]
  assign io_dram_0_wdata_bits_wstrb_34 = dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@164636.4]
  assign io_dram_0_wdata_bits_wstrb_35 = dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@164637.4]
  assign io_dram_0_wdata_bits_wstrb_36 = dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@164638.4]
  assign io_dram_0_wdata_bits_wstrb_37 = dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@164639.4]
  assign io_dram_0_wdata_bits_wstrb_38 = dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@164640.4]
  assign io_dram_0_wdata_bits_wstrb_39 = dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@164641.4]
  assign io_dram_0_wdata_bits_wstrb_40 = dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@164642.4]
  assign io_dram_0_wdata_bits_wstrb_41 = dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@164643.4]
  assign io_dram_0_wdata_bits_wstrb_42 = dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@164644.4]
  assign io_dram_0_wdata_bits_wstrb_43 = dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@164645.4]
  assign io_dram_0_wdata_bits_wstrb_44 = dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@164646.4]
  assign io_dram_0_wdata_bits_wstrb_45 = dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@164647.4]
  assign io_dram_0_wdata_bits_wstrb_46 = dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@164648.4]
  assign io_dram_0_wdata_bits_wstrb_47 = dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@164649.4]
  assign io_dram_0_wdata_bits_wstrb_48 = dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@164650.4]
  assign io_dram_0_wdata_bits_wstrb_49 = dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@164651.4]
  assign io_dram_0_wdata_bits_wstrb_50 = dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@164652.4]
  assign io_dram_0_wdata_bits_wstrb_51 = dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@164653.4]
  assign io_dram_0_wdata_bits_wstrb_52 = dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@164654.4]
  assign io_dram_0_wdata_bits_wstrb_53 = dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@164655.4]
  assign io_dram_0_wdata_bits_wstrb_54 = dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@164656.4]
  assign io_dram_0_wdata_bits_wstrb_55 = dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@164657.4]
  assign io_dram_0_wdata_bits_wstrb_56 = dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@164658.4]
  assign io_dram_0_wdata_bits_wstrb_57 = dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@164659.4]
  assign io_dram_0_wdata_bits_wstrb_58 = dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@164660.4]
  assign io_dram_0_wdata_bits_wstrb_59 = dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@164661.4]
  assign io_dram_0_wdata_bits_wstrb_60 = dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@164662.4]
  assign io_dram_0_wdata_bits_wstrb_61 = dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@164663.4]
  assign io_dram_0_wdata_bits_wstrb_62 = dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@164664.4]
  assign io_dram_0_wdata_bits_wstrb_63 = dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@164665.4]
  assign io_dram_0_wdata_bits_wlast = dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@164601.4]
  assign io_dram_0_rresp_ready = dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 195:72:@164600.4]
  assign io_dram_0_wresp_ready = dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 195:72:@164589.4]
  assign io_dram_1_cmd_valid = dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 195:72:@164777.4]
  assign io_dram_1_cmd_bits_addr = dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@164776.4]
  assign io_dram_1_cmd_bits_size = dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@164775.4]
  assign io_dram_1_cmd_bits_isWr = dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@164773.4]
  assign io_dram_1_cmd_bits_tag = dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@164772.4]
  assign io_dram_1_wdata_valid = dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 195:72:@164770.4]
  assign io_dram_1_wdata_bits_wdata_0 = dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@164762.4]
  assign io_dram_1_wdata_bits_wdata_1 = dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@164763.4]
  assign io_dram_1_wdata_bits_wdata_2 = dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@164764.4]
  assign io_dram_1_wdata_bits_wdata_3 = dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@164765.4]
  assign io_dram_1_wdata_bits_wdata_4 = dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@164766.4]
  assign io_dram_1_wdata_bits_wdata_5 = dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@164767.4]
  assign io_dram_1_wdata_bits_wdata_6 = dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@164768.4]
  assign io_dram_1_wdata_bits_wdata_7 = dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@164769.4]
  assign io_dram_1_wdata_bits_wstrb_0 = dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@164698.4]
  assign io_dram_1_wdata_bits_wstrb_1 = dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@164699.4]
  assign io_dram_1_wdata_bits_wstrb_2 = dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@164700.4]
  assign io_dram_1_wdata_bits_wstrb_3 = dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@164701.4]
  assign io_dram_1_wdata_bits_wstrb_4 = dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@164702.4]
  assign io_dram_1_wdata_bits_wstrb_5 = dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@164703.4]
  assign io_dram_1_wdata_bits_wstrb_6 = dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@164704.4]
  assign io_dram_1_wdata_bits_wstrb_7 = dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@164705.4]
  assign io_dram_1_wdata_bits_wstrb_8 = dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@164706.4]
  assign io_dram_1_wdata_bits_wstrb_9 = dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@164707.4]
  assign io_dram_1_wdata_bits_wstrb_10 = dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@164708.4]
  assign io_dram_1_wdata_bits_wstrb_11 = dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@164709.4]
  assign io_dram_1_wdata_bits_wstrb_12 = dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@164710.4]
  assign io_dram_1_wdata_bits_wstrb_13 = dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@164711.4]
  assign io_dram_1_wdata_bits_wstrb_14 = dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@164712.4]
  assign io_dram_1_wdata_bits_wstrb_15 = dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@164713.4]
  assign io_dram_1_wdata_bits_wstrb_16 = dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@164714.4]
  assign io_dram_1_wdata_bits_wstrb_17 = dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@164715.4]
  assign io_dram_1_wdata_bits_wstrb_18 = dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@164716.4]
  assign io_dram_1_wdata_bits_wstrb_19 = dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@164717.4]
  assign io_dram_1_wdata_bits_wstrb_20 = dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@164718.4]
  assign io_dram_1_wdata_bits_wstrb_21 = dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@164719.4]
  assign io_dram_1_wdata_bits_wstrb_22 = dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@164720.4]
  assign io_dram_1_wdata_bits_wstrb_23 = dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@164721.4]
  assign io_dram_1_wdata_bits_wstrb_24 = dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@164722.4]
  assign io_dram_1_wdata_bits_wstrb_25 = dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@164723.4]
  assign io_dram_1_wdata_bits_wstrb_26 = dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@164724.4]
  assign io_dram_1_wdata_bits_wstrb_27 = dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@164725.4]
  assign io_dram_1_wdata_bits_wstrb_28 = dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@164726.4]
  assign io_dram_1_wdata_bits_wstrb_29 = dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@164727.4]
  assign io_dram_1_wdata_bits_wstrb_30 = dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@164728.4]
  assign io_dram_1_wdata_bits_wstrb_31 = dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@164729.4]
  assign io_dram_1_wdata_bits_wstrb_32 = dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@164730.4]
  assign io_dram_1_wdata_bits_wstrb_33 = dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@164731.4]
  assign io_dram_1_wdata_bits_wstrb_34 = dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@164732.4]
  assign io_dram_1_wdata_bits_wstrb_35 = dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@164733.4]
  assign io_dram_1_wdata_bits_wstrb_36 = dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@164734.4]
  assign io_dram_1_wdata_bits_wstrb_37 = dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@164735.4]
  assign io_dram_1_wdata_bits_wstrb_38 = dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@164736.4]
  assign io_dram_1_wdata_bits_wstrb_39 = dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@164737.4]
  assign io_dram_1_wdata_bits_wstrb_40 = dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@164738.4]
  assign io_dram_1_wdata_bits_wstrb_41 = dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@164739.4]
  assign io_dram_1_wdata_bits_wstrb_42 = dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@164740.4]
  assign io_dram_1_wdata_bits_wstrb_43 = dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@164741.4]
  assign io_dram_1_wdata_bits_wstrb_44 = dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@164742.4]
  assign io_dram_1_wdata_bits_wstrb_45 = dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@164743.4]
  assign io_dram_1_wdata_bits_wstrb_46 = dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@164744.4]
  assign io_dram_1_wdata_bits_wstrb_47 = dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@164745.4]
  assign io_dram_1_wdata_bits_wstrb_48 = dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@164746.4]
  assign io_dram_1_wdata_bits_wstrb_49 = dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@164747.4]
  assign io_dram_1_wdata_bits_wstrb_50 = dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@164748.4]
  assign io_dram_1_wdata_bits_wstrb_51 = dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@164749.4]
  assign io_dram_1_wdata_bits_wstrb_52 = dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@164750.4]
  assign io_dram_1_wdata_bits_wstrb_53 = dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@164751.4]
  assign io_dram_1_wdata_bits_wstrb_54 = dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@164752.4]
  assign io_dram_1_wdata_bits_wstrb_55 = dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@164753.4]
  assign io_dram_1_wdata_bits_wstrb_56 = dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@164754.4]
  assign io_dram_1_wdata_bits_wstrb_57 = dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@164755.4]
  assign io_dram_1_wdata_bits_wstrb_58 = dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@164756.4]
  assign io_dram_1_wdata_bits_wstrb_59 = dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@164757.4]
  assign io_dram_1_wdata_bits_wstrb_60 = dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@164758.4]
  assign io_dram_1_wdata_bits_wstrb_61 = dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@164759.4]
  assign io_dram_1_wdata_bits_wstrb_62 = dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@164760.4]
  assign io_dram_1_wdata_bits_wstrb_63 = dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@164761.4]
  assign io_dram_1_wdata_bits_wlast = dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@164697.4]
  assign io_dram_1_rresp_ready = dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 195:72:@164696.4]
  assign io_dram_1_wresp_ready = dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 195:72:@164685.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@161470.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@161469.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@161468.4]
  assign dramArbs_0_clock = clock; // @[:@159718.4]
  assign dramArbs_0_reset = _T_558 | reset; // @[:@159719.4 Fringe.scala 187:30:@164583.4]
  assign dramArbs_0_io_enable = _T_553 & _T_557; // @[Fringe.scala 192:36:@164585.4]
  assign dramArbs_0_io_app_loads_0_cmd_valid = io_memStreams_loads_0_cmd_valid; // @[Fringe.scala 100:70:@160546.4]
  assign dramArbs_0_io_app_loads_0_cmd_bits_addr = io_memStreams_loads_0_cmd_bits_addr; // @[Fringe.scala 100:70:@160545.4]
  assign dramArbs_0_io_app_loads_0_cmd_bits_size = io_memStreams_loads_0_cmd_bits_size; // @[Fringe.scala 100:70:@160544.4]
  assign dramArbs_0_io_app_loads_0_data_ready = io_memStreams_loads_0_data_ready; // @[Fringe.scala 100:70:@160543.4]
  assign dramArbs_0_io_app_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[Fringe.scala 101:72:@160557.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[Fringe.scala 101:72:@160556.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[Fringe.scala 101:72:@160555.4]
  assign dramArbs_0_io_app_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[Fringe.scala 101:72:@160553.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[Fringe.scala 101:72:@160552.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[Fringe.scala 101:72:@160551.4]
  assign dramArbs_0_io_app_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[Fringe.scala 101:72:@160550.4]
  assign dramArbs_0_io_dram_cmd_ready = io_dram_0_cmd_ready; // @[Fringe.scala 195:72:@164682.4]
  assign dramArbs_0_io_dram_wdata_ready = io_dram_0_wdata_ready; // @[Fringe.scala 195:72:@164675.4]
  assign dramArbs_0_io_dram_rresp_valid = io_dram_0_rresp_valid; // @[Fringe.scala 195:72:@164599.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_0 = io_dram_0_rresp_bits_rdata_0; // @[Fringe.scala 195:72:@164591.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_1 = io_dram_0_rresp_bits_rdata_1; // @[Fringe.scala 195:72:@164592.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_2 = io_dram_0_rresp_bits_rdata_2; // @[Fringe.scala 195:72:@164593.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_3 = io_dram_0_rresp_bits_rdata_3; // @[Fringe.scala 195:72:@164594.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_4 = io_dram_0_rresp_bits_rdata_4; // @[Fringe.scala 195:72:@164595.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_5 = io_dram_0_rresp_bits_rdata_5; // @[Fringe.scala 195:72:@164596.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_6 = io_dram_0_rresp_bits_rdata_6; // @[Fringe.scala 195:72:@164597.4]
  assign dramArbs_0_io_dram_rresp_bits_rdata_7 = io_dram_0_rresp_bits_rdata_7; // @[Fringe.scala 195:72:@164598.4]
  assign dramArbs_0_io_dram_rresp_bits_tag = io_dram_0_rresp_bits_tag; // @[Fringe.scala 195:72:@164590.4]
  assign dramArbs_0_io_dram_wresp_valid = io_dram_0_wresp_valid; // @[Fringe.scala 195:72:@164588.4]
  assign dramArbs_0_io_dram_wresp_bits_tag = io_dram_0_wresp_bits_tag; // @[Fringe.scala 195:72:@164587.4]
  assign dramArbs_1_clock = clock; // @[:@160601.4]
  assign dramArbs_1_reset = _T_558 | reset; // @[:@160602.4 Fringe.scala 187:30:@164584.4]
  assign dramArbs_1_io_enable = _T_553 & _T_557; // @[Fringe.scala 192:36:@164586.4]
  assign dramArbs_1_io_app_loads_0_cmd_valid = 1'h0;
  assign dramArbs_1_io_app_loads_0_cmd_bits_addr = 64'h0;
  assign dramArbs_1_io_app_loads_0_cmd_bits_size = 32'h0;
  assign dramArbs_1_io_app_loads_0_data_ready = 1'h0;
  assign dramArbs_1_io_app_stores_0_cmd_valid = 1'h0;
  assign dramArbs_1_io_app_stores_0_cmd_bits_addr = 64'h0;
  assign dramArbs_1_io_app_stores_0_cmd_bits_size = 32'h0;
  assign dramArbs_1_io_app_stores_0_data_valid = 1'h0;
  assign dramArbs_1_io_app_stores_0_data_bits_wdata_0 = 32'h0;
  assign dramArbs_1_io_app_stores_0_data_bits_wstrb = 1'h0;
  assign dramArbs_1_io_app_stores_0_wresp_ready = 1'h0;
  assign dramArbs_1_io_dram_cmd_ready = io_dram_1_cmd_ready; // @[Fringe.scala 195:72:@164778.4]
  assign dramArbs_1_io_dram_wdata_ready = io_dram_1_wdata_ready; // @[Fringe.scala 195:72:@164771.4]
  assign dramArbs_1_io_dram_rresp_valid = io_dram_1_rresp_valid; // @[Fringe.scala 195:72:@164695.4]
  assign dramArbs_1_io_dram_rresp_bits_rdata_0 = io_dram_1_rresp_bits_rdata_0; // @[Fringe.scala 195:72:@164687.4]
  assign dramArbs_1_io_dram_rresp_bits_rdata_1 = io_dram_1_rresp_bits_rdata_1; // @[Fringe.scala 195:72:@164688.4]
  assign dramArbs_1_io_dram_rresp_bits_rdata_2 = io_dram_1_rresp_bits_rdata_2; // @[Fringe.scala 195:72:@164689.4]
  assign dramArbs_1_io_dram_rresp_bits_rdata_3 = io_dram_1_rresp_bits_rdata_3; // @[Fringe.scala 195:72:@164690.4]
  assign dramArbs_1_io_dram_rresp_bits_rdata_4 = io_dram_1_rresp_bits_rdata_4; // @[Fringe.scala 195:72:@164691.4]
  assign dramArbs_1_io_dram_rresp_bits_rdata_5 = io_dram_1_rresp_bits_rdata_5; // @[Fringe.scala 195:72:@164692.4]
  assign dramArbs_1_io_dram_rresp_bits_rdata_6 = io_dram_1_rresp_bits_rdata_6; // @[Fringe.scala 195:72:@164693.4]
  assign dramArbs_1_io_dram_rresp_bits_rdata_7 = io_dram_1_rresp_bits_rdata_7; // @[Fringe.scala 195:72:@164694.4]
  assign dramArbs_1_io_dram_rresp_bits_tag = io_dram_1_rresp_bits_tag; // @[Fringe.scala 195:72:@164686.4]
  assign dramArbs_1_io_dram_wresp_valid = io_dram_1_wresp_valid; // @[Fringe.scala 195:72:@164684.4]
  assign dramArbs_1_io_dram_wresp_bits_tag = io_dram_1_wresp_bits_tag; // @[Fringe.scala 195:72:@164683.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@161473.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@161472.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@161471.4]
  assign heap_io_host_0_resp_valid = _T_1097 & _T_1101; // @[Fringe.scala 204:22:@164786.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@164787.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@164788.4]
  assign regs_clock = clock; // @[:@161475.4]
  assign regs_reset = reset; // @[:@161476.4 Fringe.scala 139:14:@163523.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@163495.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@163497.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@163496.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@163498.4]
  assign regs_io_reset = _T_558 | reset; // @[Fringe.scala 138:17:@163521.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_577; // @[Fringe.scala 170:23:@163573.4]
  assign regs_io_argOuts_0_bits = {_T_593,_T_592}; // @[Fringe.scala 171:22:@163577.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@163580.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@163579.4]
  assign regs_io_argOuts_2_bits = {{32'd0}, dramArbs_0_io_debugSignals_0}; // @[Fringe.scala 179:22:@163581.4]
  assign regs_io_argOuts_3_bits = {{32'd0}, dramArbs_0_io_debugSignals_1}; // @[Fringe.scala 179:22:@163583.4]
  assign regs_io_argOuts_4_bits = {{32'd0}, dramArbs_0_io_debugSignals_2}; // @[Fringe.scala 179:22:@163585.4]
  assign regs_io_argOuts_5_bits = {{32'd0}, dramArbs_0_io_debugSignals_3}; // @[Fringe.scala 179:22:@163587.4]
  assign regs_io_argOuts_6_bits = {{32'd0}, dramArbs_0_io_debugSignals_4}; // @[Fringe.scala 179:22:@163589.4]
  assign regs_io_argOuts_7_bits = {{32'd0}, dramArbs_0_io_debugSignals_5}; // @[Fringe.scala 179:22:@163591.4]
  assign regs_io_argOuts_8_bits = {{32'd0}, dramArbs_0_io_debugSignals_6}; // @[Fringe.scala 179:22:@163593.4]
  assign regs_io_argOuts_9_bits = {{32'd0}, dramArbs_0_io_debugSignals_7}; // @[Fringe.scala 179:22:@163595.4]
  assign regs_io_argOuts_10_bits = {{32'd0}, dramArbs_0_io_debugSignals_8}; // @[Fringe.scala 179:22:@163597.4]
  assign regs_io_argOuts_11_bits = {{32'd0}, dramArbs_0_io_debugSignals_9}; // @[Fringe.scala 179:22:@163599.4]
  assign regs_io_argOuts_12_bits = {{32'd0}, dramArbs_0_io_debugSignals_10}; // @[Fringe.scala 179:22:@163601.4]
  assign regs_io_argOuts_13_bits = {{32'd0}, dramArbs_0_io_debugSignals_11}; // @[Fringe.scala 179:22:@163603.4]
  assign regs_io_argOuts_14_bits = {{32'd0}, dramArbs_0_io_debugSignals_12}; // @[Fringe.scala 179:22:@163605.4]
  assign regs_io_argOuts_15_bits = {{32'd0}, dramArbs_0_io_debugSignals_13}; // @[Fringe.scala 179:22:@163607.4]
  assign regs_io_argOuts_16_bits = {{32'd0}, dramArbs_0_io_debugSignals_14}; // @[Fringe.scala 179:22:@163609.4]
  assign regs_io_argOuts_17_bits = {{32'd0}, dramArbs_0_io_debugSignals_15}; // @[Fringe.scala 179:22:@163611.4]
  assign regs_io_argOuts_18_bits = {{32'd0}, dramArbs_0_io_debugSignals_16}; // @[Fringe.scala 179:22:@163613.4]
  assign regs_io_argOuts_19_bits = {{32'd0}, dramArbs_0_io_debugSignals_17}; // @[Fringe.scala 179:22:@163615.4]
  assign regs_io_argOuts_20_bits = {{32'd0}, dramArbs_0_io_debugSignals_18}; // @[Fringe.scala 179:22:@163617.4]
  assign regs_io_argOuts_21_bits = {{32'd0}, dramArbs_0_io_debugSignals_19}; // @[Fringe.scala 179:22:@163619.4]
  assign regs_io_argOuts_22_bits = {{32'd0}, dramArbs_0_io_debugSignals_20}; // @[Fringe.scala 179:22:@163621.4]
  assign regs_io_argOuts_23_bits = {{32'd0}, dramArbs_0_io_debugSignals_21}; // @[Fringe.scala 179:22:@163623.4]
  assign regs_io_argOuts_24_bits = {{32'd0}, dramArbs_0_io_debugSignals_22}; // @[Fringe.scala 179:22:@163625.4]
  assign regs_io_argOuts_25_bits = {{32'd0}, dramArbs_0_io_debugSignals_23}; // @[Fringe.scala 179:22:@163627.4]
  assign regs_io_argOuts_26_bits = {{32'd0}, dramArbs_0_io_debugSignals_24}; // @[Fringe.scala 179:22:@163629.4]
  assign regs_io_argOuts_27_bits = {{32'd0}, dramArbs_0_io_debugSignals_25}; // @[Fringe.scala 179:22:@163631.4]
  assign regs_io_argOuts_28_bits = {{32'd0}, dramArbs_0_io_debugSignals_26}; // @[Fringe.scala 179:22:@163633.4]
  assign regs_io_argOuts_29_bits = {{32'd0}, dramArbs_0_io_debugSignals_27}; // @[Fringe.scala 179:22:@163635.4]
  assign regs_io_argOuts_30_bits = {{32'd0}, dramArbs_0_io_debugSignals_28}; // @[Fringe.scala 179:22:@163637.4]
  assign regs_io_argOuts_31_bits = {{32'd0}, dramArbs_0_io_debugSignals_29}; // @[Fringe.scala 179:22:@163639.4]
  assign regs_io_argOuts_32_bits = {{32'd0}, dramArbs_0_io_debugSignals_30}; // @[Fringe.scala 179:22:@163641.4]
  assign regs_io_argOuts_43_bits = {{32'd0}, dramArbs_0_io_debugSignals_41}; // @[Fringe.scala 179:22:@163663.4]
  assign timeoutCtr_clock = clock; // @[:@163525.4]
  assign timeoutCtr_reset = reset; // @[:@163526.4]
  assign timeoutCtr_io_enable = _T_553 & _T_557; // @[Fringe.scala 149:24:@163540.4]
  assign depulser_clock = clock; // @[:@163544.4]
  assign depulser_reset = reset; // @[:@163545.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@163550.4]
  assign depulser_io_rst = _T_568[0]; // @[Fringe.scala 156:19:@163552.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_575 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1100 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_575 <= 1'h0;
    end else begin
      _T_575 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1100 <= 1'h0;
    end else begin
      _T_1100 <= _T_1097;
    end
  end
endmodule
module AXI4LiteToRFBridgeZCU( // @[:@164803.2]
  input         clock, // @[:@164804.4]
  input         reset, // @[:@164805.4]
  input  [39:0] io_S_AXI_AWADDR, // @[:@164806.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@164806.4]
  input         io_S_AXI_AWVALID, // @[:@164806.4]
  output        io_S_AXI_AWREADY, // @[:@164806.4]
  input  [39:0] io_S_AXI_ARADDR, // @[:@164806.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@164806.4]
  input         io_S_AXI_ARVALID, // @[:@164806.4]
  output        io_S_AXI_ARREADY, // @[:@164806.4]
  input  [63:0] io_S_AXI_WDATA, // @[:@164806.4]
  input  [7:0]  io_S_AXI_WSTRB, // @[:@164806.4]
  input         io_S_AXI_WVALID, // @[:@164806.4]
  output        io_S_AXI_WREADY, // @[:@164806.4]
  output [63:0] io_S_AXI_RDATA, // @[:@164806.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@164806.4]
  output        io_S_AXI_RVALID, // @[:@164806.4]
  input         io_S_AXI_RREADY, // @[:@164806.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@164806.4]
  output        io_S_AXI_BVALID, // @[:@164806.4]
  input         io_S_AXI_BREADY, // @[:@164806.4]
  output [39:0] io_raddr, // @[:@164806.4]
  output        io_wen, // @[:@164806.4]
  output [39:0] io_waddr, // @[:@164806.4]
  output [63:0] io_wdata, // @[:@164806.4]
  input  [63:0] io_rdata // @[:@164806.4]
);
  wire [63:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire [63:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire [39:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire [39:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire [39:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire [39:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire [63:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire [7:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire [63:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
  AXI4LiteToRFBridgeZCUVerilog d ( // @[AXI4LiteToRFBridge.scala 82:17:@164808.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 84:14:@164832.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 84:14:@164828.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 84:14:@164824.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 84:14:@164823.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 84:14:@164822.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 84:14:@164821.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 84:14:@164819.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 84:14:@164818.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 88:12:@164840.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 91:12:@164843.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 89:12:@164841.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 90:12:@164842.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 92:17:@164844.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 86:22:@164839.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 85:19:@164836.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 84:14:@164835.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 84:14:@164834.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 84:14:@164833.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 84:14:@164831.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 84:14:@164830.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 84:14:@164829.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 84:14:@164827.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 84:14:@164826.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 84:14:@164825.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 84:14:@164820.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 84:14:@164817.4]
endmodule
module MAGToAXI4Bridge( // @[:@164846.2]
  output         io_in_cmd_ready, // @[:@164849.4]
  input          io_in_cmd_valid, // @[:@164849.4]
  input  [63:0]  io_in_cmd_bits_addr, // @[:@164849.4]
  input  [31:0]  io_in_cmd_bits_size, // @[:@164849.4]
  input          io_in_cmd_bits_isWr, // @[:@164849.4]
  input  [31:0]  io_in_cmd_bits_tag, // @[:@164849.4]
  output         io_in_wdata_ready, // @[:@164849.4]
  input          io_in_wdata_valid, // @[:@164849.4]
  input  [63:0]  io_in_wdata_bits_wdata_0, // @[:@164849.4]
  input  [63:0]  io_in_wdata_bits_wdata_1, // @[:@164849.4]
  input  [63:0]  io_in_wdata_bits_wdata_2, // @[:@164849.4]
  input  [63:0]  io_in_wdata_bits_wdata_3, // @[:@164849.4]
  input  [63:0]  io_in_wdata_bits_wdata_4, // @[:@164849.4]
  input  [63:0]  io_in_wdata_bits_wdata_5, // @[:@164849.4]
  input  [63:0]  io_in_wdata_bits_wdata_6, // @[:@164849.4]
  input  [63:0]  io_in_wdata_bits_wdata_7, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_0, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_1, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_2, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_3, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_4, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_5, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_6, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_7, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_8, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_9, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_10, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_11, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_12, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_13, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_14, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_15, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_16, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_17, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_18, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_19, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_20, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_21, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_22, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_23, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_24, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_25, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_26, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_27, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_28, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_29, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_30, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_31, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_32, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_33, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_34, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_35, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_36, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_37, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_38, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_39, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_40, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_41, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_42, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_43, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_44, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_45, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_46, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_47, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_48, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_49, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_50, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_51, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_52, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_53, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_54, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_55, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_56, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_57, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_58, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_59, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_60, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_61, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_62, // @[:@164849.4]
  input          io_in_wdata_bits_wstrb_63, // @[:@164849.4]
  input          io_in_wdata_bits_wlast, // @[:@164849.4]
  input          io_in_rresp_ready, // @[:@164849.4]
  output         io_in_rresp_valid, // @[:@164849.4]
  output [63:0]  io_in_rresp_bits_rdata_0, // @[:@164849.4]
  output [63:0]  io_in_rresp_bits_rdata_1, // @[:@164849.4]
  output [63:0]  io_in_rresp_bits_rdata_2, // @[:@164849.4]
  output [63:0]  io_in_rresp_bits_rdata_3, // @[:@164849.4]
  output [63:0]  io_in_rresp_bits_rdata_4, // @[:@164849.4]
  output [63:0]  io_in_rresp_bits_rdata_5, // @[:@164849.4]
  output [63:0]  io_in_rresp_bits_rdata_6, // @[:@164849.4]
  output [63:0]  io_in_rresp_bits_rdata_7, // @[:@164849.4]
  output [31:0]  io_in_rresp_bits_tag, // @[:@164849.4]
  input          io_in_wresp_ready, // @[:@164849.4]
  output         io_in_wresp_valid, // @[:@164849.4]
  output [31:0]  io_in_wresp_bits_tag, // @[:@164849.4]
  output [31:0]  io_M_AXI_AWID, // @[:@164849.4]
  output [39:0]  io_M_AXI_AWADDR, // @[:@164849.4]
  output [7:0]   io_M_AXI_AWLEN, // @[:@164849.4]
  output         io_M_AXI_AWVALID, // @[:@164849.4]
  input          io_M_AXI_AWREADY, // @[:@164849.4]
  output [31:0]  io_M_AXI_ARID, // @[:@164849.4]
  output [39:0]  io_M_AXI_ARADDR, // @[:@164849.4]
  output [7:0]   io_M_AXI_ARLEN, // @[:@164849.4]
  output         io_M_AXI_ARVALID, // @[:@164849.4]
  input          io_M_AXI_ARREADY, // @[:@164849.4]
  output [511:0] io_M_AXI_WDATA, // @[:@164849.4]
  output [63:0]  io_M_AXI_WSTRB, // @[:@164849.4]
  output         io_M_AXI_WLAST, // @[:@164849.4]
  output         io_M_AXI_WVALID, // @[:@164849.4]
  input          io_M_AXI_WREADY, // @[:@164849.4]
  input  [31:0]  io_M_AXI_RID, // @[:@164849.4]
  input  [511:0] io_M_AXI_RDATA, // @[:@164849.4]
  input          io_M_AXI_RVALID, // @[:@164849.4]
  output         io_M_AXI_RREADY, // @[:@164849.4]
  input  [31:0]  io_M_AXI_BID, // @[:@164849.4]
  input          io_M_AXI_BVALID, // @[:@164849.4]
  output         io_M_AXI_BREADY // @[:@164849.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@164990.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@164991.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@164992.4]
  wire  _T_228; // @[MAGToAXI4Bridge.scala 35:42:@165000.4]
  wire [447:0] _T_247; // @[Cat.scala 30:58:@165024.4]
  wire [9:0] _T_257; // @[Cat.scala 30:58:@165035.4]
  wire [18:0] _T_266; // @[Cat.scala 30:58:@165044.4]
  wire [27:0] _T_275; // @[Cat.scala 30:58:@165053.4]
  wire [36:0] _T_284; // @[Cat.scala 30:58:@165062.4]
  wire [45:0] _T_293; // @[Cat.scala 30:58:@165071.4]
  wire [54:0] _T_302; // @[Cat.scala 30:58:@165080.4]
  wire [62:0] _T_310; // @[Cat.scala 30:58:@165088.4]
  assign _T_218 = io_in_cmd_bits_size - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@164990.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@164991.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@164992.4]
  assign _T_228 = io_in_cmd_bits_isWr == 1'h0; // @[MAGToAXI4Bridge.scala 35:42:@165000.4]
  assign _T_247 = {io_in_wdata_bits_wdata_7,io_in_wdata_bits_wdata_6,io_in_wdata_bits_wdata_5,io_in_wdata_bits_wdata_4,io_in_wdata_bits_wdata_3,io_in_wdata_bits_wdata_2,io_in_wdata_bits_wdata_1}; // @[Cat.scala 30:58:@165024.4]
  assign _T_257 = {io_in_wdata_bits_wstrb_63,io_in_wdata_bits_wstrb_62,io_in_wdata_bits_wstrb_61,io_in_wdata_bits_wstrb_60,io_in_wdata_bits_wstrb_59,io_in_wdata_bits_wstrb_58,io_in_wdata_bits_wstrb_57,io_in_wdata_bits_wstrb_56,io_in_wdata_bits_wstrb_55,io_in_wdata_bits_wstrb_54}; // @[Cat.scala 30:58:@165035.4]
  assign _T_266 = {_T_257,io_in_wdata_bits_wstrb_53,io_in_wdata_bits_wstrb_52,io_in_wdata_bits_wstrb_51,io_in_wdata_bits_wstrb_50,io_in_wdata_bits_wstrb_49,io_in_wdata_bits_wstrb_48,io_in_wdata_bits_wstrb_47,io_in_wdata_bits_wstrb_46,io_in_wdata_bits_wstrb_45}; // @[Cat.scala 30:58:@165044.4]
  assign _T_275 = {_T_266,io_in_wdata_bits_wstrb_44,io_in_wdata_bits_wstrb_43,io_in_wdata_bits_wstrb_42,io_in_wdata_bits_wstrb_41,io_in_wdata_bits_wstrb_40,io_in_wdata_bits_wstrb_39,io_in_wdata_bits_wstrb_38,io_in_wdata_bits_wstrb_37,io_in_wdata_bits_wstrb_36}; // @[Cat.scala 30:58:@165053.4]
  assign _T_284 = {_T_275,io_in_wdata_bits_wstrb_35,io_in_wdata_bits_wstrb_34,io_in_wdata_bits_wstrb_33,io_in_wdata_bits_wstrb_32,io_in_wdata_bits_wstrb_31,io_in_wdata_bits_wstrb_30,io_in_wdata_bits_wstrb_29,io_in_wdata_bits_wstrb_28,io_in_wdata_bits_wstrb_27}; // @[Cat.scala 30:58:@165062.4]
  assign _T_293 = {_T_284,io_in_wdata_bits_wstrb_26,io_in_wdata_bits_wstrb_25,io_in_wdata_bits_wstrb_24,io_in_wdata_bits_wstrb_23,io_in_wdata_bits_wstrb_22,io_in_wdata_bits_wstrb_21,io_in_wdata_bits_wstrb_20,io_in_wdata_bits_wstrb_19,io_in_wdata_bits_wstrb_18}; // @[Cat.scala 30:58:@165071.4]
  assign _T_302 = {_T_293,io_in_wdata_bits_wstrb_17,io_in_wdata_bits_wstrb_16,io_in_wdata_bits_wstrb_15,io_in_wdata_bits_wstrb_14,io_in_wdata_bits_wstrb_13,io_in_wdata_bits_wstrb_12,io_in_wdata_bits_wstrb_11,io_in_wdata_bits_wstrb_10,io_in_wdata_bits_wstrb_9}; // @[Cat.scala 30:58:@165080.4]
  assign _T_310 = {_T_302,io_in_wdata_bits_wstrb_8,io_in_wdata_bits_wstrb_7,io_in_wdata_bits_wstrb_6,io_in_wdata_bits_wstrb_5,io_in_wdata_bits_wstrb_4,io_in_wdata_bits_wstrb_3,io_in_wdata_bits_wstrb_2,io_in_wdata_bits_wstrb_1}; // @[Cat.scala 30:58:@165088.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? io_M_AXI_AWREADY : io_M_AXI_ARREADY; // @[MAGToAXI4Bridge.scala 36:21:@165004.4]
  assign io_in_wdata_ready = io_M_AXI_WREADY; // @[MAGToAXI4Bridge.scala 56:21:@165093.4]
  assign io_in_rresp_valid = io_M_AXI_RVALID; // @[MAGToAXI4Bridge.scala 70:21:@165121.4]
  assign io_in_rresp_bits_rdata_0 = io_M_AXI_RDATA[63:0]; // @[MAGToAXI4Bridge.scala 62:26:@165111.4]
  assign io_in_rresp_bits_rdata_1 = io_M_AXI_RDATA[127:64]; // @[MAGToAXI4Bridge.scala 62:26:@165112.4]
  assign io_in_rresp_bits_rdata_2 = io_M_AXI_RDATA[191:128]; // @[MAGToAXI4Bridge.scala 62:26:@165113.4]
  assign io_in_rresp_bits_rdata_3 = io_M_AXI_RDATA[255:192]; // @[MAGToAXI4Bridge.scala 62:26:@165114.4]
  assign io_in_rresp_bits_rdata_4 = io_M_AXI_RDATA[319:256]; // @[MAGToAXI4Bridge.scala 62:26:@165115.4]
  assign io_in_rresp_bits_rdata_5 = io_M_AXI_RDATA[383:320]; // @[MAGToAXI4Bridge.scala 62:26:@165116.4]
  assign io_in_rresp_bits_rdata_6 = io_M_AXI_RDATA[447:384]; // @[MAGToAXI4Bridge.scala 62:26:@165117.4]
  assign io_in_rresp_bits_rdata_7 = io_M_AXI_RDATA[511:448]; // @[MAGToAXI4Bridge.scala 62:26:@165118.4]
  assign io_in_rresp_bits_tag = io_M_AXI_RID; // @[MAGToAXI4Bridge.scala 73:24:@165123.4]
  assign io_in_wresp_valid = io_M_AXI_BVALID; // @[MAGToAXI4Bridge.scala 71:21:@165122.4]
  assign io_in_wresp_bits_tag = io_M_AXI_BID; // @[MAGToAXI4Bridge.scala 74:24:@165124.4]
  assign io_M_AXI_AWID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 39:21:@165005.4]
  assign io_M_AXI_AWADDR = io_in_cmd_bits_addr[39:0]; // @[MAGToAXI4Bridge.scala 40:21:@165006.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@165010.4]
  assign io_M_AXI_AWVALID = io_in_cmd_valid & io_in_cmd_bits_isWr; // @[MAGToAXI4Bridge.scala 49:21:@165018.4]
  assign io_M_AXI_ARID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 25:21:@164988.4]
  assign io_M_AXI_ARADDR = io_in_cmd_bits_addr[39:0]; // @[MAGToAXI4Bridge.scala 26:21:@164989.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@164993.4]
  assign io_M_AXI_ARVALID = io_in_cmd_valid & _T_228; // @[MAGToAXI4Bridge.scala 35:21:@165002.4]
  assign io_M_AXI_WDATA = {_T_247,io_in_wdata_bits_wdata_0}; // @[MAGToAXI4Bridge.scala 52:21:@165026.4]
  assign io_M_AXI_WSTRB = {_T_310,io_in_wdata_bits_wstrb_0}; // @[MAGToAXI4Bridge.scala 53:21:@165090.4]
  assign io_M_AXI_WLAST = io_in_wdata_bits_wlast; // @[MAGToAXI4Bridge.scala 54:21:@165091.4]
  assign io_M_AXI_WVALID = io_in_wdata_valid; // @[MAGToAXI4Bridge.scala 55:21:@165092.4]
  assign io_M_AXI_RREADY = io_in_rresp_ready; // @[MAGToAXI4Bridge.scala 64:19:@165119.4]
  assign io_M_AXI_BREADY = io_in_wresp_ready; // @[MAGToAXI4Bridge.scala 67:19:@165120.4]
endmodule
module FringeZynq( // @[:@165406.2]
  input          clock, // @[:@165407.4]
  input          reset, // @[:@165408.4]
  input          io_axil_s_clk, // @[:@165409.4]
  input  [39:0]  io_S_AXI_AWADDR, // @[:@165409.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@165409.4]
  input          io_S_AXI_AWVALID, // @[:@165409.4]
  output         io_S_AXI_AWREADY, // @[:@165409.4]
  input  [39:0]  io_S_AXI_ARADDR, // @[:@165409.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@165409.4]
  input          io_S_AXI_ARVALID, // @[:@165409.4]
  output         io_S_AXI_ARREADY, // @[:@165409.4]
  input  [63:0]  io_S_AXI_WDATA, // @[:@165409.4]
  input  [7:0]   io_S_AXI_WSTRB, // @[:@165409.4]
  input          io_S_AXI_WVALID, // @[:@165409.4]
  output         io_S_AXI_WREADY, // @[:@165409.4]
  output [63:0]  io_S_AXI_RDATA, // @[:@165409.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@165409.4]
  output         io_S_AXI_RVALID, // @[:@165409.4]
  input          io_S_AXI_RREADY, // @[:@165409.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@165409.4]
  output         io_S_AXI_BVALID, // @[:@165409.4]
  input          io_S_AXI_BREADY, // @[:@165409.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@165409.4]
  output [39:0]  io_M_AXI_0_AWADDR, // @[:@165409.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@165409.4]
  output         io_M_AXI_0_AWVALID, // @[:@165409.4]
  input          io_M_AXI_0_AWREADY, // @[:@165409.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@165409.4]
  output [39:0]  io_M_AXI_0_ARADDR, // @[:@165409.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@165409.4]
  output         io_M_AXI_0_ARVALID, // @[:@165409.4]
  input          io_M_AXI_0_ARREADY, // @[:@165409.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@165409.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@165409.4]
  output         io_M_AXI_0_WLAST, // @[:@165409.4]
  output         io_M_AXI_0_WVALID, // @[:@165409.4]
  input          io_M_AXI_0_WREADY, // @[:@165409.4]
  input  [31:0]  io_M_AXI_0_RID, // @[:@165409.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@165409.4]
  input          io_M_AXI_0_RVALID, // @[:@165409.4]
  output         io_M_AXI_0_RREADY, // @[:@165409.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@165409.4]
  input          io_M_AXI_0_BVALID, // @[:@165409.4]
  output         io_M_AXI_0_BREADY, // @[:@165409.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@165409.4]
  output [39:0]  io_M_AXI_1_AWADDR, // @[:@165409.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@165409.4]
  output         io_M_AXI_1_AWVALID, // @[:@165409.4]
  input          io_M_AXI_1_AWREADY, // @[:@165409.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@165409.4]
  output [39:0]  io_M_AXI_1_ARADDR, // @[:@165409.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@165409.4]
  output         io_M_AXI_1_ARVALID, // @[:@165409.4]
  input          io_M_AXI_1_ARREADY, // @[:@165409.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@165409.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@165409.4]
  output         io_M_AXI_1_WLAST, // @[:@165409.4]
  output         io_M_AXI_1_WVALID, // @[:@165409.4]
  input          io_M_AXI_1_WREADY, // @[:@165409.4]
  input  [31:0]  io_M_AXI_1_RID, // @[:@165409.4]
  input  [511:0] io_M_AXI_1_RDATA, // @[:@165409.4]
  input          io_M_AXI_1_RVALID, // @[:@165409.4]
  output         io_M_AXI_1_RREADY, // @[:@165409.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@165409.4]
  input          io_M_AXI_1_BVALID, // @[:@165409.4]
  output         io_M_AXI_1_BREADY, // @[:@165409.4]
  output         io_enable, // @[:@165409.4]
  input          io_done, // @[:@165409.4]
  output         io_reset, // @[:@165409.4]
  output [63:0]  io_argIns_0, // @[:@165409.4]
  output [63:0]  io_argIns_1, // @[:@165409.4]
  input          io_argOuts_0_valid, // @[:@165409.4]
  input  [63:0]  io_argOuts_0_bits, // @[:@165409.4]
  output [63:0]  io_argEchos_0, // @[:@165409.4]
  output         io_memStreams_loads_0_cmd_ready, // @[:@165409.4]
  input          io_memStreams_loads_0_cmd_valid, // @[:@165409.4]
  input  [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@165409.4]
  input  [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@165409.4]
  input          io_memStreams_loads_0_data_ready, // @[:@165409.4]
  output         io_memStreams_loads_0_data_valid, // @[:@165409.4]
  output [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@165409.4]
  output         io_memStreams_stores_0_cmd_ready, // @[:@165409.4]
  input          io_memStreams_stores_0_cmd_valid, // @[:@165409.4]
  input  [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@165409.4]
  input  [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@165409.4]
  output         io_memStreams_stores_0_data_ready, // @[:@165409.4]
  input          io_memStreams_stores_0_data_valid, // @[:@165409.4]
  input  [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@165409.4]
  input          io_memStreams_stores_0_data_bits_wstrb, // @[:@165409.4]
  input          io_memStreams_stores_0_wresp_ready, // @[:@165409.4]
  output         io_memStreams_stores_0_wresp_valid, // @[:@165409.4]
  output         io_memStreams_stores_0_wresp_bits, // @[:@165409.4]
  input          io_heap_0_req_valid, // @[:@165409.4]
  input          io_heap_0_req_bits_allocDealloc, // @[:@165409.4]
  input  [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@165409.4]
  output         io_heap_0_resp_valid, // @[:@165409.4]
  output         io_heap_0_resp_bits_allocDealloc, // @[:@165409.4]
  output [63:0]  io_heap_0_resp_bits_sizeAddr // @[:@165409.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 70:28:@165752.4]
  wire [39:0] fringeCommon_io_raddr; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 70:28:@165752.4]
  wire [39:0] fringeCommon_io_waddr; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_argIns_1; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_argEchos_0; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_memStreams_loads_0_cmd_ready; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_memStreams_loads_0_cmd_valid; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_memStreams_loads_0_cmd_bits_addr; // @[FringeZynq.scala 70:28:@165752.4]
  wire [31:0] fringeCommon_io_memStreams_loads_0_cmd_bits_size; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_memStreams_loads_0_data_ready; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_memStreams_loads_0_data_valid; // @[FringeZynq.scala 70:28:@165752.4]
  wire [31:0] fringeCommon_io_memStreams_loads_0_data_bits_rdata_0; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 70:28:@165752.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 70:28:@165752.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_cmd_ready; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 70:28:@165752.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 70:28:@165752.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_ready; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_rresp_valid; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_rresp_bits_rdata_0; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_rresp_bits_rdata_1; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_rresp_bits_rdata_2; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_rresp_bits_rdata_3; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_rresp_bits_rdata_4; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_rresp_bits_rdata_5; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_rresp_bits_rdata_6; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_0_rresp_bits_rdata_7; // @[FringeZynq.scala 70:28:@165752.4]
  wire [31:0] fringeCommon_io_dram_0_rresp_bits_tag; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_0_wresp_valid; // @[FringeZynq.scala 70:28:@165752.4]
  wire [31:0] fringeCommon_io_dram_0_wresp_bits_tag; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_cmd_ready; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 70:28:@165752.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 70:28:@165752.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_ready; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_rresp_valid; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_rresp_bits_rdata_0; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_rresp_bits_rdata_1; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_rresp_bits_rdata_2; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_rresp_bits_rdata_3; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_rresp_bits_rdata_4; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_rresp_bits_rdata_5; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_rresp_bits_rdata_6; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_dram_1_rresp_bits_rdata_7; // @[FringeZynq.scala 70:28:@165752.4]
  wire [31:0] fringeCommon_io_dram_1_rresp_bits_tag; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_dram_1_wresp_valid; // @[FringeZynq.scala 70:28:@165752.4]
  wire [31:0] fringeCommon_io_dram_1_wresp_bits_tag; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 70:28:@165752.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 70:28:@165752.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 70:28:@165752.4]
  wire  AXI4LiteToRFBridgeZCU_clock; // @[FringeZynq.scala 105:31:@166028.4]
  wire  AXI4LiteToRFBridgeZCU_reset; // @[FringeZynq.scala 105:31:@166028.4]
  wire [39:0] AXI4LiteToRFBridgeZCU_io_S_AXI_AWADDR; // @[FringeZynq.scala 105:31:@166028.4]
  wire [2:0] AXI4LiteToRFBridgeZCU_io_S_AXI_AWPROT; // @[FringeZynq.scala 105:31:@166028.4]
  wire  AXI4LiteToRFBridgeZCU_io_S_AXI_AWVALID; // @[FringeZynq.scala 105:31:@166028.4]
  wire  AXI4LiteToRFBridgeZCU_io_S_AXI_AWREADY; // @[FringeZynq.scala 105:31:@166028.4]
  wire [39:0] AXI4LiteToRFBridgeZCU_io_S_AXI_ARADDR; // @[FringeZynq.scala 105:31:@166028.4]
  wire [2:0] AXI4LiteToRFBridgeZCU_io_S_AXI_ARPROT; // @[FringeZynq.scala 105:31:@166028.4]
  wire  AXI4LiteToRFBridgeZCU_io_S_AXI_ARVALID; // @[FringeZynq.scala 105:31:@166028.4]
  wire  AXI4LiteToRFBridgeZCU_io_S_AXI_ARREADY; // @[FringeZynq.scala 105:31:@166028.4]
  wire [63:0] AXI4LiteToRFBridgeZCU_io_S_AXI_WDATA; // @[FringeZynq.scala 105:31:@166028.4]
  wire [7:0] AXI4LiteToRFBridgeZCU_io_S_AXI_WSTRB; // @[FringeZynq.scala 105:31:@166028.4]
  wire  AXI4LiteToRFBridgeZCU_io_S_AXI_WVALID; // @[FringeZynq.scala 105:31:@166028.4]
  wire  AXI4LiteToRFBridgeZCU_io_S_AXI_WREADY; // @[FringeZynq.scala 105:31:@166028.4]
  wire [63:0] AXI4LiteToRFBridgeZCU_io_S_AXI_RDATA; // @[FringeZynq.scala 105:31:@166028.4]
  wire [1:0] AXI4LiteToRFBridgeZCU_io_S_AXI_RRESP; // @[FringeZynq.scala 105:31:@166028.4]
  wire  AXI4LiteToRFBridgeZCU_io_S_AXI_RVALID; // @[FringeZynq.scala 105:31:@166028.4]
  wire  AXI4LiteToRFBridgeZCU_io_S_AXI_RREADY; // @[FringeZynq.scala 105:31:@166028.4]
  wire [1:0] AXI4LiteToRFBridgeZCU_io_S_AXI_BRESP; // @[FringeZynq.scala 105:31:@166028.4]
  wire  AXI4LiteToRFBridgeZCU_io_S_AXI_BVALID; // @[FringeZynq.scala 105:31:@166028.4]
  wire  AXI4LiteToRFBridgeZCU_io_S_AXI_BREADY; // @[FringeZynq.scala 105:31:@166028.4]
  wire [39:0] AXI4LiteToRFBridgeZCU_io_raddr; // @[FringeZynq.scala 105:31:@166028.4]
  wire  AXI4LiteToRFBridgeZCU_io_wen; // @[FringeZynq.scala 105:31:@166028.4]
  wire [39:0] AXI4LiteToRFBridgeZCU_io_waddr; // @[FringeZynq.scala 105:31:@166028.4]
  wire [63:0] AXI4LiteToRFBridgeZCU_io_wdata; // @[FringeZynq.scala 105:31:@166028.4]
  wire [63:0] AXI4LiteToRFBridgeZCU_io_rdata; // @[FringeZynq.scala 105:31:@166028.4]
  wire  MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_cmd_valid; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_cmd_bits_addr; // @[FringeZynq.scala 136:27:@166133.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_size; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_cmd_bits_isWr; // @[FringeZynq.scala 136:27:@166133.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_tag; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_valid; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wlast; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_rresp_ready; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_rresp_valid; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_0; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_1; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_2; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_3; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_4; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_5; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_6; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_in_rresp_bits_rdata_7; // @[FringeZynq.scala 136:27:@166133.4]
  wire [31:0] MAGToAXI4Bridge_io_in_rresp_bits_tag; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wresp_ready; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 136:27:@166133.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 136:27:@166133.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 136:27:@166133.4]
  wire [39:0] MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 136:27:@166133.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWREADY; // @[FringeZynq.scala 136:27:@166133.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 136:27:@166133.4]
  wire [39:0] MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 136:27:@166133.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARREADY; // @[FringeZynq.scala 136:27:@166133.4]
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 136:27:@166133.4]
  wire [63:0] MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WREADY; // @[FringeZynq.scala 136:27:@166133.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_RID; // @[FringeZynq.scala 136:27:@166133.4]
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_RDATA; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_M_AXI_RVALID; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 136:27:@166133.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_BID; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BVALID; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 136:27:@166133.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_valid; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_cmd_bits_addr; // @[FringeZynq.scala 136:27:@166273.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_size; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_bits_isWr; // @[FringeZynq.scala 136:27:@166273.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_tag; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_valid; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wlast; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_rresp_ready; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_rresp_valid; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_0; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_1; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_2; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_3; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_4; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_5; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_6; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_7; // @[FringeZynq.scala 136:27:@166273.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_rresp_bits_tag; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_ready; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 136:27:@166273.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 136:27:@166273.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 136:27:@166273.4]
  wire [39:0] MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 136:27:@166273.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWREADY; // @[FringeZynq.scala 136:27:@166273.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 136:27:@166273.4]
  wire [39:0] MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 136:27:@166273.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARREADY; // @[FringeZynq.scala 136:27:@166273.4]
  wire [511:0] MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 136:27:@166273.4]
  wire [63:0] MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WREADY; // @[FringeZynq.scala 136:27:@166273.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_RID; // @[FringeZynq.scala 136:27:@166273.4]
  wire [511:0] MAGToAXI4Bridge_1_io_M_AXI_RDATA; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_RVALID; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 136:27:@166273.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_BID; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BVALID; // @[FringeZynq.scala 136:27:@166273.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 136:27:@166273.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 70:28:@165752.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argIns_1(fringeCommon_io_argIns_1),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_argEchos_0(fringeCommon_io_argEchos_0),
    .io_memStreams_loads_0_cmd_ready(fringeCommon_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(fringeCommon_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(fringeCommon_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(fringeCommon_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(fringeCommon_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(fringeCommon_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(fringeCommon_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_stores_0_cmd_ready(fringeCommon_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(fringeCommon_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(fringeCommon_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(fringeCommon_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(fringeCommon_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(fringeCommon_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(fringeCommon_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(fringeCommon_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(fringeCommon_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(fringeCommon_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(fringeCommon_io_memStreams_stores_0_wresp_bits),
    .io_dram_0_cmd_ready(fringeCommon_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(fringeCommon_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(fringeCommon_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(fringeCommon_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_isWr(fringeCommon_io_dram_0_cmd_bits_isWr),
    .io_dram_0_cmd_bits_tag(fringeCommon_io_dram_0_cmd_bits_tag),
    .io_dram_0_wdata_ready(fringeCommon_io_dram_0_wdata_ready),
    .io_dram_0_wdata_valid(fringeCommon_io_dram_0_wdata_valid),
    .io_dram_0_wdata_bits_wdata_0(fringeCommon_io_dram_0_wdata_bits_wdata_0),
    .io_dram_0_wdata_bits_wdata_1(fringeCommon_io_dram_0_wdata_bits_wdata_1),
    .io_dram_0_wdata_bits_wdata_2(fringeCommon_io_dram_0_wdata_bits_wdata_2),
    .io_dram_0_wdata_bits_wdata_3(fringeCommon_io_dram_0_wdata_bits_wdata_3),
    .io_dram_0_wdata_bits_wdata_4(fringeCommon_io_dram_0_wdata_bits_wdata_4),
    .io_dram_0_wdata_bits_wdata_5(fringeCommon_io_dram_0_wdata_bits_wdata_5),
    .io_dram_0_wdata_bits_wdata_6(fringeCommon_io_dram_0_wdata_bits_wdata_6),
    .io_dram_0_wdata_bits_wdata_7(fringeCommon_io_dram_0_wdata_bits_wdata_7),
    .io_dram_0_wdata_bits_wstrb_0(fringeCommon_io_dram_0_wdata_bits_wstrb_0),
    .io_dram_0_wdata_bits_wstrb_1(fringeCommon_io_dram_0_wdata_bits_wstrb_1),
    .io_dram_0_wdata_bits_wstrb_2(fringeCommon_io_dram_0_wdata_bits_wstrb_2),
    .io_dram_0_wdata_bits_wstrb_3(fringeCommon_io_dram_0_wdata_bits_wstrb_3),
    .io_dram_0_wdata_bits_wstrb_4(fringeCommon_io_dram_0_wdata_bits_wstrb_4),
    .io_dram_0_wdata_bits_wstrb_5(fringeCommon_io_dram_0_wdata_bits_wstrb_5),
    .io_dram_0_wdata_bits_wstrb_6(fringeCommon_io_dram_0_wdata_bits_wstrb_6),
    .io_dram_0_wdata_bits_wstrb_7(fringeCommon_io_dram_0_wdata_bits_wstrb_7),
    .io_dram_0_wdata_bits_wstrb_8(fringeCommon_io_dram_0_wdata_bits_wstrb_8),
    .io_dram_0_wdata_bits_wstrb_9(fringeCommon_io_dram_0_wdata_bits_wstrb_9),
    .io_dram_0_wdata_bits_wstrb_10(fringeCommon_io_dram_0_wdata_bits_wstrb_10),
    .io_dram_0_wdata_bits_wstrb_11(fringeCommon_io_dram_0_wdata_bits_wstrb_11),
    .io_dram_0_wdata_bits_wstrb_12(fringeCommon_io_dram_0_wdata_bits_wstrb_12),
    .io_dram_0_wdata_bits_wstrb_13(fringeCommon_io_dram_0_wdata_bits_wstrb_13),
    .io_dram_0_wdata_bits_wstrb_14(fringeCommon_io_dram_0_wdata_bits_wstrb_14),
    .io_dram_0_wdata_bits_wstrb_15(fringeCommon_io_dram_0_wdata_bits_wstrb_15),
    .io_dram_0_wdata_bits_wstrb_16(fringeCommon_io_dram_0_wdata_bits_wstrb_16),
    .io_dram_0_wdata_bits_wstrb_17(fringeCommon_io_dram_0_wdata_bits_wstrb_17),
    .io_dram_0_wdata_bits_wstrb_18(fringeCommon_io_dram_0_wdata_bits_wstrb_18),
    .io_dram_0_wdata_bits_wstrb_19(fringeCommon_io_dram_0_wdata_bits_wstrb_19),
    .io_dram_0_wdata_bits_wstrb_20(fringeCommon_io_dram_0_wdata_bits_wstrb_20),
    .io_dram_0_wdata_bits_wstrb_21(fringeCommon_io_dram_0_wdata_bits_wstrb_21),
    .io_dram_0_wdata_bits_wstrb_22(fringeCommon_io_dram_0_wdata_bits_wstrb_22),
    .io_dram_0_wdata_bits_wstrb_23(fringeCommon_io_dram_0_wdata_bits_wstrb_23),
    .io_dram_0_wdata_bits_wstrb_24(fringeCommon_io_dram_0_wdata_bits_wstrb_24),
    .io_dram_0_wdata_bits_wstrb_25(fringeCommon_io_dram_0_wdata_bits_wstrb_25),
    .io_dram_0_wdata_bits_wstrb_26(fringeCommon_io_dram_0_wdata_bits_wstrb_26),
    .io_dram_0_wdata_bits_wstrb_27(fringeCommon_io_dram_0_wdata_bits_wstrb_27),
    .io_dram_0_wdata_bits_wstrb_28(fringeCommon_io_dram_0_wdata_bits_wstrb_28),
    .io_dram_0_wdata_bits_wstrb_29(fringeCommon_io_dram_0_wdata_bits_wstrb_29),
    .io_dram_0_wdata_bits_wstrb_30(fringeCommon_io_dram_0_wdata_bits_wstrb_30),
    .io_dram_0_wdata_bits_wstrb_31(fringeCommon_io_dram_0_wdata_bits_wstrb_31),
    .io_dram_0_wdata_bits_wstrb_32(fringeCommon_io_dram_0_wdata_bits_wstrb_32),
    .io_dram_0_wdata_bits_wstrb_33(fringeCommon_io_dram_0_wdata_bits_wstrb_33),
    .io_dram_0_wdata_bits_wstrb_34(fringeCommon_io_dram_0_wdata_bits_wstrb_34),
    .io_dram_0_wdata_bits_wstrb_35(fringeCommon_io_dram_0_wdata_bits_wstrb_35),
    .io_dram_0_wdata_bits_wstrb_36(fringeCommon_io_dram_0_wdata_bits_wstrb_36),
    .io_dram_0_wdata_bits_wstrb_37(fringeCommon_io_dram_0_wdata_bits_wstrb_37),
    .io_dram_0_wdata_bits_wstrb_38(fringeCommon_io_dram_0_wdata_bits_wstrb_38),
    .io_dram_0_wdata_bits_wstrb_39(fringeCommon_io_dram_0_wdata_bits_wstrb_39),
    .io_dram_0_wdata_bits_wstrb_40(fringeCommon_io_dram_0_wdata_bits_wstrb_40),
    .io_dram_0_wdata_bits_wstrb_41(fringeCommon_io_dram_0_wdata_bits_wstrb_41),
    .io_dram_0_wdata_bits_wstrb_42(fringeCommon_io_dram_0_wdata_bits_wstrb_42),
    .io_dram_0_wdata_bits_wstrb_43(fringeCommon_io_dram_0_wdata_bits_wstrb_43),
    .io_dram_0_wdata_bits_wstrb_44(fringeCommon_io_dram_0_wdata_bits_wstrb_44),
    .io_dram_0_wdata_bits_wstrb_45(fringeCommon_io_dram_0_wdata_bits_wstrb_45),
    .io_dram_0_wdata_bits_wstrb_46(fringeCommon_io_dram_0_wdata_bits_wstrb_46),
    .io_dram_0_wdata_bits_wstrb_47(fringeCommon_io_dram_0_wdata_bits_wstrb_47),
    .io_dram_0_wdata_bits_wstrb_48(fringeCommon_io_dram_0_wdata_bits_wstrb_48),
    .io_dram_0_wdata_bits_wstrb_49(fringeCommon_io_dram_0_wdata_bits_wstrb_49),
    .io_dram_0_wdata_bits_wstrb_50(fringeCommon_io_dram_0_wdata_bits_wstrb_50),
    .io_dram_0_wdata_bits_wstrb_51(fringeCommon_io_dram_0_wdata_bits_wstrb_51),
    .io_dram_0_wdata_bits_wstrb_52(fringeCommon_io_dram_0_wdata_bits_wstrb_52),
    .io_dram_0_wdata_bits_wstrb_53(fringeCommon_io_dram_0_wdata_bits_wstrb_53),
    .io_dram_0_wdata_bits_wstrb_54(fringeCommon_io_dram_0_wdata_bits_wstrb_54),
    .io_dram_0_wdata_bits_wstrb_55(fringeCommon_io_dram_0_wdata_bits_wstrb_55),
    .io_dram_0_wdata_bits_wstrb_56(fringeCommon_io_dram_0_wdata_bits_wstrb_56),
    .io_dram_0_wdata_bits_wstrb_57(fringeCommon_io_dram_0_wdata_bits_wstrb_57),
    .io_dram_0_wdata_bits_wstrb_58(fringeCommon_io_dram_0_wdata_bits_wstrb_58),
    .io_dram_0_wdata_bits_wstrb_59(fringeCommon_io_dram_0_wdata_bits_wstrb_59),
    .io_dram_0_wdata_bits_wstrb_60(fringeCommon_io_dram_0_wdata_bits_wstrb_60),
    .io_dram_0_wdata_bits_wstrb_61(fringeCommon_io_dram_0_wdata_bits_wstrb_61),
    .io_dram_0_wdata_bits_wstrb_62(fringeCommon_io_dram_0_wdata_bits_wstrb_62),
    .io_dram_0_wdata_bits_wstrb_63(fringeCommon_io_dram_0_wdata_bits_wstrb_63),
    .io_dram_0_wdata_bits_wlast(fringeCommon_io_dram_0_wdata_bits_wlast),
    .io_dram_0_rresp_ready(fringeCommon_io_dram_0_rresp_ready),
    .io_dram_0_rresp_valid(fringeCommon_io_dram_0_rresp_valid),
    .io_dram_0_rresp_bits_rdata_0(fringeCommon_io_dram_0_rresp_bits_rdata_0),
    .io_dram_0_rresp_bits_rdata_1(fringeCommon_io_dram_0_rresp_bits_rdata_1),
    .io_dram_0_rresp_bits_rdata_2(fringeCommon_io_dram_0_rresp_bits_rdata_2),
    .io_dram_0_rresp_bits_rdata_3(fringeCommon_io_dram_0_rresp_bits_rdata_3),
    .io_dram_0_rresp_bits_rdata_4(fringeCommon_io_dram_0_rresp_bits_rdata_4),
    .io_dram_0_rresp_bits_rdata_5(fringeCommon_io_dram_0_rresp_bits_rdata_5),
    .io_dram_0_rresp_bits_rdata_6(fringeCommon_io_dram_0_rresp_bits_rdata_6),
    .io_dram_0_rresp_bits_rdata_7(fringeCommon_io_dram_0_rresp_bits_rdata_7),
    .io_dram_0_rresp_bits_tag(fringeCommon_io_dram_0_rresp_bits_tag),
    .io_dram_0_wresp_ready(fringeCommon_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(fringeCommon_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag(fringeCommon_io_dram_0_wresp_bits_tag),
    .io_dram_1_cmd_ready(fringeCommon_io_dram_1_cmd_ready),
    .io_dram_1_cmd_valid(fringeCommon_io_dram_1_cmd_valid),
    .io_dram_1_cmd_bits_addr(fringeCommon_io_dram_1_cmd_bits_addr),
    .io_dram_1_cmd_bits_size(fringeCommon_io_dram_1_cmd_bits_size),
    .io_dram_1_cmd_bits_isWr(fringeCommon_io_dram_1_cmd_bits_isWr),
    .io_dram_1_cmd_bits_tag(fringeCommon_io_dram_1_cmd_bits_tag),
    .io_dram_1_wdata_ready(fringeCommon_io_dram_1_wdata_ready),
    .io_dram_1_wdata_valid(fringeCommon_io_dram_1_wdata_valid),
    .io_dram_1_wdata_bits_wdata_0(fringeCommon_io_dram_1_wdata_bits_wdata_0),
    .io_dram_1_wdata_bits_wdata_1(fringeCommon_io_dram_1_wdata_bits_wdata_1),
    .io_dram_1_wdata_bits_wdata_2(fringeCommon_io_dram_1_wdata_bits_wdata_2),
    .io_dram_1_wdata_bits_wdata_3(fringeCommon_io_dram_1_wdata_bits_wdata_3),
    .io_dram_1_wdata_bits_wdata_4(fringeCommon_io_dram_1_wdata_bits_wdata_4),
    .io_dram_1_wdata_bits_wdata_5(fringeCommon_io_dram_1_wdata_bits_wdata_5),
    .io_dram_1_wdata_bits_wdata_6(fringeCommon_io_dram_1_wdata_bits_wdata_6),
    .io_dram_1_wdata_bits_wdata_7(fringeCommon_io_dram_1_wdata_bits_wdata_7),
    .io_dram_1_wdata_bits_wstrb_0(fringeCommon_io_dram_1_wdata_bits_wstrb_0),
    .io_dram_1_wdata_bits_wstrb_1(fringeCommon_io_dram_1_wdata_bits_wstrb_1),
    .io_dram_1_wdata_bits_wstrb_2(fringeCommon_io_dram_1_wdata_bits_wstrb_2),
    .io_dram_1_wdata_bits_wstrb_3(fringeCommon_io_dram_1_wdata_bits_wstrb_3),
    .io_dram_1_wdata_bits_wstrb_4(fringeCommon_io_dram_1_wdata_bits_wstrb_4),
    .io_dram_1_wdata_bits_wstrb_5(fringeCommon_io_dram_1_wdata_bits_wstrb_5),
    .io_dram_1_wdata_bits_wstrb_6(fringeCommon_io_dram_1_wdata_bits_wstrb_6),
    .io_dram_1_wdata_bits_wstrb_7(fringeCommon_io_dram_1_wdata_bits_wstrb_7),
    .io_dram_1_wdata_bits_wstrb_8(fringeCommon_io_dram_1_wdata_bits_wstrb_8),
    .io_dram_1_wdata_bits_wstrb_9(fringeCommon_io_dram_1_wdata_bits_wstrb_9),
    .io_dram_1_wdata_bits_wstrb_10(fringeCommon_io_dram_1_wdata_bits_wstrb_10),
    .io_dram_1_wdata_bits_wstrb_11(fringeCommon_io_dram_1_wdata_bits_wstrb_11),
    .io_dram_1_wdata_bits_wstrb_12(fringeCommon_io_dram_1_wdata_bits_wstrb_12),
    .io_dram_1_wdata_bits_wstrb_13(fringeCommon_io_dram_1_wdata_bits_wstrb_13),
    .io_dram_1_wdata_bits_wstrb_14(fringeCommon_io_dram_1_wdata_bits_wstrb_14),
    .io_dram_1_wdata_bits_wstrb_15(fringeCommon_io_dram_1_wdata_bits_wstrb_15),
    .io_dram_1_wdata_bits_wstrb_16(fringeCommon_io_dram_1_wdata_bits_wstrb_16),
    .io_dram_1_wdata_bits_wstrb_17(fringeCommon_io_dram_1_wdata_bits_wstrb_17),
    .io_dram_1_wdata_bits_wstrb_18(fringeCommon_io_dram_1_wdata_bits_wstrb_18),
    .io_dram_1_wdata_bits_wstrb_19(fringeCommon_io_dram_1_wdata_bits_wstrb_19),
    .io_dram_1_wdata_bits_wstrb_20(fringeCommon_io_dram_1_wdata_bits_wstrb_20),
    .io_dram_1_wdata_bits_wstrb_21(fringeCommon_io_dram_1_wdata_bits_wstrb_21),
    .io_dram_1_wdata_bits_wstrb_22(fringeCommon_io_dram_1_wdata_bits_wstrb_22),
    .io_dram_1_wdata_bits_wstrb_23(fringeCommon_io_dram_1_wdata_bits_wstrb_23),
    .io_dram_1_wdata_bits_wstrb_24(fringeCommon_io_dram_1_wdata_bits_wstrb_24),
    .io_dram_1_wdata_bits_wstrb_25(fringeCommon_io_dram_1_wdata_bits_wstrb_25),
    .io_dram_1_wdata_bits_wstrb_26(fringeCommon_io_dram_1_wdata_bits_wstrb_26),
    .io_dram_1_wdata_bits_wstrb_27(fringeCommon_io_dram_1_wdata_bits_wstrb_27),
    .io_dram_1_wdata_bits_wstrb_28(fringeCommon_io_dram_1_wdata_bits_wstrb_28),
    .io_dram_1_wdata_bits_wstrb_29(fringeCommon_io_dram_1_wdata_bits_wstrb_29),
    .io_dram_1_wdata_bits_wstrb_30(fringeCommon_io_dram_1_wdata_bits_wstrb_30),
    .io_dram_1_wdata_bits_wstrb_31(fringeCommon_io_dram_1_wdata_bits_wstrb_31),
    .io_dram_1_wdata_bits_wstrb_32(fringeCommon_io_dram_1_wdata_bits_wstrb_32),
    .io_dram_1_wdata_bits_wstrb_33(fringeCommon_io_dram_1_wdata_bits_wstrb_33),
    .io_dram_1_wdata_bits_wstrb_34(fringeCommon_io_dram_1_wdata_bits_wstrb_34),
    .io_dram_1_wdata_bits_wstrb_35(fringeCommon_io_dram_1_wdata_bits_wstrb_35),
    .io_dram_1_wdata_bits_wstrb_36(fringeCommon_io_dram_1_wdata_bits_wstrb_36),
    .io_dram_1_wdata_bits_wstrb_37(fringeCommon_io_dram_1_wdata_bits_wstrb_37),
    .io_dram_1_wdata_bits_wstrb_38(fringeCommon_io_dram_1_wdata_bits_wstrb_38),
    .io_dram_1_wdata_bits_wstrb_39(fringeCommon_io_dram_1_wdata_bits_wstrb_39),
    .io_dram_1_wdata_bits_wstrb_40(fringeCommon_io_dram_1_wdata_bits_wstrb_40),
    .io_dram_1_wdata_bits_wstrb_41(fringeCommon_io_dram_1_wdata_bits_wstrb_41),
    .io_dram_1_wdata_bits_wstrb_42(fringeCommon_io_dram_1_wdata_bits_wstrb_42),
    .io_dram_1_wdata_bits_wstrb_43(fringeCommon_io_dram_1_wdata_bits_wstrb_43),
    .io_dram_1_wdata_bits_wstrb_44(fringeCommon_io_dram_1_wdata_bits_wstrb_44),
    .io_dram_1_wdata_bits_wstrb_45(fringeCommon_io_dram_1_wdata_bits_wstrb_45),
    .io_dram_1_wdata_bits_wstrb_46(fringeCommon_io_dram_1_wdata_bits_wstrb_46),
    .io_dram_1_wdata_bits_wstrb_47(fringeCommon_io_dram_1_wdata_bits_wstrb_47),
    .io_dram_1_wdata_bits_wstrb_48(fringeCommon_io_dram_1_wdata_bits_wstrb_48),
    .io_dram_1_wdata_bits_wstrb_49(fringeCommon_io_dram_1_wdata_bits_wstrb_49),
    .io_dram_1_wdata_bits_wstrb_50(fringeCommon_io_dram_1_wdata_bits_wstrb_50),
    .io_dram_1_wdata_bits_wstrb_51(fringeCommon_io_dram_1_wdata_bits_wstrb_51),
    .io_dram_1_wdata_bits_wstrb_52(fringeCommon_io_dram_1_wdata_bits_wstrb_52),
    .io_dram_1_wdata_bits_wstrb_53(fringeCommon_io_dram_1_wdata_bits_wstrb_53),
    .io_dram_1_wdata_bits_wstrb_54(fringeCommon_io_dram_1_wdata_bits_wstrb_54),
    .io_dram_1_wdata_bits_wstrb_55(fringeCommon_io_dram_1_wdata_bits_wstrb_55),
    .io_dram_1_wdata_bits_wstrb_56(fringeCommon_io_dram_1_wdata_bits_wstrb_56),
    .io_dram_1_wdata_bits_wstrb_57(fringeCommon_io_dram_1_wdata_bits_wstrb_57),
    .io_dram_1_wdata_bits_wstrb_58(fringeCommon_io_dram_1_wdata_bits_wstrb_58),
    .io_dram_1_wdata_bits_wstrb_59(fringeCommon_io_dram_1_wdata_bits_wstrb_59),
    .io_dram_1_wdata_bits_wstrb_60(fringeCommon_io_dram_1_wdata_bits_wstrb_60),
    .io_dram_1_wdata_bits_wstrb_61(fringeCommon_io_dram_1_wdata_bits_wstrb_61),
    .io_dram_1_wdata_bits_wstrb_62(fringeCommon_io_dram_1_wdata_bits_wstrb_62),
    .io_dram_1_wdata_bits_wstrb_63(fringeCommon_io_dram_1_wdata_bits_wstrb_63),
    .io_dram_1_wdata_bits_wlast(fringeCommon_io_dram_1_wdata_bits_wlast),
    .io_dram_1_rresp_ready(fringeCommon_io_dram_1_rresp_ready),
    .io_dram_1_rresp_valid(fringeCommon_io_dram_1_rresp_valid),
    .io_dram_1_rresp_bits_rdata_0(fringeCommon_io_dram_1_rresp_bits_rdata_0),
    .io_dram_1_rresp_bits_rdata_1(fringeCommon_io_dram_1_rresp_bits_rdata_1),
    .io_dram_1_rresp_bits_rdata_2(fringeCommon_io_dram_1_rresp_bits_rdata_2),
    .io_dram_1_rresp_bits_rdata_3(fringeCommon_io_dram_1_rresp_bits_rdata_3),
    .io_dram_1_rresp_bits_rdata_4(fringeCommon_io_dram_1_rresp_bits_rdata_4),
    .io_dram_1_rresp_bits_rdata_5(fringeCommon_io_dram_1_rresp_bits_rdata_5),
    .io_dram_1_rresp_bits_rdata_6(fringeCommon_io_dram_1_rresp_bits_rdata_6),
    .io_dram_1_rresp_bits_rdata_7(fringeCommon_io_dram_1_rresp_bits_rdata_7),
    .io_dram_1_rresp_bits_tag(fringeCommon_io_dram_1_rresp_bits_tag),
    .io_dram_1_wresp_ready(fringeCommon_io_dram_1_wresp_ready),
    .io_dram_1_wresp_valid(fringeCommon_io_dram_1_wresp_valid),
    .io_dram_1_wresp_bits_tag(fringeCommon_io_dram_1_wresp_bits_tag),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridgeZCU AXI4LiteToRFBridgeZCU ( // @[FringeZynq.scala 105:31:@166028.4]
    .clock(AXI4LiteToRFBridgeZCU_clock),
    .reset(AXI4LiteToRFBridgeZCU_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridgeZCU_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridgeZCU_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridgeZCU_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridgeZCU_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridgeZCU_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridgeZCU_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridgeZCU_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridgeZCU_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridgeZCU_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridgeZCU_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridgeZCU_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridgeZCU_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridgeZCU_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridgeZCU_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridgeZCU_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridgeZCU_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridgeZCU_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridgeZCU_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridgeZCU_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridgeZCU_io_raddr),
    .io_wen(AXI4LiteToRFBridgeZCU_io_wen),
    .io_waddr(AXI4LiteToRFBridgeZCU_io_waddr),
    .io_wdata(AXI4LiteToRFBridgeZCU_io_wdata),
    .io_rdata(AXI4LiteToRFBridgeZCU_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 136:27:@166133.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_io_in_rresp_ready),
    .io_in_rresp_valid(MAGToAXI4Bridge_io_in_rresp_valid),
    .io_in_rresp_bits_rdata_0(MAGToAXI4Bridge_io_in_rresp_bits_rdata_0),
    .io_in_rresp_bits_rdata_1(MAGToAXI4Bridge_io_in_rresp_bits_rdata_1),
    .io_in_rresp_bits_rdata_2(MAGToAXI4Bridge_io_in_rresp_bits_rdata_2),
    .io_in_rresp_bits_rdata_3(MAGToAXI4Bridge_io_in_rresp_bits_rdata_3),
    .io_in_rresp_bits_rdata_4(MAGToAXI4Bridge_io_in_rresp_bits_rdata_4),
    .io_in_rresp_bits_rdata_5(MAGToAXI4Bridge_io_in_rresp_bits_rdata_5),
    .io_in_rresp_bits_rdata_6(MAGToAXI4Bridge_io_in_rresp_bits_rdata_6),
    .io_in_rresp_bits_rdata_7(MAGToAXI4Bridge_io_in_rresp_bits_rdata_7),
    .io_in_rresp_bits_tag(MAGToAXI4Bridge_io_in_rresp_bits_tag),
    .io_in_wresp_ready(MAGToAXI4Bridge_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_io_M_AXI_WREADY),
    .io_M_AXI_RID(MAGToAXI4Bridge_io_M_AXI_RID),
    .io_M_AXI_RDATA(MAGToAXI4Bridge_io_M_AXI_RDATA),
    .io_M_AXI_RVALID(MAGToAXI4Bridge_io_M_AXI_RVALID),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_1 ( // @[FringeZynq.scala 136:27:@166273.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_1_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_1_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_1_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_1_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_1_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_1_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_1_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_1_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_1_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_1_io_in_rresp_ready),
    .io_in_rresp_valid(MAGToAXI4Bridge_1_io_in_rresp_valid),
    .io_in_rresp_bits_rdata_0(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_0),
    .io_in_rresp_bits_rdata_1(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_1),
    .io_in_rresp_bits_rdata_2(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_2),
    .io_in_rresp_bits_rdata_3(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_3),
    .io_in_rresp_bits_rdata_4(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_4),
    .io_in_rresp_bits_rdata_5(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_5),
    .io_in_rresp_bits_rdata_6(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_6),
    .io_in_rresp_bits_rdata_7(MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_7),
    .io_in_rresp_bits_tag(MAGToAXI4Bridge_1_io_in_rresp_bits_tag),
    .io_in_wresp_ready(MAGToAXI4Bridge_1_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_1_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_1_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_1_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_1_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_1_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_1_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_1_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_1_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_1_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_1_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_1_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_1_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_1_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_1_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_1_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_1_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_1_io_M_AXI_WREADY),
    .io_M_AXI_RID(MAGToAXI4Bridge_1_io_M_AXI_RID),
    .io_M_AXI_RDATA(MAGToAXI4Bridge_1_io_M_AXI_RDATA),
    .io_M_AXI_RVALID(MAGToAXI4Bridge_1_io_M_AXI_RVALID),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_1_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_1_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_1_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_1_io_M_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridgeZCU_io_S_AXI_AWREADY; // @[FringeZynq.scala 106:28:@166046.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridgeZCU_io_S_AXI_ARREADY; // @[FringeZynq.scala 106:28:@166042.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridgeZCU_io_S_AXI_WREADY; // @[FringeZynq.scala 106:28:@166038.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridgeZCU_io_S_AXI_RDATA; // @[FringeZynq.scala 106:28:@166037.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridgeZCU_io_S_AXI_RRESP; // @[FringeZynq.scala 106:28:@166036.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridgeZCU_io_S_AXI_RVALID; // @[FringeZynq.scala 106:28:@166035.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridgeZCU_io_S_AXI_BRESP; // @[FringeZynq.scala 106:28:@166033.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridgeZCU_io_S_AXI_BVALID; // @[FringeZynq.scala 106:28:@166032.4]
  assign io_M_AXI_0_AWID = MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 138:10:@166272.4]
  assign io_M_AXI_0_AWADDR = MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 138:10:@166270.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 138:10:@166269.4]
  assign io_M_AXI_0_AWVALID = MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 138:10:@166262.4]
  assign io_M_AXI_0_ARID = MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 138:10:@166260.4]
  assign io_M_AXI_0_ARADDR = MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 138:10:@166258.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 138:10:@166257.4]
  assign io_M_AXI_0_ARVALID = MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 138:10:@166250.4]
  assign io_M_AXI_0_WDATA = MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 138:10:@166248.4]
  assign io_M_AXI_0_WSTRB = MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 138:10:@166247.4]
  assign io_M_AXI_0_WLAST = MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 138:10:@166246.4]
  assign io_M_AXI_0_WVALID = MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 138:10:@166245.4]
  assign io_M_AXI_0_RREADY = MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 138:10:@166237.4]
  assign io_M_AXI_0_BREADY = MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 138:10:@166232.4]
  assign io_M_AXI_1_AWID = MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 138:10:@166412.4]
  assign io_M_AXI_1_AWADDR = MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 138:10:@166410.4]
  assign io_M_AXI_1_AWLEN = MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 138:10:@166409.4]
  assign io_M_AXI_1_AWVALID = MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 138:10:@166402.4]
  assign io_M_AXI_1_ARID = MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 138:10:@166400.4]
  assign io_M_AXI_1_ARADDR = MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 138:10:@166398.4]
  assign io_M_AXI_1_ARLEN = MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 138:10:@166397.4]
  assign io_M_AXI_1_ARVALID = MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 138:10:@166390.4]
  assign io_M_AXI_1_WDATA = MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 138:10:@166388.4]
  assign io_M_AXI_1_WSTRB = MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 138:10:@166387.4]
  assign io_M_AXI_1_WLAST = MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 138:10:@166386.4]
  assign io_M_AXI_1_WVALID = MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 138:10:@166385.4]
  assign io_M_AXI_1_RREADY = MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 138:10:@166377.4]
  assign io_M_AXI_1_BREADY = MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 138:10:@166372.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 120:13:@166058.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 124:12:@166062.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 126:13:@166063.4]
  assign io_argIns_1 = fringeCommon_io_argIns_1; // @[FringeZynq.scala 126:13:@166064.4]
  assign io_argEchos_0 = fringeCommon_io_argEchos_0; // @[FringeZynq.scala 72:28:@166027.4]
  assign io_memStreams_loads_0_cmd_ready = fringeCommon_io_memStreams_loads_0_cmd_ready; // @[FringeZynq.scala 131:17:@166126.4]
  assign io_memStreams_loads_0_data_valid = fringeCommon_io_memStreams_loads_0_data_valid; // @[FringeZynq.scala 131:17:@166121.4]
  assign io_memStreams_loads_0_data_bits_rdata_0 = fringeCommon_io_memStreams_loads_0_data_bits_rdata_0; // @[FringeZynq.scala 131:17:@166120.4]
  assign io_memStreams_stores_0_cmd_ready = fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 131:17:@166119.4]
  assign io_memStreams_stores_0_data_ready = fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 131:17:@166115.4]
  assign io_memStreams_stores_0_wresp_valid = fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 131:17:@166110.4]
  assign io_memStreams_stores_0_wresp_bits = fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 131:17:@166109.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 132:11:@166129.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 132:11:@166128.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 132:11:@166127.4]
  assign fringeCommon_clock = clock; // @[:@165753.4]
  assign fringeCommon_reset = reset; // @[:@165754.4 FringeZynq.scala 122:22:@166061.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridgeZCU_io_raddr; // @[FringeZynq.scala 110:27:@166052.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridgeZCU_io_wen; // @[FringeZynq.scala 111:27:@166053.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridgeZCU_io_waddr; // @[FringeZynq.scala 112:27:@166054.4]
  assign fringeCommon_io_wdata = AXI4LiteToRFBridgeZCU_io_wdata; // @[FringeZynq.scala 113:27:@166055.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 121:24:@166059.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 127:27:@166066.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 127:27:@166065.4]
  assign fringeCommon_io_memStreams_loads_0_cmd_valid = io_memStreams_loads_0_cmd_valid; // @[FringeZynq.scala 131:17:@166125.4]
  assign fringeCommon_io_memStreams_loads_0_cmd_bits_addr = io_memStreams_loads_0_cmd_bits_addr; // @[FringeZynq.scala 131:17:@166124.4]
  assign fringeCommon_io_memStreams_loads_0_cmd_bits_size = io_memStreams_loads_0_cmd_bits_size; // @[FringeZynq.scala 131:17:@166123.4]
  assign fringeCommon_io_memStreams_loads_0_data_ready = io_memStreams_loads_0_data_ready; // @[FringeZynq.scala 131:17:@166122.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 131:17:@166118.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 131:17:@166117.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 131:17:@166116.4]
  assign fringeCommon_io_memStreams_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 131:17:@166114.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 131:17:@166113.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 131:17:@166112.4]
  assign fringeCommon_io_memStreams_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 131:17:@166111.4]
  assign fringeCommon_io_dram_0_cmd_ready = MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 137:21:@166231.4]
  assign fringeCommon_io_dram_0_wdata_ready = MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 137:21:@166224.4]
  assign fringeCommon_io_dram_0_rresp_valid = MAGToAXI4Bridge_io_in_rresp_valid; // @[FringeZynq.scala 137:21:@166148.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_0 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_0; // @[FringeZynq.scala 137:21:@166140.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_1 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_1; // @[FringeZynq.scala 137:21:@166141.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_2 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_2; // @[FringeZynq.scala 137:21:@166142.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_3 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_3; // @[FringeZynq.scala 137:21:@166143.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_4 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_4; // @[FringeZynq.scala 137:21:@166144.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_5 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_5; // @[FringeZynq.scala 137:21:@166145.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_6 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_6; // @[FringeZynq.scala 137:21:@166146.4]
  assign fringeCommon_io_dram_0_rresp_bits_rdata_7 = MAGToAXI4Bridge_io_in_rresp_bits_rdata_7; // @[FringeZynq.scala 137:21:@166147.4]
  assign fringeCommon_io_dram_0_rresp_bits_tag = MAGToAXI4Bridge_io_in_rresp_bits_tag; // @[FringeZynq.scala 137:21:@166139.4]
  assign fringeCommon_io_dram_0_wresp_valid = MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 137:21:@166137.4]
  assign fringeCommon_io_dram_0_wresp_bits_tag = MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 137:21:@166136.4]
  assign fringeCommon_io_dram_1_cmd_ready = MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 137:21:@166371.4]
  assign fringeCommon_io_dram_1_wdata_ready = MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 137:21:@166364.4]
  assign fringeCommon_io_dram_1_rresp_valid = MAGToAXI4Bridge_1_io_in_rresp_valid; // @[FringeZynq.scala 137:21:@166288.4]
  assign fringeCommon_io_dram_1_rresp_bits_rdata_0 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_0; // @[FringeZynq.scala 137:21:@166280.4]
  assign fringeCommon_io_dram_1_rresp_bits_rdata_1 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_1; // @[FringeZynq.scala 137:21:@166281.4]
  assign fringeCommon_io_dram_1_rresp_bits_rdata_2 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_2; // @[FringeZynq.scala 137:21:@166282.4]
  assign fringeCommon_io_dram_1_rresp_bits_rdata_3 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_3; // @[FringeZynq.scala 137:21:@166283.4]
  assign fringeCommon_io_dram_1_rresp_bits_rdata_4 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_4; // @[FringeZynq.scala 137:21:@166284.4]
  assign fringeCommon_io_dram_1_rresp_bits_rdata_5 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_5; // @[FringeZynq.scala 137:21:@166285.4]
  assign fringeCommon_io_dram_1_rresp_bits_rdata_6 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_6; // @[FringeZynq.scala 137:21:@166286.4]
  assign fringeCommon_io_dram_1_rresp_bits_rdata_7 = MAGToAXI4Bridge_1_io_in_rresp_bits_rdata_7; // @[FringeZynq.scala 137:21:@166287.4]
  assign fringeCommon_io_dram_1_rresp_bits_tag = MAGToAXI4Bridge_1_io_in_rresp_bits_tag; // @[FringeZynq.scala 137:21:@166279.4]
  assign fringeCommon_io_dram_1_wresp_valid = MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 137:21:@166277.4]
  assign fringeCommon_io_dram_1_wresp_bits_tag = MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 137:21:@166276.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 132:11:@166132.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 132:11:@166131.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 132:11:@166130.4]
  assign AXI4LiteToRFBridgeZCU_clock = io_axil_s_clk; // @[:@166029.4 FringeZynq.scala 107:25:@166051.4]
  assign AXI4LiteToRFBridgeZCU_reset = reset; // @[:@166030.4]
  assign AXI4LiteToRFBridgeZCU_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 106:28:@166049.4]
  assign AXI4LiteToRFBridgeZCU_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 106:28:@166048.4]
  assign AXI4LiteToRFBridgeZCU_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 106:28:@166047.4]
  assign AXI4LiteToRFBridgeZCU_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 106:28:@166045.4]
  assign AXI4LiteToRFBridgeZCU_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 106:28:@166044.4]
  assign AXI4LiteToRFBridgeZCU_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 106:28:@166043.4]
  assign AXI4LiteToRFBridgeZCU_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 106:28:@166041.4]
  assign AXI4LiteToRFBridgeZCU_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 106:28:@166040.4]
  assign AXI4LiteToRFBridgeZCU_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 106:28:@166039.4]
  assign AXI4LiteToRFBridgeZCU_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 106:28:@166034.4]
  assign AXI4LiteToRFBridgeZCU_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 106:28:@166031.4]
  assign AXI4LiteToRFBridgeZCU_io_rdata = fringeCommon_io_rdata; // @[FringeZynq.scala 114:28:@166056.4]
  assign MAGToAXI4Bridge_io_in_cmd_valid = fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 137:21:@166230.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_addr = fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 137:21:@166229.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_size = fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 137:21:@166228.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_isWr = fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 137:21:@166226.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag = fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 137:21:@166225.4]
  assign MAGToAXI4Bridge_io_in_wdata_valid = fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 137:21:@166223.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 137:21:@166215.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 137:21:@166216.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 137:21:@166217.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 137:21:@166218.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 137:21:@166219.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 137:21:@166220.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 137:21:@166221.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 137:21:@166222.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 137:21:@166151.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 137:21:@166152.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 137:21:@166153.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 137:21:@166154.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 137:21:@166155.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 137:21:@166156.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 137:21:@166157.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 137:21:@166158.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 137:21:@166159.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 137:21:@166160.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 137:21:@166161.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 137:21:@166162.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 137:21:@166163.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 137:21:@166164.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 137:21:@166165.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 137:21:@166166.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 137:21:@166167.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 137:21:@166168.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 137:21:@166169.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 137:21:@166170.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 137:21:@166171.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 137:21:@166172.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 137:21:@166173.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 137:21:@166174.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 137:21:@166175.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 137:21:@166176.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 137:21:@166177.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 137:21:@166178.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 137:21:@166179.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 137:21:@166180.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 137:21:@166181.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 137:21:@166182.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 137:21:@166183.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 137:21:@166184.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 137:21:@166185.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 137:21:@166186.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 137:21:@166187.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 137:21:@166188.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 137:21:@166189.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 137:21:@166190.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 137:21:@166191.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 137:21:@166192.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 137:21:@166193.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 137:21:@166194.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 137:21:@166195.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 137:21:@166196.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 137:21:@166197.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 137:21:@166198.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 137:21:@166199.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 137:21:@166200.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 137:21:@166201.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 137:21:@166202.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 137:21:@166203.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 137:21:@166204.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 137:21:@166205.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 137:21:@166206.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 137:21:@166207.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 137:21:@166208.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 137:21:@166209.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 137:21:@166210.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 137:21:@166211.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 137:21:@166212.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 137:21:@166213.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 137:21:@166214.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wlast = fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 137:21:@166150.4]
  assign MAGToAXI4Bridge_io_in_rresp_ready = fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 137:21:@166149.4]
  assign MAGToAXI4Bridge_io_in_wresp_ready = fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 137:21:@166138.4]
  assign MAGToAXI4Bridge_io_M_AXI_AWREADY = io_M_AXI_0_AWREADY; // @[FringeZynq.scala 138:10:@166261.4]
  assign MAGToAXI4Bridge_io_M_AXI_ARREADY = io_M_AXI_0_ARREADY; // @[FringeZynq.scala 138:10:@166249.4]
  assign MAGToAXI4Bridge_io_M_AXI_WREADY = io_M_AXI_0_WREADY; // @[FringeZynq.scala 138:10:@166244.4]
  assign MAGToAXI4Bridge_io_M_AXI_RID = io_M_AXI_0_RID; // @[FringeZynq.scala 138:10:@166243.4]
  assign MAGToAXI4Bridge_io_M_AXI_RDATA = io_M_AXI_0_RDATA; // @[FringeZynq.scala 138:10:@166241.4]
  assign MAGToAXI4Bridge_io_M_AXI_RVALID = io_M_AXI_0_RVALID; // @[FringeZynq.scala 138:10:@166238.4]
  assign MAGToAXI4Bridge_io_M_AXI_BID = io_M_AXI_0_BID; // @[FringeZynq.scala 138:10:@166236.4]
  assign MAGToAXI4Bridge_io_M_AXI_BVALID = io_M_AXI_0_BVALID; // @[FringeZynq.scala 138:10:@166233.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_valid = fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 137:21:@166370.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_addr = fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 137:21:@166369.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_size = fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 137:21:@166368.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_isWr = fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 137:21:@166366.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_tag = fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 137:21:@166365.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_valid = fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 137:21:@166363.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 137:21:@166355.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 137:21:@166356.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 137:21:@166357.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 137:21:@166358.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 137:21:@166359.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 137:21:@166360.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 137:21:@166361.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 137:21:@166362.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 137:21:@166291.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 137:21:@166292.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 137:21:@166293.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 137:21:@166294.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 137:21:@166295.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 137:21:@166296.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 137:21:@166297.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 137:21:@166298.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 137:21:@166299.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 137:21:@166300.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 137:21:@166301.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 137:21:@166302.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 137:21:@166303.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 137:21:@166304.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 137:21:@166305.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 137:21:@166306.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 137:21:@166307.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 137:21:@166308.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 137:21:@166309.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 137:21:@166310.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 137:21:@166311.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 137:21:@166312.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 137:21:@166313.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 137:21:@166314.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 137:21:@166315.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 137:21:@166316.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 137:21:@166317.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 137:21:@166318.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 137:21:@166319.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 137:21:@166320.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 137:21:@166321.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 137:21:@166322.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 137:21:@166323.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 137:21:@166324.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 137:21:@166325.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 137:21:@166326.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 137:21:@166327.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 137:21:@166328.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 137:21:@166329.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 137:21:@166330.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 137:21:@166331.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 137:21:@166332.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 137:21:@166333.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 137:21:@166334.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 137:21:@166335.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 137:21:@166336.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 137:21:@166337.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 137:21:@166338.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 137:21:@166339.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 137:21:@166340.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 137:21:@166341.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 137:21:@166342.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 137:21:@166343.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 137:21:@166344.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 137:21:@166345.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 137:21:@166346.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 137:21:@166347.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 137:21:@166348.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 137:21:@166349.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 137:21:@166350.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 137:21:@166351.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 137:21:@166352.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 137:21:@166353.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 137:21:@166354.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wlast = fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 137:21:@166290.4]
  assign MAGToAXI4Bridge_1_io_in_rresp_ready = fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 137:21:@166289.4]
  assign MAGToAXI4Bridge_1_io_in_wresp_ready = fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 137:21:@166278.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_AWREADY = io_M_AXI_1_AWREADY; // @[FringeZynq.scala 138:10:@166401.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_ARREADY = io_M_AXI_1_ARREADY; // @[FringeZynq.scala 138:10:@166389.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_WREADY = io_M_AXI_1_WREADY; // @[FringeZynq.scala 138:10:@166384.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_RID = io_M_AXI_1_RID; // @[FringeZynq.scala 138:10:@166383.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_RDATA = io_M_AXI_1_RDATA; // @[FringeZynq.scala 138:10:@166381.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_RVALID = io_M_AXI_1_RVALID; // @[FringeZynq.scala 138:10:@166378.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BID = io_M_AXI_1_BID; // @[FringeZynq.scala 138:10:@166376.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BVALID = io_M_AXI_1_BVALID; // @[FringeZynq.scala 138:10:@166373.4]
endmodule
module SpatialIP( // @[:@166414.2]
  input          clock, // @[:@166415.4]
  input          reset, // @[:@166416.4]
  input          io_raddr, // @[:@166417.4]
  input          io_wen, // @[:@166417.4]
  input          io_waddr, // @[:@166417.4]
  input          io_wdata, // @[:@166417.4]
  output         io_rdata, // @[:@166417.4]
  input          io_axil_s_clk, // @[:@166417.4]
  input  [39:0]  io_S_AXI_AWADDR, // @[:@166417.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@166417.4]
  input          io_S_AXI_AWVALID, // @[:@166417.4]
  output         io_S_AXI_AWREADY, // @[:@166417.4]
  input  [39:0]  io_S_AXI_ARADDR, // @[:@166417.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@166417.4]
  input          io_S_AXI_ARVALID, // @[:@166417.4]
  output         io_S_AXI_ARREADY, // @[:@166417.4]
  input  [63:0]  io_S_AXI_WDATA, // @[:@166417.4]
  input  [7:0]   io_S_AXI_WSTRB, // @[:@166417.4]
  input          io_S_AXI_WVALID, // @[:@166417.4]
  output         io_S_AXI_WREADY, // @[:@166417.4]
  output [63:0]  io_S_AXI_RDATA, // @[:@166417.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@166417.4]
  output         io_S_AXI_RVALID, // @[:@166417.4]
  input          io_S_AXI_RREADY, // @[:@166417.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@166417.4]
  output         io_S_AXI_BVALID, // @[:@166417.4]
  input          io_S_AXI_BREADY, // @[:@166417.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@166417.4]
  output [31:0]  io_M_AXI_0_AWUSER, // @[:@166417.4]
  output [39:0]  io_M_AXI_0_AWADDR, // @[:@166417.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@166417.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@166417.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@166417.4]
  output         io_M_AXI_0_AWLOCK, // @[:@166417.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@166417.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@166417.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@166417.4]
  output         io_M_AXI_0_AWVALID, // @[:@166417.4]
  input          io_M_AXI_0_AWREADY, // @[:@166417.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@166417.4]
  output [31:0]  io_M_AXI_0_ARUSER, // @[:@166417.4]
  output [39:0]  io_M_AXI_0_ARADDR, // @[:@166417.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@166417.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@166417.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@166417.4]
  output         io_M_AXI_0_ARLOCK, // @[:@166417.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@166417.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@166417.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@166417.4]
  output         io_M_AXI_0_ARVALID, // @[:@166417.4]
  input          io_M_AXI_0_ARREADY, // @[:@166417.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@166417.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@166417.4]
  output         io_M_AXI_0_WLAST, // @[:@166417.4]
  output         io_M_AXI_0_WVALID, // @[:@166417.4]
  input          io_M_AXI_0_WREADY, // @[:@166417.4]
  input  [31:0]  io_M_AXI_0_RID, // @[:@166417.4]
  input  [39:0]  io_M_AXI_0_RUSER, // @[:@166417.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@166417.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@166417.4]
  input          io_M_AXI_0_RLAST, // @[:@166417.4]
  input          io_M_AXI_0_RVALID, // @[:@166417.4]
  output         io_M_AXI_0_RREADY, // @[:@166417.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@166417.4]
  input  [31:0]  io_M_AXI_0_BUSER, // @[:@166417.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@166417.4]
  input          io_M_AXI_0_BVALID, // @[:@166417.4]
  output         io_M_AXI_0_BREADY, // @[:@166417.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@166417.4]
  output [31:0]  io_M_AXI_1_AWUSER, // @[:@166417.4]
  output [39:0]  io_M_AXI_1_AWADDR, // @[:@166417.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@166417.4]
  output [2:0]   io_M_AXI_1_AWSIZE, // @[:@166417.4]
  output [1:0]   io_M_AXI_1_AWBURST, // @[:@166417.4]
  output         io_M_AXI_1_AWLOCK, // @[:@166417.4]
  output [3:0]   io_M_AXI_1_AWCACHE, // @[:@166417.4]
  output [2:0]   io_M_AXI_1_AWPROT, // @[:@166417.4]
  output [3:0]   io_M_AXI_1_AWQOS, // @[:@166417.4]
  output         io_M_AXI_1_AWVALID, // @[:@166417.4]
  input          io_M_AXI_1_AWREADY, // @[:@166417.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@166417.4]
  output [31:0]  io_M_AXI_1_ARUSER, // @[:@166417.4]
  output [39:0]  io_M_AXI_1_ARADDR, // @[:@166417.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@166417.4]
  output [2:0]   io_M_AXI_1_ARSIZE, // @[:@166417.4]
  output [1:0]   io_M_AXI_1_ARBURST, // @[:@166417.4]
  output         io_M_AXI_1_ARLOCK, // @[:@166417.4]
  output [3:0]   io_M_AXI_1_ARCACHE, // @[:@166417.4]
  output [2:0]   io_M_AXI_1_ARPROT, // @[:@166417.4]
  output [3:0]   io_M_AXI_1_ARQOS, // @[:@166417.4]
  output         io_M_AXI_1_ARVALID, // @[:@166417.4]
  input          io_M_AXI_1_ARREADY, // @[:@166417.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@166417.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@166417.4]
  output         io_M_AXI_1_WLAST, // @[:@166417.4]
  output         io_M_AXI_1_WVALID, // @[:@166417.4]
  input          io_M_AXI_1_WREADY, // @[:@166417.4]
  input  [31:0]  io_M_AXI_1_RID, // @[:@166417.4]
  input  [39:0]  io_M_AXI_1_RUSER, // @[:@166417.4]
  input  [511:0] io_M_AXI_1_RDATA, // @[:@166417.4]
  input  [1:0]   io_M_AXI_1_RRESP, // @[:@166417.4]
  input          io_M_AXI_1_RLAST, // @[:@166417.4]
  input          io_M_AXI_1_RVALID, // @[:@166417.4]
  output         io_M_AXI_1_RREADY, // @[:@166417.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@166417.4]
  input  [31:0]  io_M_AXI_1_BUSER, // @[:@166417.4]
  input  [1:0]   io_M_AXI_1_BRESP, // @[:@166417.4]
  input          io_M_AXI_1_BVALID, // @[:@166417.4]
  output         io_M_AXI_1_BREADY, // @[:@166417.4]
  input          io_TOP_AXI_AWID, // @[:@166417.4]
  input          io_TOP_AXI_AWUSER, // @[:@166417.4]
  input  [39:0]  io_TOP_AXI_AWADDR, // @[:@166417.4]
  input  [7:0]   io_TOP_AXI_AWLEN, // @[:@166417.4]
  input  [2:0]   io_TOP_AXI_AWSIZE, // @[:@166417.4]
  input  [1:0]   io_TOP_AXI_AWBURST, // @[:@166417.4]
  input          io_TOP_AXI_AWLOCK, // @[:@166417.4]
  input  [3:0]   io_TOP_AXI_AWCACHE, // @[:@166417.4]
  input  [2:0]   io_TOP_AXI_AWPROT, // @[:@166417.4]
  input  [3:0]   io_TOP_AXI_AWQOS, // @[:@166417.4]
  input          io_TOP_AXI_AWVALID, // @[:@166417.4]
  input          io_TOP_AXI_AWREADY, // @[:@166417.4]
  input          io_TOP_AXI_ARID, // @[:@166417.4]
  input          io_TOP_AXI_ARUSER, // @[:@166417.4]
  input  [39:0]  io_TOP_AXI_ARADDR, // @[:@166417.4]
  input  [7:0]   io_TOP_AXI_ARLEN, // @[:@166417.4]
  input  [2:0]   io_TOP_AXI_ARSIZE, // @[:@166417.4]
  input  [1:0]   io_TOP_AXI_ARBURST, // @[:@166417.4]
  input          io_TOP_AXI_ARLOCK, // @[:@166417.4]
  input  [3:0]   io_TOP_AXI_ARCACHE, // @[:@166417.4]
  input  [2:0]   io_TOP_AXI_ARPROT, // @[:@166417.4]
  input  [3:0]   io_TOP_AXI_ARQOS, // @[:@166417.4]
  input          io_TOP_AXI_ARVALID, // @[:@166417.4]
  input          io_TOP_AXI_ARREADY, // @[:@166417.4]
  input  [63:0]  io_TOP_AXI_WDATA, // @[:@166417.4]
  input  [63:0]  io_TOP_AXI_WSTRB, // @[:@166417.4]
  input          io_TOP_AXI_WLAST, // @[:@166417.4]
  input          io_TOP_AXI_WVALID, // @[:@166417.4]
  input          io_TOP_AXI_WREADY, // @[:@166417.4]
  input          io_TOP_AXI_RID, // @[:@166417.4]
  input          io_TOP_AXI_RUSER, // @[:@166417.4]
  input  [63:0]  io_TOP_AXI_RDATA, // @[:@166417.4]
  input  [1:0]   io_TOP_AXI_RRESP, // @[:@166417.4]
  input          io_TOP_AXI_RLAST, // @[:@166417.4]
  input          io_TOP_AXI_RVALID, // @[:@166417.4]
  input          io_TOP_AXI_RREADY, // @[:@166417.4]
  input          io_TOP_AXI_BID, // @[:@166417.4]
  input          io_TOP_AXI_BUSER, // @[:@166417.4]
  input  [1:0]   io_TOP_AXI_BRESP, // @[:@166417.4]
  input          io_TOP_AXI_BVALID, // @[:@166417.4]
  input          io_TOP_AXI_BREADY, // @[:@166417.4]
  input          io_DWIDTH_AXI_AWID, // @[:@166417.4]
  input          io_DWIDTH_AXI_AWUSER, // @[:@166417.4]
  input  [39:0]  io_DWIDTH_AXI_AWADDR, // @[:@166417.4]
  input  [7:0]   io_DWIDTH_AXI_AWLEN, // @[:@166417.4]
  input  [2:0]   io_DWIDTH_AXI_AWSIZE, // @[:@166417.4]
  input  [1:0]   io_DWIDTH_AXI_AWBURST, // @[:@166417.4]
  input          io_DWIDTH_AXI_AWLOCK, // @[:@166417.4]
  input  [3:0]   io_DWIDTH_AXI_AWCACHE, // @[:@166417.4]
  input  [2:0]   io_DWIDTH_AXI_AWPROT, // @[:@166417.4]
  input  [3:0]   io_DWIDTH_AXI_AWQOS, // @[:@166417.4]
  input          io_DWIDTH_AXI_AWVALID, // @[:@166417.4]
  input          io_DWIDTH_AXI_AWREADY, // @[:@166417.4]
  input          io_DWIDTH_AXI_ARID, // @[:@166417.4]
  input          io_DWIDTH_AXI_ARUSER, // @[:@166417.4]
  input  [39:0]  io_DWIDTH_AXI_ARADDR, // @[:@166417.4]
  input  [7:0]   io_DWIDTH_AXI_ARLEN, // @[:@166417.4]
  input  [2:0]   io_DWIDTH_AXI_ARSIZE, // @[:@166417.4]
  input  [1:0]   io_DWIDTH_AXI_ARBURST, // @[:@166417.4]
  input          io_DWIDTH_AXI_ARLOCK, // @[:@166417.4]
  input  [3:0]   io_DWIDTH_AXI_ARCACHE, // @[:@166417.4]
  input  [2:0]   io_DWIDTH_AXI_ARPROT, // @[:@166417.4]
  input  [3:0]   io_DWIDTH_AXI_ARQOS, // @[:@166417.4]
  input          io_DWIDTH_AXI_ARVALID, // @[:@166417.4]
  input          io_DWIDTH_AXI_ARREADY, // @[:@166417.4]
  input  [63:0]  io_DWIDTH_AXI_WDATA, // @[:@166417.4]
  input  [63:0]  io_DWIDTH_AXI_WSTRB, // @[:@166417.4]
  input          io_DWIDTH_AXI_WLAST, // @[:@166417.4]
  input          io_DWIDTH_AXI_WVALID, // @[:@166417.4]
  input          io_DWIDTH_AXI_WREADY, // @[:@166417.4]
  input          io_DWIDTH_AXI_RID, // @[:@166417.4]
  input          io_DWIDTH_AXI_RUSER, // @[:@166417.4]
  input  [63:0]  io_DWIDTH_AXI_RDATA, // @[:@166417.4]
  input  [1:0]   io_DWIDTH_AXI_RRESP, // @[:@166417.4]
  input          io_DWIDTH_AXI_RLAST, // @[:@166417.4]
  input          io_DWIDTH_AXI_RVALID, // @[:@166417.4]
  input          io_DWIDTH_AXI_RREADY, // @[:@166417.4]
  input          io_DWIDTH_AXI_BID, // @[:@166417.4]
  input          io_DWIDTH_AXI_BUSER, // @[:@166417.4]
  input  [1:0]   io_DWIDTH_AXI_BRESP, // @[:@166417.4]
  input          io_DWIDTH_AXI_BVALID, // @[:@166417.4]
  input          io_DWIDTH_AXI_BREADY, // @[:@166417.4]
  input          io_PROTOCOL_AXI_AWID, // @[:@166417.4]
  input          io_PROTOCOL_AXI_AWUSER, // @[:@166417.4]
  input  [39:0]  io_PROTOCOL_AXI_AWADDR, // @[:@166417.4]
  input  [7:0]   io_PROTOCOL_AXI_AWLEN, // @[:@166417.4]
  input  [2:0]   io_PROTOCOL_AXI_AWSIZE, // @[:@166417.4]
  input  [1:0]   io_PROTOCOL_AXI_AWBURST, // @[:@166417.4]
  input          io_PROTOCOL_AXI_AWLOCK, // @[:@166417.4]
  input  [3:0]   io_PROTOCOL_AXI_AWCACHE, // @[:@166417.4]
  input  [2:0]   io_PROTOCOL_AXI_AWPROT, // @[:@166417.4]
  input  [3:0]   io_PROTOCOL_AXI_AWQOS, // @[:@166417.4]
  input          io_PROTOCOL_AXI_AWVALID, // @[:@166417.4]
  input          io_PROTOCOL_AXI_AWREADY, // @[:@166417.4]
  input          io_PROTOCOL_AXI_ARID, // @[:@166417.4]
  input          io_PROTOCOL_AXI_ARUSER, // @[:@166417.4]
  input  [39:0]  io_PROTOCOL_AXI_ARADDR, // @[:@166417.4]
  input  [7:0]   io_PROTOCOL_AXI_ARLEN, // @[:@166417.4]
  input  [2:0]   io_PROTOCOL_AXI_ARSIZE, // @[:@166417.4]
  input  [1:0]   io_PROTOCOL_AXI_ARBURST, // @[:@166417.4]
  input          io_PROTOCOL_AXI_ARLOCK, // @[:@166417.4]
  input  [3:0]   io_PROTOCOL_AXI_ARCACHE, // @[:@166417.4]
  input  [2:0]   io_PROTOCOL_AXI_ARPROT, // @[:@166417.4]
  input  [3:0]   io_PROTOCOL_AXI_ARQOS, // @[:@166417.4]
  input          io_PROTOCOL_AXI_ARVALID, // @[:@166417.4]
  input          io_PROTOCOL_AXI_ARREADY, // @[:@166417.4]
  input  [63:0]  io_PROTOCOL_AXI_WDATA, // @[:@166417.4]
  input  [63:0]  io_PROTOCOL_AXI_WSTRB, // @[:@166417.4]
  input          io_PROTOCOL_AXI_WLAST, // @[:@166417.4]
  input          io_PROTOCOL_AXI_WVALID, // @[:@166417.4]
  input          io_PROTOCOL_AXI_WREADY, // @[:@166417.4]
  input          io_PROTOCOL_AXI_RID, // @[:@166417.4]
  input          io_PROTOCOL_AXI_RUSER, // @[:@166417.4]
  input  [63:0]  io_PROTOCOL_AXI_RDATA, // @[:@166417.4]
  input  [1:0]   io_PROTOCOL_AXI_RRESP, // @[:@166417.4]
  input          io_PROTOCOL_AXI_RLAST, // @[:@166417.4]
  input          io_PROTOCOL_AXI_RVALID, // @[:@166417.4]
  input          io_PROTOCOL_AXI_RREADY, // @[:@166417.4]
  input          io_PROTOCOL_AXI_BID, // @[:@166417.4]
  input          io_PROTOCOL_AXI_BUSER, // @[:@166417.4]
  input  [1:0]   io_PROTOCOL_AXI_BRESP, // @[:@166417.4]
  input          io_PROTOCOL_AXI_BVALID, // @[:@166417.4]
  input          io_PROTOCOL_AXI_BREADY, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_AWID, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_AWUSER, // @[:@166417.4]
  input  [39:0]  io_CLOCKCONVERT_AXI_AWADDR, // @[:@166417.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_AWLEN, // @[:@166417.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWSIZE, // @[:@166417.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_AWBURST, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_AWLOCK, // @[:@166417.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWCACHE, // @[:@166417.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWPROT, // @[:@166417.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWQOS, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_AWVALID, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_AWREADY, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_ARID, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_ARUSER, // @[:@166417.4]
  input  [39:0]  io_CLOCKCONVERT_AXI_ARADDR, // @[:@166417.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_ARLEN, // @[:@166417.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARSIZE, // @[:@166417.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_ARBURST, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_ARLOCK, // @[:@166417.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARCACHE, // @[:@166417.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARPROT, // @[:@166417.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARQOS, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_ARVALID, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_ARREADY, // @[:@166417.4]
  input  [63:0]  io_CLOCKCONVERT_AXI_WDATA, // @[:@166417.4]
  input  [63:0]  io_CLOCKCONVERT_AXI_WSTRB, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_WLAST, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_WVALID, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_WREADY, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_RID, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_RUSER, // @[:@166417.4]
  input  [63:0]  io_CLOCKCONVERT_AXI_RDATA, // @[:@166417.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_RRESP, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_RLAST, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_RVALID, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_RREADY, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_BID, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_BUSER, // @[:@166417.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_BRESP, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_BVALID, // @[:@166417.4]
  input          io_CLOCKCONVERT_AXI_BREADY // @[:@166417.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@166419.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@166419.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@166419.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@166419.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@166419.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@166419.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@166419.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@166419.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@166419.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@166419.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@166419.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@166419.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@166419.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@166419.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@166419.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@166419.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@166419.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@166419.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@166419.4]
  wire  FringeZynq_clock; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_reset; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_axil_s_clk; // @[Zynq.scala 18:24:@166514.4]
  wire [39:0] FringeZynq_io_S_AXI_AWADDR; // @[Zynq.scala 18:24:@166514.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 18:24:@166514.4]
  wire [39:0] FringeZynq_io_S_AXI_ARADDR; // @[Zynq.scala 18:24:@166514.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 18:24:@166514.4]
  wire [63:0] FringeZynq_io_S_AXI_WDATA; // @[Zynq.scala 18:24:@166514.4]
  wire [7:0] FringeZynq_io_S_AXI_WSTRB; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 18:24:@166514.4]
  wire [63:0] FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 18:24:@166514.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[Zynq.scala 18:24:@166514.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[Zynq.scala 18:24:@166514.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 18:24:@166514.4]
  wire [39:0] FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 18:24:@166514.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_0_AWREADY; // @[Zynq.scala 18:24:@166514.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 18:24:@166514.4]
  wire [39:0] FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 18:24:@166514.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_0_ARREADY; // @[Zynq.scala 18:24:@166514.4]
  wire [511:0] FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 18:24:@166514.4]
  wire [63:0] FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_0_WREADY; // @[Zynq.scala 18:24:@166514.4]
  wire [31:0] FringeZynq_io_M_AXI_0_RID; // @[Zynq.scala 18:24:@166514.4]
  wire [511:0] FringeZynq_io_M_AXI_0_RDATA; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_0_RVALID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 18:24:@166514.4]
  wire [31:0] FringeZynq_io_M_AXI_0_BID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_0_BVALID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 18:24:@166514.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 18:24:@166514.4]
  wire [39:0] FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 18:24:@166514.4]
  wire [7:0] FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_1_AWREADY; // @[Zynq.scala 18:24:@166514.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 18:24:@166514.4]
  wire [39:0] FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 18:24:@166514.4]
  wire [7:0] FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_1_ARREADY; // @[Zynq.scala 18:24:@166514.4]
  wire [511:0] FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 18:24:@166514.4]
  wire [63:0] FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_1_WREADY; // @[Zynq.scala 18:24:@166514.4]
  wire [31:0] FringeZynq_io_M_AXI_1_RID; // @[Zynq.scala 18:24:@166514.4]
  wire [511:0] FringeZynq_io_M_AXI_1_RDATA; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_1_RVALID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 18:24:@166514.4]
  wire [31:0] FringeZynq_io_M_AXI_1_BID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_1_BVALID; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_enable; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_done; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_reset; // @[Zynq.scala 18:24:@166514.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[Zynq.scala 18:24:@166514.4]
  wire [63:0] FringeZynq_io_argIns_1; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[Zynq.scala 18:24:@166514.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[Zynq.scala 18:24:@166514.4]
  wire [63:0] FringeZynq_io_argEchos_0; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_memStreams_loads_0_cmd_ready; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_memStreams_loads_0_cmd_valid; // @[Zynq.scala 18:24:@166514.4]
  wire [63:0] FringeZynq_io_memStreams_loads_0_cmd_bits_addr; // @[Zynq.scala 18:24:@166514.4]
  wire [31:0] FringeZynq_io_memStreams_loads_0_cmd_bits_size; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_memStreams_loads_0_data_ready; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_memStreams_loads_0_data_valid; // @[Zynq.scala 18:24:@166514.4]
  wire [31:0] FringeZynq_io_memStreams_loads_0_data_bits_rdata_0; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 18:24:@166514.4]
  wire [63:0] FringeZynq_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 18:24:@166514.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_memStreams_stores_0_data_valid; // @[Zynq.scala 18:24:@166514.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 18:24:@166514.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 18:24:@166514.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 18:24:@166514.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 18:24:@166514.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@166419.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  FringeZynq FringeZynq ( // @[Zynq.scala 18:24:@166514.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_axil_s_clk(FringeZynq_io_axil_s_clk),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWID(FringeZynq_io_M_AXI_0_AWID),
    .io_M_AXI_0_AWADDR(FringeZynq_io_M_AXI_0_AWADDR),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_AWVALID(FringeZynq_io_M_AXI_0_AWVALID),
    .io_M_AXI_0_AWREADY(FringeZynq_io_M_AXI_0_AWREADY),
    .io_M_AXI_0_ARID(FringeZynq_io_M_AXI_0_ARID),
    .io_M_AXI_0_ARADDR(FringeZynq_io_M_AXI_0_ARADDR),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_M_AXI_0_ARVALID(FringeZynq_io_M_AXI_0_ARVALID),
    .io_M_AXI_0_ARREADY(FringeZynq_io_M_AXI_0_ARREADY),
    .io_M_AXI_0_WDATA(FringeZynq_io_M_AXI_0_WDATA),
    .io_M_AXI_0_WSTRB(FringeZynq_io_M_AXI_0_WSTRB),
    .io_M_AXI_0_WLAST(FringeZynq_io_M_AXI_0_WLAST),
    .io_M_AXI_0_WVALID(FringeZynq_io_M_AXI_0_WVALID),
    .io_M_AXI_0_WREADY(FringeZynq_io_M_AXI_0_WREADY),
    .io_M_AXI_0_RID(FringeZynq_io_M_AXI_0_RID),
    .io_M_AXI_0_RDATA(FringeZynq_io_M_AXI_0_RDATA),
    .io_M_AXI_0_RVALID(FringeZynq_io_M_AXI_0_RVALID),
    .io_M_AXI_0_RREADY(FringeZynq_io_M_AXI_0_RREADY),
    .io_M_AXI_0_BID(FringeZynq_io_M_AXI_0_BID),
    .io_M_AXI_0_BVALID(FringeZynq_io_M_AXI_0_BVALID),
    .io_M_AXI_0_BREADY(FringeZynq_io_M_AXI_0_BREADY),
    .io_M_AXI_1_AWID(FringeZynq_io_M_AXI_1_AWID),
    .io_M_AXI_1_AWADDR(FringeZynq_io_M_AXI_1_AWADDR),
    .io_M_AXI_1_AWLEN(FringeZynq_io_M_AXI_1_AWLEN),
    .io_M_AXI_1_AWVALID(FringeZynq_io_M_AXI_1_AWVALID),
    .io_M_AXI_1_AWREADY(FringeZynq_io_M_AXI_1_AWREADY),
    .io_M_AXI_1_ARID(FringeZynq_io_M_AXI_1_ARID),
    .io_M_AXI_1_ARADDR(FringeZynq_io_M_AXI_1_ARADDR),
    .io_M_AXI_1_ARLEN(FringeZynq_io_M_AXI_1_ARLEN),
    .io_M_AXI_1_ARVALID(FringeZynq_io_M_AXI_1_ARVALID),
    .io_M_AXI_1_ARREADY(FringeZynq_io_M_AXI_1_ARREADY),
    .io_M_AXI_1_WDATA(FringeZynq_io_M_AXI_1_WDATA),
    .io_M_AXI_1_WSTRB(FringeZynq_io_M_AXI_1_WSTRB),
    .io_M_AXI_1_WLAST(FringeZynq_io_M_AXI_1_WLAST),
    .io_M_AXI_1_WVALID(FringeZynq_io_M_AXI_1_WVALID),
    .io_M_AXI_1_WREADY(FringeZynq_io_M_AXI_1_WREADY),
    .io_M_AXI_1_RID(FringeZynq_io_M_AXI_1_RID),
    .io_M_AXI_1_RDATA(FringeZynq_io_M_AXI_1_RDATA),
    .io_M_AXI_1_RVALID(FringeZynq_io_M_AXI_1_RVALID),
    .io_M_AXI_1_RREADY(FringeZynq_io_M_AXI_1_RREADY),
    .io_M_AXI_1_BID(FringeZynq_io_M_AXI_1_BID),
    .io_M_AXI_1_BVALID(FringeZynq_io_M_AXI_1_BVALID),
    .io_M_AXI_1_BREADY(FringeZynq_io_M_AXI_1_BREADY),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argIns_1(FringeZynq_io_argIns_1),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_argEchos_0(FringeZynq_io_argEchos_0),
    .io_memStreams_loads_0_cmd_ready(FringeZynq_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(FringeZynq_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(FringeZynq_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(FringeZynq_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(FringeZynq_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(FringeZynq_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(FringeZynq_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_stores_0_cmd_ready(FringeZynq_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(FringeZynq_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(FringeZynq_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(FringeZynq_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(FringeZynq_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(FringeZynq_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(FringeZynq_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(FringeZynq_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(FringeZynq_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(FringeZynq_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(FringeZynq_io_memStreams_stores_0_wresp_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 21:21:@166532.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 21:21:@166528.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 21:21:@166524.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 21:21:@166523.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 21:21:@166522.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 21:21:@166521.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 21:21:@166519.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 21:21:@166518.4]
  assign io_M_AXI_0_AWID = FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 25:14:@166577.4]
  assign io_M_AXI_0_AWUSER = 32'h0; // @[Zynq.scala 25:14:@166576.4]
  assign io_M_AXI_0_AWADDR = FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 25:14:@166575.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 25:14:@166574.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[Zynq.scala 25:14:@166573.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[Zynq.scala 25:14:@166572.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[Zynq.scala 25:14:@166571.4]
  assign io_M_AXI_0_AWCACHE = 4'hf; // @[Zynq.scala 25:14:@166570.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[Zynq.scala 25:14:@166569.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[Zynq.scala 25:14:@166568.4]
  assign io_M_AXI_0_AWVALID = FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 25:14:@166567.4]
  assign io_M_AXI_0_ARID = FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 25:14:@166565.4]
  assign io_M_AXI_0_ARUSER = 32'h0; // @[Zynq.scala 25:14:@166564.4]
  assign io_M_AXI_0_ARADDR = FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 25:14:@166563.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 25:14:@166562.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[Zynq.scala 25:14:@166561.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[Zynq.scala 25:14:@166560.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[Zynq.scala 25:14:@166559.4]
  assign io_M_AXI_0_ARCACHE = 4'hf; // @[Zynq.scala 25:14:@166558.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[Zynq.scala 25:14:@166557.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[Zynq.scala 25:14:@166556.4]
  assign io_M_AXI_0_ARVALID = FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 25:14:@166555.4]
  assign io_M_AXI_0_WDATA = FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 25:14:@166553.4]
  assign io_M_AXI_0_WSTRB = FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 25:14:@166552.4]
  assign io_M_AXI_0_WLAST = FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 25:14:@166551.4]
  assign io_M_AXI_0_WVALID = FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 25:14:@166550.4]
  assign io_M_AXI_0_RREADY = FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 25:14:@166542.4]
  assign io_M_AXI_0_BREADY = FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 25:14:@166537.4]
  assign io_M_AXI_1_AWID = FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 25:14:@166618.4]
  assign io_M_AXI_1_AWUSER = 32'h0; // @[Zynq.scala 25:14:@166617.4]
  assign io_M_AXI_1_AWADDR = FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 25:14:@166616.4]
  assign io_M_AXI_1_AWLEN = FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 25:14:@166615.4]
  assign io_M_AXI_1_AWSIZE = 3'h6; // @[Zynq.scala 25:14:@166614.4]
  assign io_M_AXI_1_AWBURST = 2'h1; // @[Zynq.scala 25:14:@166613.4]
  assign io_M_AXI_1_AWLOCK = 1'h0; // @[Zynq.scala 25:14:@166612.4]
  assign io_M_AXI_1_AWCACHE = 4'hf; // @[Zynq.scala 25:14:@166611.4]
  assign io_M_AXI_1_AWPROT = 3'h0; // @[Zynq.scala 25:14:@166610.4]
  assign io_M_AXI_1_AWQOS = 4'h0; // @[Zynq.scala 25:14:@166609.4]
  assign io_M_AXI_1_AWVALID = FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 25:14:@166608.4]
  assign io_M_AXI_1_ARID = FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 25:14:@166606.4]
  assign io_M_AXI_1_ARUSER = 32'h0; // @[Zynq.scala 25:14:@166605.4]
  assign io_M_AXI_1_ARADDR = FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 25:14:@166604.4]
  assign io_M_AXI_1_ARLEN = FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 25:14:@166603.4]
  assign io_M_AXI_1_ARSIZE = 3'h6; // @[Zynq.scala 25:14:@166602.4]
  assign io_M_AXI_1_ARBURST = 2'h1; // @[Zynq.scala 25:14:@166601.4]
  assign io_M_AXI_1_ARLOCK = 1'h0; // @[Zynq.scala 25:14:@166600.4]
  assign io_M_AXI_1_ARCACHE = 4'hf; // @[Zynq.scala 25:14:@166599.4]
  assign io_M_AXI_1_ARPROT = 3'h0; // @[Zynq.scala 25:14:@166598.4]
  assign io_M_AXI_1_ARQOS = 4'h0; // @[Zynq.scala 25:14:@166597.4]
  assign io_M_AXI_1_ARVALID = FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 25:14:@166596.4]
  assign io_M_AXI_1_WDATA = FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 25:14:@166594.4]
  assign io_M_AXI_1_WSTRB = FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 25:14:@166593.4]
  assign io_M_AXI_1_WLAST = FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 25:14:@166592.4]
  assign io_M_AXI_1_WVALID = FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 25:14:@166591.4]
  assign io_M_AXI_1_RREADY = FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 25:14:@166583.4]
  assign io_M_AXI_1_BREADY = FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 25:14:@166578.4]
  assign accel_clock = clock; // @[:@166420.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@166421.4 Zynq.scala 55:17:@166860.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[Zynq.scala 52:21:@166855.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = FringeZynq_io_memStreams_loads_0_cmd_ready; // @[Zynq.scala 50:26:@166848.4]
  assign accel_io_memStreams_loads_0_data_valid = FringeZynq_io_memStreams_loads_0_data_valid; // @[Zynq.scala 50:26:@166843.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = FringeZynq_io_memStreams_loads_0_data_bits_rdata_0; // @[Zynq.scala 50:26:@166842.4]
  assign accel_io_memStreams_stores_0_cmd_ready = FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 50:26:@166841.4]
  assign accel_io_memStreams_stores_0_data_ready = FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 50:26:@166837.4]
  assign accel_io_memStreams_stores_0_wresp_valid = FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 50:26:@166832.4]
  assign accel_io_memStreams_stores_0_wresp_bits = FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 50:26:@166831.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[Zynq.scala 50:26:@166830.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[Zynq.scala 50:26:@166819.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 64'h0; // @[Zynq.scala 50:26:@166811.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 64'h0; // @[Zynq.scala 50:26:@166812.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 64'h0; // @[Zynq.scala 50:26:@166813.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 64'h0; // @[Zynq.scala 50:26:@166814.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 64'h0; // @[Zynq.scala 50:26:@166815.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 64'h0; // @[Zynq.scala 50:26:@166816.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 64'h0; // @[Zynq.scala 50:26:@166817.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 64'h0; // @[Zynq.scala 50:26:@166818.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[Zynq.scala 50:26:@166810.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[Zynq.scala 50:26:@166791.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[Zynq.scala 50:26:@166790.4]
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 51:20:@166851.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 51:20:@166850.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 51:20:@166849.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[Zynq.scala 35:21:@166784.4]
  assign accel_io_argIns_1 = FringeZynq_io_argIns_1; // @[Zynq.scala 35:21:@166785.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = FringeZynq_io_argEchos_0; // @[Zynq.scala 41:24:@166788.4]
  assign FringeZynq_clock = clock; // @[:@166515.4]
  assign FringeZynq_reset = reset == 1'h0; // @[:@166516.4 Zynq.scala 54:18:@166859.4]
  assign FringeZynq_io_axil_s_clk = io_axil_s_clk; // @[Zynq.scala 22:26:@166536.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[Zynq.scala 21:21:@166535.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[Zynq.scala 21:21:@166534.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[Zynq.scala 21:21:@166533.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[Zynq.scala 21:21:@166531.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[Zynq.scala 21:21:@166530.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[Zynq.scala 21:21:@166529.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[Zynq.scala 21:21:@166527.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[Zynq.scala 21:21:@166526.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[Zynq.scala 21:21:@166525.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[Zynq.scala 21:21:@166520.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[Zynq.scala 21:21:@166517.4]
  assign FringeZynq_io_M_AXI_0_AWREADY = io_M_AXI_0_AWREADY; // @[Zynq.scala 25:14:@166566.4]
  assign FringeZynq_io_M_AXI_0_ARREADY = io_M_AXI_0_ARREADY; // @[Zynq.scala 25:14:@166554.4]
  assign FringeZynq_io_M_AXI_0_WREADY = io_M_AXI_0_WREADY; // @[Zynq.scala 25:14:@166549.4]
  assign FringeZynq_io_M_AXI_0_RID = io_M_AXI_0_RID; // @[Zynq.scala 25:14:@166548.4]
  assign FringeZynq_io_M_AXI_0_RDATA = io_M_AXI_0_RDATA; // @[Zynq.scala 25:14:@166546.4]
  assign FringeZynq_io_M_AXI_0_RVALID = io_M_AXI_0_RVALID; // @[Zynq.scala 25:14:@166543.4]
  assign FringeZynq_io_M_AXI_0_BID = io_M_AXI_0_BID; // @[Zynq.scala 25:14:@166541.4]
  assign FringeZynq_io_M_AXI_0_BVALID = io_M_AXI_0_BVALID; // @[Zynq.scala 25:14:@166538.4]
  assign FringeZynq_io_M_AXI_1_AWREADY = io_M_AXI_1_AWREADY; // @[Zynq.scala 25:14:@166607.4]
  assign FringeZynq_io_M_AXI_1_ARREADY = io_M_AXI_1_ARREADY; // @[Zynq.scala 25:14:@166595.4]
  assign FringeZynq_io_M_AXI_1_WREADY = io_M_AXI_1_WREADY; // @[Zynq.scala 25:14:@166590.4]
  assign FringeZynq_io_M_AXI_1_RID = io_M_AXI_1_RID; // @[Zynq.scala 25:14:@166589.4]
  assign FringeZynq_io_M_AXI_1_RDATA = io_M_AXI_1_RDATA; // @[Zynq.scala 25:14:@166587.4]
  assign FringeZynq_io_M_AXI_1_RVALID = io_M_AXI_1_RVALID; // @[Zynq.scala 25:14:@166584.4]
  assign FringeZynq_io_M_AXI_1_BID = io_M_AXI_1_BID; // @[Zynq.scala 25:14:@166582.4]
  assign FringeZynq_io_M_AXI_1_BVALID = io_M_AXI_1_BVALID; // @[Zynq.scala 25:14:@166579.4]
  assign FringeZynq_io_done = accel_io_done; // @[Zynq.scala 53:20:@166856.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[Zynq.scala 38:26:@166787.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[Zynq.scala 37:25:@166786.4]
  assign FringeZynq_io_memStreams_loads_0_cmd_valid = accel_io_memStreams_loads_0_cmd_valid; // @[Zynq.scala 50:26:@166847.4]
  assign FringeZynq_io_memStreams_loads_0_cmd_bits_addr = accel_io_memStreams_loads_0_cmd_bits_addr; // @[Zynq.scala 50:26:@166846.4]
  assign FringeZynq_io_memStreams_loads_0_cmd_bits_size = accel_io_memStreams_loads_0_cmd_bits_size; // @[Zynq.scala 50:26:@166845.4]
  assign FringeZynq_io_memStreams_loads_0_data_ready = accel_io_memStreams_loads_0_data_ready; // @[Zynq.scala 50:26:@166844.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_valid = accel_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 50:26:@166840.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_addr = accel_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 50:26:@166839.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_size = accel_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 50:26:@166838.4]
  assign FringeZynq_io_memStreams_stores_0_data_valid = accel_io_memStreams_stores_0_data_valid; // @[Zynq.scala 50:26:@166836.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wdata_0 = accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 50:26:@166835.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wstrb = accel_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 50:26:@166834.4]
  assign FringeZynq_io_memStreams_stores_0_wresp_ready = accel_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 50:26:@166833.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[Zynq.scala 51:20:@166854.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 51:20:@166853.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 51:20:@166852.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module SRAMVerilogDualRead
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr0,
    input [AWIDTH-1:0] raddr1,
    input [AWIDTH-1:0] waddr,
    input raddrEn0,
    input raddrEn1,
    input waddrEn,
    input wen,
    input backpressure0,
    input backpressure1,
    input [DWIDTH-1:0] wdata,
    output reg [DWIDTH-1:0] rdata0,
    output reg [DWIDTH-1:0] rdata1
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk)
    begin
            if (wen)
            begin
                mem[waddr] <= wdata;
            end
            if (backpressure0) rdata0 <= mem[raddr0];
    end


    always @(posedge clk)
    begin
        if (backpressure1) rdata1 <= mem[raddr1];
    end
endmodule




